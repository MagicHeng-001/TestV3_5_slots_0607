// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:11 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hXbprmQnQs4JFb1NrMoxcICjbCGGN0MRm91FORk3t5Vz6tpMeEWvqHR60PgKiEIe
MkX3LZA4IzGv+sr0W8NNI0Rxc1rbgMxP0ziCBmCEkN/qmPwIWCp7qZZ1mM1DmNCZ
KD6kGDEmblR3dvszVHgtpDQUNPjy3SKVQ5IIxJ/M+3w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34720)
w2zs700Xc9ADEMfgmo8spYi3TNQhQmOXc6lC8ZeQ2EgssZd5FtoZdEerLy2jvtRS
yuqC8J9YJEcPX+hUOxP2Yp/nD9yEGrR9ThQqRtXjhjPAuLimxggghMnYXAQYrX40
ztXTaNoz6q96Ki20N5uMs8iS8QKkdYKxdhG92bX35IQDb2YDEN7IKNuUirO6Mh/u
aE8AyZKEn8+JcCVy8kYkFpIqhATYlt9SB/1/WYC2qZ/sQl0rKPDUh/RZ5bKblOIR
fZkgPwS7/7NHq4H+jetAJY0nutRLO4Po3x/goB+uHvMmcJGsgZbgkCADkYmI9mDl
MzQF2U6u7LAqcFBJeLdWFJvf3aSGfpdodsA+KxhIrwZXDVQQtOzxZZY7TPt9nY22
657sCZjUOBAFTnNd3BG3ckNiL71k+1kjd/LpcEkguqSIWk2r5Bz1bT2uc0aMhf8j
j61bb8nbFQG0sUw5oHyoIFk2NPg6v1Nv/pICFdZuhp4kby+OjfvmDvzgSWQ61LOF
mHzNt766suXzCBu2a+q/HIk+sIcoQq1tcbk6QY8cJBqP8OTAon3JLIihnJCcQKOC
1KCY0X+7dNzRfKipRytVVY16eFhgnQlathy5TWNURCRxpGr3SQCdT1mPhnKBao5X
0LGtPR6Ugt2xYk4c1mR1tC59nUP+GX4k+7ZWzZCs2dodHKMxt2UUoDeEwgVlpgcT
T/eDmbsA5zvyipOYwS/ixGPB0qyBniMqMkxhMA48X5Oyn63yC8IEPtgbXywXjuZ0
hHReG61m0Zj9GBxSWlO0JwxG9oQLp+GMcGshDGWl8EFXjYAcfgGuwC9AVUo1rDb7
YAd9ZdUg9kg1rUjMmn/oRFbXNFv3SKm0Kb1Cz5ytwSOeIFeRq7zIY/qRCUItBhPR
FGw2wtPn+s6o5QwdHBsOpWP+i3ywS3TyCKHBRKGXu31lrJRz1lFYRQNMPq7dmSmU
SrBezzezA81UIm2eqr85ugAZV3LbUr/fgJvhBufaF1pwO4EIM0B8Ua3+RUgFLwkW
lwaYj6umyOi7MhorCBVVvMyc4QfEYfwj5iwyd6Jv0Mql9UMS0CHgqA8uOH1EuhgS
2rJHEtjGdbYMRIxmR+pO7dSq9fp77181NoLgQHR31yDrYb+kWO50TK/aKDtGnfzC
cDJjmxa33ebYmfflPdvsbIOPoAxNLkUDoVA4Y2CWIimAlKK2tSLL30YhRVKbQBNJ
qQPmtVN3S/FyIjIbzrpyypOBV835uEhghkR8aOI0F9wSEi7QQ0aXuO3X8CJ72ke5
yXlDyIS1H+T2DPrnzjSrm/FpKIZaT+b/CRSAsIhZEbljLDwvev1CczK+TEYXtutC
jff7URdc9GbT3ZTsXzcHgY8F7cNphYek2TAbrvtjNEiKLDQJ0bp6GgIzaamvbeMJ
UWnmqDXRuWD5a4Yfojua65wurW5FU+HxfPe5TN9tIcNaVper8kWiDVo/BX3vETDH
hCv0309TCQkb6rcJYZNhIIsV1EFUmASeZ8WuDHZSrW1HsV59V6bdhCyyoWUD2IZp
ZTmst+CRH3zYf/G1/k6cdKuyeF6dhpFZiglehx/X3Vj6o6jnEf6fphYx844oVpS8
K/5vr6zhIenyXjy/tp5qukbxCImM0Cpdrt7TWB3K0XdrvCwe/oht4/ZoUHVXyiCV
XkkNWVMXNBPL2r+NyuUq1fPr8xINRjC7PFL3AXovrMWN/zPT2WeY3KwvuTiFM0oz
l1NiseerM1R3qcBEaz6gjLMDDkqFBMQenSLEOq8qPRTXiFwSgjsl5sFQUkX6YMjg
B3u8/NKfhodvynV1/h5/uWIc47xvGuAbGgr9BS7oT37EDBxJNGqTTE7ohV9fkjpj
zW9y5PDVixLK3l2WDkBCiTLNgQI3aunxbJ1Ll/3B5FggrG/8HuvRcDdm4rB/7lgC
QMT9dBkU0Xt8fg75DoEd8AclDiEWOWvF6TiHxnxtqi1HOK5IAzlabSFYwZUuj+Hl
S8KPeinQnuCKULFEPf10yjvtqO27tDSGpsn8QlbD7uY1D+8Dqzevth6CxnzeuMR5
pH4VFsg26A63jtvQ//4dn8CNEbmEXcBW8ZnjX9TYVmPv/y8SJtLXqajUbZ5/4y1+
v+TbTUuxnxfiyrWfJAUU2ysqnn+GjyShmvlpgGQX8PQuS9TSMefObofSsyIUZ7Ot
nF06glKL3T/doh5oLWQIfSq4ZW7BSo9WjIhbEhyqzPyIGK03UJCyIeOZ4a6reJsD
+H51w3/DWzjcq1XNM1UbY0eFFKd1hU8QaVCVtDmZ+sZq4zW8Gj+JB6DEw1YIhYBB
dC4jaGPki73ZyHDgQhrpGLwFhzWyQ6nTaNNGIPlWuRpHgUr7buEjcHDGAy5dNJ8u
sWLhkMZvH+3KRBQzZbIVkRCQ+cpP+9+GE+zzR1uuuVcpAb/iSVUln0qG1tO+ZPhW
yjk2IfZ3XoL4zo0yTqGJoaebuUtGTi1DBBa40SyNWSfQuXE5A9AqHuqiB7BspRs1
nZ2FSToIKCeIFxBU2Zh516NiRDLTLTH6grNLnGKN5gcRQTwHSHIyxDPRwPZUEc6e
+bVfCVRdW3BJ9dik3PQKA3A0ORIg1TLhXKzAgds4/JVTct6HFquRHh0qv2TGqfDO
u3mlcsUyU050rIo0YA62iGhjcgDpJJp0GFNJs5ya/RezFP+MQY/H6aylTnWx3kuK
SBGgBMYp7Ase0LqWgaLh7/He5F49rXJj88iCCc8KYPSyjMgYgtE9x7u+44u0VGd/
/YiCryrttDBLiIgEzTztLAv0jqu1kMKsZ8J6n0+7GwQEDt0DFDDyoa1IidcdYHCD
s+O7s7mg0+hVH0UXkB3LGEXXoBK49R5sZVFIYRGV+Ghw4+vUVNIfqVyULJgS1sqc
vz3fcN5OLMFzNHq2iCcrssvep5e2M4HoU2frrOTe+Kk1gdORRA+8eBznS4BV29sH
mO9BggaiPDmbWLcqVUUgAnB/9PVqrxaTXGXB1hi71HRJqLr3C69SKONH16qvp+fq
88/SeksF8WcHofruSth+wuK4cm+ueIjbGWZIb0VOtHpuPxK1CHnBGZWe077KdupD
G9NuIJTmg5TyAttrLtAnYfmv45eZaVCUXbZOg+U0CS4+xCFljhS+oqOOkojo2pFD
HxTcimqssIqhxUut/lJ7BwvROeTtNSWBNblD1wVFdOPxM8rIBhzZlOFXWG+66tcm
+GrC/tUH6ir+jBAB1KBxi9g3lqjKgISEcsrLcYdkXeksP2tX/ZUedj20HuPkvX7s
Y3zc27xM3z1V0uXl6NqeeRLN7N9atNfI7UNyVCwn7FhhMv2ManPOOytEJyxVx86D
sNaJ0SLQ3p9bt8Emnle6aa1ifcGlBgjVoGjq2wxWvvVoU9PWqW75bcgYHCJ7HD1S
yxR6WMJ3mhOR93sMZYQOysQG6fxSMjZCHrjzELdykIG4cJws00gWBQeK27I9KGO5
GqpBch+dIk+Sce7YiKaIpNyV7fNBKVAHHeWIaavLA383cWX2+OhmUODyF763xJil
FhQ8alvmvMM2yv5U+IFbs+dFNIG4mBtC3l/gswB9YN1evM/G2gDWyE4+9zT6wRni
5TgFv/ZHFNyXGY3eBpCcAm1y6KmdolWjZMuILB1ETIgpil89I1F6AVpY8BbUB3n3
/QnGwzJwmkdhA6f6eNptvTZl5ng22/pcL1lEx8gZCKqDM84pZxyP/U34DlT9paNT
BvgpWZjjMjc+a/mKvfUYhTK7zcYH7+xbdzKKatWkS23YsgXqY/nraRt4Vfp2jKob
ECTstjC3WfXQfbfvR+jh+l1lJf7dG6x2FAb+jj35Fz9hDToBD4LYtSuvU+08pXUH
gNx6QfCv5ZGOCYGEa4XEfQziOzD2jDPrIdFvtqa22ePZ7u0LB7UhW/gnAXmDeXMc
A4+1zSWIY1DL2M3itqEk4H63c/LoqKDge3mdiggc7Rw+lbwZevDcO7TAj7ph9yRY
B+7U9LyEJnNF/JqM5743SxwyVsUNPoCQ7C6BQcR3NO6yk1jtAQGBCbK2BEoEiRJ8
YPvl8hik5z43QJXaCBclkFQE44FFPPD/VqYZmp+VbjnIz71jOZvMXohAsIT4ZnxN
6SLTtz86C1eNGRot79DbwOkJjNk7A4OVMBgx6ERc78RL9hJpTvoZbwKyx8GZJFTK
lTP2M+5tjFA87z0AozoBWhiARs+anznRctxKFm7nBOZ5iN5YlS5Az4fvAa6zaffE
79/Q9O2ctgaWQ2ias2pzAeBOopPkGNm92aErbPsZSl6qi4ulFd2P1BW52npDhxrP
94mJwFTY1VbQ21ietFxYKyME5aMZUtDF9uJK2wz32ph/zhKK2KnwLHmgE/8sbUZ6
E8CdESBr8PycW+vEmLj1l+7xL4NtQPE+xRDfsn37879XD4eLpuybYscpZoqpmdhH
AeXiWVXm2+TXFfSgKbh61Xj72mCb7vYgRmvZguhsRUs3DdbcdSerkAkrqx6BIWoh
n/n9ngOpnfQIaBHXBQvMBBQht17eVuB/Cfgib8MvyPl69osBKKMsP5hJCVWN1Y72
rJkgbwEvA4SYSP7eCsGZFse7O0Gccus2DQM0zZ4OX9E83wbtqZm/SLPQPvCUEITL
tGUGzTqijI65K/Cj27fdF//4aCIdimxua2+8fkMFIPGXyG5owgo6vuc3uMF90fhq
OgNwITI3P8eK8z9xPFPH3HDTRKSmLA5NHDgE/hwUMMJOb6f4y/A04JHd7OnUqYlO
ldUPI9EOKiypwJ8UXRI9PRnNf3wBDM0vIB/YfUDENVjMGiOkGwzhWSpVgPhO2xR2
+SFcmRu9WYJu7QxDYmi07jb5YbNRvaSoVAc55BU9ptj4xYwMdaTgB71tRtVZt2ay
L6LP1rsowVukRHRsMVWov4OXmbPko1RrkBoLJgGq8O6GaiPPLJV17ZyeLXoui2aD
eJ99vyv2Oeq8FwItqF5j2ZG9D8ufNQtd7+mN+OqUVt6T5s3rh3fBKTSDjPeHPysq
IqoMk55kTiSOmvR4JbIk2xZaGlZSnSCA+HLFQiUFJu1sgemySZYDo8dEzqSMUL96
p+rOSWM9JIwZDs1dv8QE7yJNUO/lA0BBpnmcg/xDThBb+M1Vj32O4648Vfqcwlp5
VWLmNnDcNCqKxiZEB40ku+HtutrRjxTHc361aQKcyq0AAiGvxOb6RtQRcpge8B95
D1+OVhMy9NUiMHswfs/4UP4qdgfmdJlJIZ2jimVKUimhpK6xuC+WobRNdId01HR2
TKTMJN9kkxjvNemYM2Y9wOZele2D14nGNQfgaIdSDhWbXNXBzxbVR5IL5r2HQ3oM
/NlGrbp1E7XBuJQsx2RKji/Ap4gzCN156wyMVH62qbekUjcSzMBM6LtvV+4rejCZ
4A0v3B6a+1OXw0/cn5OOS31fXPRSrEw7R9ZJMoZYuDVyYvnbn1beTYLxqjG2p/S7
XcGaIRGsa0fW9YBcU7SSDmfYEJIMTrTOR+TqQC+Qs4YcaUago11q0cVhHEaoxYvM
ay4RxTitJFTfZ9p8eDUvGOBgcQWCLwP4DqHe1Z2HY87b3sOWaGqtwRCJF92gNX/+
o9KMw8PAKYL4X22gHyYnUnKTWsfjgighFEYBJed9VZMJ7gT8psgQNh76ujChAmfg
dJAerFYt/HWOUOCKzH/7fA0wQpOHyJC7n+AdluqQojdZ8F5uZj6DUAYQuMul3+J/
LCws97BuMP1Jb0PC3S4aEr6T5c/ApNP6bEyro4GCtAQ3O9zkPDaeEWfsnOoQR1wW
6rS6WKj5doiyww0O0AfE3G8o02mlJ0dLVZg7EhixhYQ9kUYJuCrt7p/oKQ2Nce3b
pf2qeJ88hx0L153GTZwsKDiangFpt6K1KEcKQhewRoaiNoLMZMuxxGS+7WHGhdMQ
rlByJgEQ74DuFbSYNlbdhd1q4/cdlC9V4Z6Xp5t+JihiaJ6AuhlddVga7IHbaNeT
VRmlb1yvZNmg7Z746XmOY5H7LGFQALKn4T9pc4mOEv9z+sjqY457s3DCWBDvJTuq
46jb2Eu02uoSbSBNlwHsgOuvGG5JK4QFlvzAwg37NPBQhavZLgJjXeYnjcjhar/P
Lk0CklgFP3qP6O0n/eWDGXBAwU4TZxzok8cpca0Vnz5dlm0liWav0I0I2ZjF6AkQ
PuMN3XUvAwYr6ih3CLQygqd4hlaUKhD2nZkQOPBw9GuiPssbsUpOF3ku3gApHoSq
/MHO0k2GWDHNv81qpfAZXhkne8vepSsArEh+GvQS91wjtFbllNByDR+Aey52XKcv
G1vkgdh2t/Ivu/nvdQ4/kFSXSH3NG2+15cHi+63jt/7+JQjAwA+keZxiSMZfDv+6
fCOALW7X7GuTf4UlTV8iBlMCd1YkEVULzEz3uRxAZRMWoWufOiuipt6Dk2CF4M1s
kHHa5JvQu+3Bpl5hj9c2rMxL1DS/jESP8rcMLB2zFJZoEVaE2yvL4Wz0t6ro/Y3S
Z90g5bzE9svI8EQudL4kx3hQLf2NytJliNbDjIEOoLzG0RBKUmN0CttKWysWJeOj
gqfIjxFSEziSDCEbUq6R349vhGAPk2AxiNIO0ZgewAVpNPevVEhVeLDVYde4kE/V
l2tWD1rDlEtqGucaNg0jSl6I1tQFPYnSXPggtKYxYPq26VE/68CgAEiFt/7wwxUh
SnSry8j3cC5Lexz57COK2iu6pxB3Fx/pZME+nIIsxcyF2qaqhaONG3mg5e3twRB5
4EGAQBBdJ+BROeL9MexKcGQzyiWGCrwjNWGO4flOZggpt0aPsm4E6rjBAhQ8WV4i
7/zUpEP0dIpSM1+UBZ2YTIMWx4pRZUORhTv73bjkHm7oGETmJSRAfxKyfeEn41ML
hgYiDTc2Pe+XqLw1wJxqMLcxXCqDyKGPVNc73zrLXgrYumCU2SXPp1hBapTJFG3E
8oo7Hht9Pvfudz9WP1WDm1zEtG5j+aKJ3JgaBP2C5I7Ckbsk85utlOBbcBC6fPBm
L3Yo4xOn7I2h/TXVRSvte19V27oo2tg7/MSYTIPQyarBJi7RR+7blrQlvWMh2W56
KLus8ptDU3p8eSlCPK9u8CbmV0LcznQS5LBjMNIFNX+A1QPn2BrpB791+5Zm8ERj
ZLIGP7FfTomxhBDs4qVrYmDo3wzLtbfiVgUe6Yt7uv1sziAjv52aMzPDjTw3KAMd
FgpmFbasQn8vfC+QcJ6mjSbukP4HZ1uKKMAuFST6GdgngNugXF4wjdr6pWsjzg82
p0avOAn4n4FRAF1xefQxnEXOYcTt0M1MeBLGhHdlyGb4bGYPDGN3mWO0cruACOJO
jubLDoSUL5xJszpU1fo3F5wQq7+eFzoRkeWj4IMtHw0rC9Ws+mmUkVE1Yxjh2GCg
D15dG6g+E9ZKpnXBuKqIz/dnEXi4/Rl89YSI9IwsFnDvJgR6nvIsGbkIVugEm8yw
M36dD3kujktfLJdHfl8jHdiKXAF0U4UXNGxKKyiQHMJQ8X+Q/Au9QIztZtsd0qQQ
xoeWAu6fFcew0krw8RlwDS45eXvfkqqe62gh8mVjcIhVabt0C/v+9ZShFyujPmg+
OUn38PN2Eq5PFqu01CXK4Hp+ynlLutN6VterKYKU9/a7hs6aYl3vn+UNzd69FwHY
BVK6c47/HRLUX9lrZ9Tuq1MhGkU7sOj8j2l0KlskFO+ubb3E/jrY+9Sz3KwhcnpU
E8GsAAyYNR0deckamQVbAKjP9YOhiTFBD2Sj1Ui78jwPLSC5QkLw0wROdjW/IXxG
KBgNQUcvvmmwWtTh6n9g21TK5DmEcYc65a8AG14YrHhVRbWPRujTBsg7IpWJr1lW
GZsqTqtZ1jZzbaZoOSeyDPtntfhWua8snfuO3U8hVz+fO/QTB3cuwz3AZHWpmRcE
Mru31fILDay6CHQLZ4/LycqkwIH15pZV4UryEEMOcM3QkyLHcdmi/heVmNatIQln
UQNt0FDHlTotsz8utQmOykeOq/5LeaPCy0OG0ajfL3IrizFItiHljD0r3TdrUjlN
8amAKddDIXc5NCesLf14Z2o9fdEwnrg1xuc17fgUrSJOaVOef7q4XoOIK11fjmnH
viVoJIz3+JFqC7xpiWRNeqdACXBraPTdBKtwVOH4vxNPkNbz+rvrJnKPtH+YpMhd
yqaBxKpA2SFfjmoNZMD1iqzv81WgQ0vUge1jt5D6azTfHzRHCOn1QH7f5E+H0uM+
V0sexUiM+VJP0w8GtVFPRuj9B1aifU9SGCqW88eRvIkphAoj88fzRNw8etPVjJH4
YzYJdgXcav7x9Kqv9lnCJqNnqD1pFjj4jfUSabH74NYa10a2pKGtxokxX9B7X/wv
sOInb0zh/JFhE2OsPEoY8m42W1TrA1cAiomohSYoummbrPBwvI9DbtlXk3v54Ssl
E8i1kyc/RUITIFJSJOz4j02X9gVpo0m4TBsvRx1fVmU8brYZPaHxJpUUJY8asEr/
ESVxJqq0vRmwJb0owZXjZwT25HjxXALMjxOvd1xGVQVMW5gMl1Ad9PQ6RxEpIJZp
JLRU5EhtWeGvhHtX0NmiWMZXvmrvYT3evBN9d+lg8yp7X/JaM85V2k6ebl7bZkmR
yKWpXpPI3JPDCmq8NjLD2gM0HPFAcNeKsNAJaqMcZBh30ZylciDGF74Bu79wxFT5
oxEh+RXxOPLC6Am5DX1Lr6aYDerbe+Prk3gH0wiq54cVcyemM4UScExv8UK9ToxM
Epv4L82/vFOlwb/qJWlSx0oYllyOuvbMtKOKMn4Hrp1tk4DwcCtpkmeQGqwGSDu5
VQpPfYjBBfLkgWYeOBV9vz3mVObFB2Gsip5yCi/ourtC2UGwhhCpa3nw5z9qNmUK
u12LyN32oqKUXFUwCDG0fpzYbaaDW+mDg/K4K8aTvLYFBjZRFjLrHLuhhvV4eE0R
X8MUamCD6L2yEKuIABJktEnU0SgHA/VKwR2gTDcbR4rrzWmE3DwZlJEkTFrRjOFg
CZkq5kPTfCiw6i6xiMvLUzYsLyX8f9Y7VOC5kc1hQzrE5n+FePTjmmYM69PTMPbe
3Koga83R8JdCJooVsDCuPNG4WiSuuaZhdrJOxseXOz0BFe9PrK+4njoLi+gdhZFS
YWtL1I0EI9DGHgNyhRWcfGlMHxoFlDBtBa0rxc29+fP5QsHWyYx7F70cPIUxAY7O
suF7mcypNeR8qmY/rLIDiObn05qEyxip4iiH1MmABPb2ZxoXERMeCQ3L9yhb88/c
f2S/z9eXxLixpOWWJtyPWgDZC9ea3u4fQnftEaggSfD2dYMYnhXrDY203yNvVDnU
uT0YQ1gWkWD02RXIYiTePbOJd9js1vKGl3MnJizFsvW1hSZXagS2Xec4F7aC1MGo
GBqQ6zAREEbj9R7De5hfsRUsdy7hVgllkjt7BYJz/Ll89a/VbtnzYh3JF8kmMpSI
vsGX5CSPzNxcLJsQA8hHw23Ti97XW2slqIsi4An7K+rVD0WOB7dgMUK+UlOWUb2D
1pK6mSNbDsOwzwinwqQYGFG/5f5cP88HvPhPi6H9+428VdRjwaqJr/Lncklt7PXP
cfqGkBI6FxT3yAk68itaE+PD2y9sAy7VhVoy8p4LesJT+qeFarY+YqQvqgsbdq9Z
7n+Vz6YbFcWnGygE+uD7s5dMqg1iBucGN7U2sWvm+BVhV+/nnilUIlY/A7H2MzWW
9e94J9C8wFMHjWeERkfdrQAPm2nXjNClBnQ/MQkmZDLKuCxl5gintZdNPUUrtXZu
B4175OFF0iVBYMsL1GM2QY1O/GHpmfsGgBNjab0tbC+oD/qdWKjkuBlEg2RUbJsV
g9scSgNcowzw9KUe5Z0kUprK2QRPy+bdvlzuNkt8snHfXbmljEvVV80Kje4MzE58
rOAkgvUxYV9yaT9JFHIcbHFqPMI6SjCjGeuu0RhWcAzM3JfN4K+lsCwUhVFUDPPw
BWVzQ4ueD5LJMfD9ynrwTu/lQuUb9RAepHfHsOQ9AKWw2A4OyTVlHDWniHbniTPr
PK/7FjF5H4P6f9sifGHH644mtYtOohjdWgpoHZwpG0+sdZ56gP39kfqtyRWB7ikP
rS7zuYCEDs1BEfstVUEIPflqP7dF/u2cH72fZTpTd94AMAq5UgC/2/Qg7ydbYskg
5Sl1DIHvnZyUSANVHzf1PEs7vcrcCE1Z5j1v6htmZi2LBNgCu6mdpmV4iFDH1OSJ
a43Yf/m1XDKAtHlwnLs2ap0yWGyheVDNV3CcwyQv4lOHpE7QwrUPqxQdwNWTCwxz
AsbgBcKKgYZPssBYV4lQEouyar1wwghplt31g377aX5k/tjDr2xz2KGIhgayvPaU
O/5/WEi2e/OOIruFRfGcMoB0tCK0F+tCnbmkQZyhNN4OhOFwxZzkUYcjIGf14TNl
/p+Aq6bhoSNN1TOV18Gs0y97gio6CIWOOX0wt+rD3G7AQuLfO6np/veoD/rlCsQJ
vu7OOYUoTM4yuKPxr5bxNxIJFtXSUaeEc/XM7xq3hJgLjZr5SnE3OQK+9rZj4wn3
R5vLlC6S1TBjvjp3xJbLCOnnp6naMD65ttuCkOH6NeYIqNe5jPrEmQao6t09dYW+
GXW0KGdLWQJWJGLoJPY77chTVVQKwHOCf0HjH2OXPM/rTKxmgEfi/N+4kW4B41Hb
5FalSHOmaRKDcNkYE/VJEuGGDucfYcESmufTTcOaC2JBfQjJ49cn6tIuJyr5Ogq5
aIeE5qvWvc9kNkvaqj1UZQMwiNhnZCYkqekNjUajx1w/Z1Ub/MS0Nc/Mp1YckhfT
yIIo67miHbwRPLj7PBlBDdr4bs9qMeXkaikrKIUN90GrHzb5XlRCIOaFomOU05oC
QVprCel10IQHlEBWKfVxA6H5WZ3Op/xGGWLou2IuhhZWwo0UxSUZfFJLDZPc4ylM
/kNwWAXVjS5yYjGDV4mH27mfr7SZKvOpo67gOq9kSlTvrACResKE4SxkzzLCA06U
OhrUOYsekTHPvKBKIm7TfC8NQhdmpv489fzdDjl32M8ElGtOJ9W5xAj/yeg8UiS4
16w6Ro6tEyqJmQfhoO+TooK2txPZL1jOvzpxcdSsC57ZWgMdbCk1/DRIJ7gDqPXn
ZFCWZiLaYkt43FcLHIjyMi+ngjtoH9yNQbjemVEJOozg+hWNhHFepwv771hjwbbs
cSoGPIAorSB2A3mepygoTDT9pQh2JOyXjJ7IdgHsl/vTIwLKuBLAxO7XaIrIQhww
phex//VmEear7Hx4JUsciM8pO0oGtpkcXY2RtV9e1WKuH35DUjO3o9AePD+wLIdb
xJZSHH6jOcY/ctW1TnDGBLxnRvQz3WEttDRPisHsq+/RM9+SVGdUW+1iyl1lFWbI
O7csvfGxfH0AqBGhwQ0y8G737AvZkHFlBJe8MrE4NBNzcaZnbVefmKbgx/S//p2M
4Byd+to/IPQFvdFeInlTZI9kPFm3F/1CX3ip6gVBODcQJ40nYIo2t6Fqi//e1e9X
cnx7ja1sVx3ystL+5oCGDZxQyn2Pgkq8h2edEcgbqueAsR4M2AE7fPLj+uFI1VUY
AjleO3fNkAJH2Mx/EYlrJA+rEhqeeVYlx1/YU9QmKTaUcqYdMtVqImi35MRh+OJG
6TKsarF7EH3PR+E/BEp9LLFbg3+2G3u9rN761J13xh7YLywVCJuXOnVG8Xv5J6ft
xlcV2TX3cv0AmRpxy1XuTa5xkbmC5CGnqGzJguYn7ewfHOKBuFhA+QfACcR/mMA4
qMlWM9PxH9jIiVUhsWQ/1R/cghITQSp1l4XlHiDKcWc1hNPaXWdKsi5G4xFOn2Ww
3rA41mumFcXf87/6Z67Jr1WXmTCTQgUsgDXxMjo2Vx8LQvLgQpy5BZiQH3wuLuax
45d3vTG6HIV+QGfWcdnxxFUBV5oh6ff6SRgssGDh0RovkhvByaD0PZbLS7u4/16A
N1lWRsiGCVOhcxk98ja7TfC1j/qcBgKI3u7fhVz0QDDRKOxeovkYSvQ/0bsnJRsB
pc7PKeP90WBj7p2+xdzxniEXDxZuVlcW3dzwvMckH7eDqnjvgPjhAPMnCYmQKOvU
s8q+81q0eIV9kpe2pck+30P//dK4hwsWVsBmtwiF3R+FF+VvlXO2oysf0ARH3UI9
NMsf/pxlTVqlIqFdEi8xH1O3RP7K5ljgoNsSbavPmKRj6+gzvk5SRbqsaVGqu7K/
nmXyzp0VoQPheGExsTLvdr9YwoRcWHT7c5hJv8AejvYrL+LWfB3NaRTE0OeZ8kOf
hoULgymS0ZRF/IcrDhcvujb7iCfP410Fkn4Llovs/KHhLU7M2yMvS/E3afox3IUR
BOiL57j0tOIB/l/He+tgaOa0HrAt0SUmmLtWIn/wycvoDG9YGQDw9SfLRCHcwUWj
ZXI7xVWX+qy/75fWZtrkgzBe70ynxb3jxWDhVc7jH3zFUKrSDdFYT2GGfLIpp/bN
gjhZtsu2hOaQA2cTf/HA1jpdUWwVaKN0sUP/z4vyYhQjTrCdAN+65qYzdkQ/1cZ5
GSKftXjoFL2K3ehYmWcwnQ4sRutgE+sdFTBwwaVK8dSLoh58aKReE3/asAOCRIXA
TeaQI720wCIlzXndrbMpJ7D6O1AheKt0T8+enVa1KIOEwFaq2OOJeBB1vfdRUCxU
y8NnKPv6qI/ioLE6SaEvEoXVHBGW3Yqk9rdDZGQRWqEtXU+4crSpxJ4Ohd1viafw
dHsOPWEkLO6kEE453taxpHXG1N0q01ef559DvPoxzgaMyE5LV0Ltopx/dPmeBfoP
1mMuu77z82PjrFOrLIJBaL6fjKHcU7hLeCDOpuPlR36clt6fnfkpL95SVttPSNKo
Eof4KrZ+5yYo/o9IF69a49Ym3vrO81XRVNjnoW2x7vl5DOABi/wiVtpHuco2FTen
RbOuSsGk92in9fG7unIp1XM1e+zTRxkYA/Xn1ueHowkWfbRfw46jnTBxg9OtYBzp
pXsZ50WbuworMYaw8TP5OfFP0/kvQ8D5yjhFanbWwB1EKwUESgw372DXi5VSMN2J
YK7DiH2k853u1b92sW+f8fdCM57w5hCN0vCMW4gnI6+LOpyu9BRj+zSrEu9HU2jj
+6uyGYJgG998LftsfWoTvGMZkN5algdhKLk586X0PFkNPw7C4/8kKu6kDSQ9B9DK
eWnbxEAI0nxERoWFf/KOEKtTRAd5lico57bK9QoENj/5XcJc0cOs96gpcQrJ1LjC
SJ+d09hyak0LtW3pBdNoBTLwXLwiaBpCZi2mZL2j0Kt3dP62+0DowMUCgGJftxNC
LFjhC+kdPFz6yLvB9ZXFaP1o04jkgLB8VhsXmYC/Cw7YpHRiwcXcObQzcyQ+x+z7
t5NiVkUqDfDsohKUhTE0kjh59haH0qqWssq+2uk8a1pv5nWArqC4F4j5svMt1eXd
pSobKveRDC+7Zn06DHzENvfgLPpufWMwHOke6fmI4uT5ZMflX3t1V+8auFlwKwuu
GxUUV6BJiw8GKgfWKXsZY76DJ3nlyT6SJjk8jtn8/INe5X8wJVllgMFWFKn1HINa
+oQiRTsC7FhOOJc1KdSiGKlxP5J5aHIe6EFEk9TRUXLb0wFGEucorgyAcuu8Hqra
029cZmcMDssoCAM64dYjgL5eFTuE4ZN8X5Sk7L/enxxymMgR62fYXr0SIDjv9xK6
iRRxRfXTRTKQaP4qD2u1xVxxcI5MiFqpz9hnE09wns5/E4HYuYN8Qa+ThBwNC6dw
j5GJ1JL/kdJ4tQZbhndRg5jqTX8qx6jKXx38GjwYvtqOckOo88w/gpVY4KQpuNPR
g3hwsLtoZzBsMImgIl2QIduGOLipzxiAAhDfv2L2aHfF+dRPEbfeBOt07Y71BCWT
q4pGSpLqFph+hRbJMywUjuuwFojgFcXoAXLqkTi+GV2yxy6K4McOEgiQEeiAhhEy
rOQZXtg3kZTVzhE9M4w7mxY+3ibZF/vlXgHFhBwSCxp947RhiichmzmtsxLbKtXr
XfF2vC5LINrvoyTrchp+yH1TqxyNXU+EA5T0QGDvxNhs4S3ZbDqKnhR3u90CDwTE
fdrArJ8UCiTr1a7u1mfg/tMnCBYfJKjZcr0wGtOYSzRuutqGCMHAXTMOQrXwSL4U
LJjcmgEvOfF9SDpCD8qRgF+fHNxudiX3WSLhRdPeuu4nD45MIklsGmy4/AbxhQ85
AqRkXf5av6w/04eK4QQAsBxo9hJWCr1YgqwH6W+ZYWg1nSqLAn510frwl+G0bPXN
cs7r3ZwNgtNwE5zxUudxN4Dtd30yUMFoyoAbVb5qgQv1/ybrCzeTHFUoTiUzp4D3
wOQfzxT414/rYrYkblV3Lco1IF4Vwxc6ozbH21R0zsClcpqRInt3K0KzJBmNLxN0
EMIgS5AO3XThLyTOovD8AIvUu4q+ltmbmP/t0dgtq5EvrOFSZ6Am+nTFxAK8apAc
aZr2NpMUe9TudjsbFFI/+d54dp+H4EONcxV98n2h89+fn7MEXOkFwEcOqRFK2e1/
/n5xUHhGH4HLv4PXeZveUxBwAZtNvsHq0Ws0YLKqDA1zbIs3zgjbjfk/chCEIvpX
V3jgFfFoyVWRKFnVBV+/z3NMPedLmu865Ubj7R89APa+aY5F/0lgt1KllY8CGzJV
MdpHtaFagOR8gWxHQ3RYnU2LuUIbwgJ1JQ0PI1Wb+IxgFnA4cZgxU12SM5lREkwS
6p9GB73Qr82ckTDb7WxUtTygR1V8pFWVGLSlHrZpA+q6ElnjbCMDbJin+AgQ2jJx
K6F12gy1CpC+okjJGQMgRaffYFKGoH5nJ4QTq+Yw/uoS5qBMPi8Lq9jhuPa+tB1r
YsVZ9x62tGvg3KE3/vF8L2KY1zvdL9n55dWcRnHMGbp28+sJAzKm+GC7xPwHV8bM
yEp9zGzdlGc9Q676+LqozrmxozFzTKZ8pEx0nxuvIKgCwBCnW/AogT7Kw24XVOLI
umLggZbjkUJKpg4y5lktMUZGTt7Ou6NE6exhD+31YAG260t1LoQKWSvXWSWlS7zZ
Qxr1mOBWWfGp6/V2j9eXGHseCUopPxCMgF0qlbbOd/8oZCrlhQYzz8o+q2anNdo1
RLZ8FBb09QTJbhORDs3nosCYMKWOHG0/l6oIxeGwg9IrIfrpDUUGdXbGsjvVJHFt
hDptcEzDa+z9MgjTsdBNwfmI1NCH1tlNq92FQnM2cxhXD6gYTrOTljsNuUoz11hg
jrgqMsMpweQQoPtvzcpGbj3czV1Wtzmz7ITn83erEoGehgiyuz3ErTzQbNRZQtvN
wmTzfAvfKlqqXAff0ezzPFL2ZOAggJ5mNEcVaHpfQ5Ri9cXQKhXe2Ad8MRjndCns
ppYfmjuOWWnQ/aQns5JcHkxeCfEifAhQuxiC5ZGG4FuAXNe940LIRR48KM1xMYvo
HyhND3/r0HW5+pS6jj9GDtD4GljZhykcrEpeGBu/Dbb+ffhG0vNPz62vutVLG3z1
VIyzl4zkX1cpxBpwdvFRGH7FOlq/A/bMJ/GFmQgaY+raj/B9hOXkVaXD6th1am6F
SpZpOT4pdaR8DpwM5B2I8CfHrRDkCIptsi9oTrP08bUWX6o4ojiIfB3+0aJ+wxwV
zeY3rS996svEZB7pYix0OWKNdHlWzGZFjca17wYzCxDRy2w+s9hURp5d+N/DcGgZ
pbdSyjNeQcdir7NL6e19KqSd1KjY2ZhzjP/09UdNSjENfPrN9JoqEKrvdiu+UPYn
hMbd5TBCEmLsUQQ5IV6RRLSF28tuZTDkE7gKRCEtK+fzL9FRxy0d6HDMRU4if+54
yy6jpj46F3RvV0GAAdEIpgvXYvTmUM+k1x5w+pO/gaZsG/DWT7rkAEvQPiu8RJlL
Ncpk6RmUWzxzjxIeJ+yRqOdlGCOSE3pdmS4hLwc1vS36yzSoWM/iRPvyVkQO8mgu
+nDBeVYGeRZQODbHWvyGy18cNrA2Y09i5y1y7qxXVyZZyVgMRdVxCiK6Ub/0sQEd
ZzVmnVZm4fx5jw0q/QMZgPWY1BWre3GGi5TvMZj/LDM7Yx9lWQHVQJcf329vzOCf
LvGPl64L86rmygCE8yLVTmhI84Cgwjc22ZTM4G8yjl8ghgl7wQDGOfi5e2ZoK3Gu
j0tU8stDN/cE3jTuhDTVFkLDn4AbJ1KG8ToS6R18ojnckHiLAifjSCfoXoYeZLCj
+xTXu2rFD2vq9f8oxiJ5U1EIY0lF2rWrKqJEepnthhc/9x6vim2nCYdKN33+asKw
t5KCjsuRMe2U95SiagFTfjOVD6YkPXAxxPkhGzdJt43IX4mwxWHnVqSUp95GAVs9
lIiq8ONuV+xFfVjlnbpGpJUCtc4vcpIXeXvLbGg4q3AI7D8XCncA/lvaYuJzGaH6
wFgDGOuANURPAf9qA9UmwJORL2EpJFW4JcYpJMpu/PmtYHqFKE72a35hROYzTgG0
szyhFSP/+SZIUaovUrvE3wx9sxtc/s3t+4Y0TtA7Lt8rDONhoMVvVxSA4tNjlbfd
93KuPJ+yJaNHJKgOrvOsGQedmGTr4G75Wx2vDfRZ1NLWnYJd2MZXjst88zurZa86
CwLA/u4gZX7HME9B6bq3ossfdzZ/RavkXFQN6kJU+NMrIEamKtnd+UHgB3GwM58I
PrfMw9HUMzGyK9rGgkU77eSkVEWtdOfMMkitckjCBIUbL5piAPI99liQLPawwuU0
K3GVQHg2Ae4elUS8o0UQo8wCu6MK6yM00NcAn3z4fG6QGDkQZQz4KDN6Eohhpkpj
qNBiBYkj+Irw+Cf/bUEdEg1hfPqkkEm7Hg0KFPQmJcOn2rKaUYDjuWL2SyvcXqyB
ZIe+gMaC2g6oJOi7YWk41/Vh/BH5ygGXozTQHy+ZBa6rzp8BLc1cjXI1CiIlpTyD
eIq2at9BpwV/+mHoMzOZVEAN7lZnF+2we3uLtL6GCinrsiEaaultvxoDlimcp3mO
KqEO69XhgwNvVjHbsB2fWGYmc+LtE9zqbK18F4eUQW7enpIqPL8RbJCHnl8GDkTA
kqIEDebdAfzxhGqCPyWHcyYHsoGg55XmAo/8fekFen8Db3rPUDlhZccFw1m3N7Pf
r4SfwN3T4jyqHOrj/AFJx6ZDDTklC7NAdndu1txqQBYhNInI8zSsAkGf2ZDXfZi0
YpJVRGQ8Acqs8tRfoEPeI3Nw1hEgf+S8oYWrLgOsSTWQpVwJcRzp78dw9phKiSZr
dJYehwbaOo/LzyywW9yK6Nd16kAhbYsIK2UG2otK5vpWqPCA5cP0JLRSqXUZppN7
K+SfeI+WfdrUiyUgdcYl0wfdruGAuhiGgIpG71mQtJV8TJYCG/gxEhD97nu8qDQl
R25Y/2E6zL+sx9vyfPtwqKvms9N2SegLGdjA7nB/gmnVBmMKczUlrtAIQlKllLkI
hPF5cdEvWdVh7osvIkoNswLrgDytlr6SY0KJ5v5TQAcrjmOc/mDuZlBrbWQr/Yoo
OY7TaBsqiM/pbmq+x/8B+pqLMRrlhZFbnAJLRD2HeaH8x0T8IZJRyZTEpCWlZZCG
GzpgurP3XrcaOMngDMRsxiljwHjTo/P7EHnNlfVwiUqyhXVwkTyb9TZwTkBgf2Ev
nz1jxrzysqYjn/3srx05RxL+nu6Jtpz/PBr4iLsz566dCl0aMXJp7J0jPi+HnihD
0gmUfEBcgTkp9/HCUpl2Xu1CCXehDHEnlqV9styxzYj4AhfBnj0U2NMAPh7LZ29d
buNleolqK1h7LnlXkTqc2WFTu58aRHhzzYgxXHPiFaDVqIq/iYu15k0bmc3vtIF+
iWaXwHOBbG+MszxxmMJ/bS9k/Om4QfQsq+FGp7XD8VZ016po+pN8zmt8ZVViJJTP
QQBQW5GeUJGpSavjrQOfyiORKpY5KY5zqO3qu6pSjJrjko+W68u4N8hwuTJsuS72
uUbD7hvsdpCZ9RLn+VUc4/xwAcJF1rnQf5H3jWDHwTuCfK2F2ysrGjtz9oNcYNW2
TdftOBAjn63rWfRKpDDYH4hhKjOlO9PDM/mMiX/WWfnpEaZ3o/R+KFnnWhSwO9Id
QXPP5ATbpLTYjg3TtTV/v1LJj8KvIo5ZuEEAfJBnRllmHS0XfpVdLwaY4GCL7sf4
Lv5a8VzTFkSWqzdKBgsDckRhY3H2zmEzAFHSOuMBTiGP5tx4f0cDuCizl8QdPaF6
AcC+mQaJjvaTHPxtRAbKWQK8SpjpKHI6w/mxf/vYfeYoz1j1boJrOwSFe7opgel7
M5PdUTf0E6DX91j3DMP6PFSoi5+O8pGSakFeKBR94NR9E+MZeY5rY5TnkuU5XpTS
MSQXcRSIQjatENSlCKDW5xHU8mXCGshKflJvb7VZkAL7xetwqUjIVtLblCx16ynb
JjUhjGJgx2S4Xi4muh+6iwKip6MTcN6PzuwwxVhcW/7LtIv7Cr6+quWe9gwnQ/z2
7WEcJYaoCX451uBx81jjeuy5qP2M6tvjUkYKEVc5iCG1VBpz3p2OZvs0JsHFMx6E
MSWiFXJvmCGgBl6QGne/7JwepYAPbigpOFdIjygOEJHl9l1Kpuui+W7DoQq3gUGH
TFgYGJdhewjzgBOYl2PDHSDa8V68EggXhHE1J81VdJ6aEUtyV911ACfiaBafeTcT
uZAWn0aeiF34XVZQS50onYZehV8X1/TyqxeLiTFwUSwkuqnuUswOgyU5xaUsEtK4
6wm8Zh9ONz2TtaW/xnwTzXHI8k3JAFAlmTzff58NC7whb6qPdYiJ5lpbLV9POKxj
w7NTg0X9UuP7CgkMzcbbOgzPaLAEyer/QBvXR2F2Qkwy68FLzgW88bF81d0A8XMQ
Yr+zyaUX6v0AwImNoqQdikR48ABtywWoJ2WB70CcmZUHTxU8oVhBnGz3MEbSAy8q
ugeEdoaffQta58d+Sz1wUkNqMpTJUB3kFvoyMaiSLvJtz/s+5nTcYlXWbRZ3Bhh3
odR9xZ3eO6T9tT7rMujo2+WJVBJTDJ+c0abz3ebmLvHgv6150D0v7oGPKLCrkrRg
ZwOogWXCbF763y6TLq8A7bgouH/MXj+Ghh7PqFxKsqiSF93hwb5rP3uDeHOaUEw/
X3YMyVI70IsZGrY6HRJChD3iSj37pbfBrWkT44ypp5uqgFWy0VYMhMJeC7NcLYAW
yx99eIzMo1a++4eXT9SHYBCKiXpMzOezLKUqIWoDNLTPDYCywEXuFUh29aWikYnb
Pm4q43X3/Q+ngFljCahOsfm0nlge0+JQJCsCJpKk7ERO/gV34w2cBy8gsedWkLh8
Qd3YCkcOeB/FAXWppBgx8xNejIgFYg4mlAx9hsdil7U4pjsr7rRIOcDtYTsP8MQi
me5oHPPd2r/7Otzr4uXFML2Pqkw8RpaLJ1NnLSpaxSgLe1Vf36epo6I6lt718FYt
UK4AbtcaFJcvALGv8hpsmTcXwOIVM+qd3RiXnOwVATKKbR7TUO+zZrAp5GGls9x3
l4XLK2JJa9f8V7FRi+aytMioC9rDJi40q4ebUfKI/sY25hAmGz/v+wiyDq9heB4Q
IX4zq2gaqaQGQuzz3sWDnwmp84zuDuYCL7jEqkf7VRbKm4Tnpl9rjYs/KS0dLuPY
JSDtiMPyxK+U5VcB7f6Dxai0ZiHXgEB9hkwN/te5/+a4GKBZgBftDG3EbBTVQVIj
Z4/WZHiS6NN54t3j2LJMWozEjKLl0sU6cn/5E9gjOHkcXyji6t4lzEWOroLWvhOL
oxlaOArJizfmMvfk1bAOx/wsNiGITyElmkfsLHvIj61nFJhpWKV0KIKEY3iVgoCl
GRUZV2rp4pEHypxBvkGuKbTc6jujqEQZPTWeQ3Fi+/focNt9sIqLs0Uo2AFarF4o
8d6TjXB6XPU7Lyd1m6OWFtJOaYtDKfXxcLRW8vkxIIA1EHhTlNKHSJ3iHh473uid
CFOARQ6vMZzeibjL/Ha1CDoTJZZT5URLwlPVIB3jFu2tFDOzJ4LgSZL5saF6HKQs
LOZVk4FQUvLDUo49U9ze8yOw2wrIT/EC/TG/MyEWDq5Iixmfa/jG7OZgAf5Ii+Yj
xWeyanvV6npbq42+Z1Z4qdnBtP4ezCqsfXMNFnkNH9tR6Ap8Fw3fSgCRhyYUHGYF
rnrtAfTFb24mPp8MLFd7CIr7NDfh339cp6q5AFYErjLSqYYYWDrnM+n2oi5HKi7r
TzuecBQ0OPNX5gOGInxJs1hSEgskjXqboU09eXKEnc8TKZQ4ouF2wfW9yUjPNpbo
dWVM1oGKHr1uagHktIbtcb0+u1ZPmQ5FS0Ifnf/hhBy+a6Hmj8Rv7ZmrkKHO2Oir
Q+ZeE3/WYaUQMsh7qKh216dOEP/lJVCB3/pNqR9co1K+olYCVOpM0sPfr2YRrzMt
okDtwjLSWy+cFNcu5jSvB5O4A3DJhUIDuzLEYwU02sDFRixC0WEUKoEUfcwxHvmI
Yl5VRnlSkQ2Gudyy5Kl11Rcc2dikLm/H/lxw3mCIeXW4l2RZzOuRZ30eO3WZSy0U
pJbZUXv/bvGy2ZimAkBB9jsAxXPEE+lYjTUaWGFiE2GiTRUYTSad/5V6adW5viU9
hJR5mveEe+b4cN6aVR1+8xdhEY22pRvYvKkBzKoGmxaTAZcJ8bT6f0NFk/ApUqTW
1EVA8rRyxZls1OLxGT0dOTBfddEbH/Kkw61/T0jsb13034Wvw62FlmF6uwinTGhb
3IVAGqTnuw+/+0ps7eZwAq/g9YKewTOBJjSjl/6/geuRESg2CVY0oo0zvYsabgF6
m+4EtcE8+13VeCXWxgeZF3do8qwkyrg1tdAq+2iww+bdOLUNE3TTt1K5OwbeYBX9
Vi5cY4bs9CUpyRdjYzWVc3mt3baOkOE7tfY7ln4h6x/82YI4slJNN1BbMdMX15zV
aldvuiiEOYuf1IsMzbKSrxUk/foMXXFBfljPaWztBdy5kCpANB5fCVTzbRhzyvft
Aswq72MNg3mLSux+K6DkIjp9axRdLTsw7EahxhsLpVTLZ8DM6VNF/WvoLeUbin7+
SpKmDPapt3UnyWxW+LC4uY2T5BZXHxT9YVLKWtKGhsK1NZ7unJfTs9HikMBNl6C2
tX8pZgS9c89WTQegaKSxkWtjrR6aLZ1tlxwzbi6yu7lkiTOuV0fmYq+1bWC7iUU/
/BXTZwZ9FaFt/T8fdEw9PItXdBwyrgJdJn+9H+s1oEgQi3SAygAuvsusyxiBl6Hm
3WuJLNCA21ogMRaOp7sa6vQXUc7BWGbJrdkqpLi0dMvfbF0oTkucEI3qZV71CMXL
wbXuLXj6k6VU1G+PlpUfKF5CCSoZCHz5pZWs0tjj14dtL16osqSDecO5fCV3LVXU
ToES70p4GzPIwQby0MD40h+eud11w3ztRpyhkfmai2QjCH1gglc0Pak5b352Wgmz
D2UdJAbMA0NAm7QLttR9A5Uqlmj3zCpWSLipey9KUKH/HMzgYN26JUvQH9rnMrOJ
MctI8EUbkqS7RY9RfUziSk4HSoPCbL/bIzPlpdZ2JLmPoqX8dPtple8q2OUaMGhP
6FgSSkaz5KaVMZ7fTCjcozmePuthCpua/+JexWqAxHlexXL6yaGTnnCjifaYbsR5
WDdz0FdnocG9RSC2q7bfM6iswLCbLBz6FKAeNomlaibxTV7WRt/+zCDh9VmbWhsN
nBsE0zv7pXaNb/Pap5sG1QomhSG963UmlR3ymTHS7bh9PDJJZ2V9SXLQNquYPa4I
zjO/kRIEUjKqF7j8FAxbvUkv8x+M8iIAMFRw9bbdgQ7C7jXVPAt2EPcpcYIrK3Io
p2oUzbn+tudTKkxrwEh4LKhOHU+meftQ+LKUirsDkXq6xVPtPxLIZ4nf9+bcRRIQ
Xmn0AoswfPcqCuIXCh1N2Iz9Dbig28K+zXpn+3LbG8BLSvbocvrEwkLaAsIM2MBx
qsEQQ3oBSQEPUDkXJXZrsUN7SAK3opPAQ/yPyYb8FPpFnREt8e7MDiwtjXVVw6qB
Iz6vZ8wSjM+LBN70UWc/bKPoOAHi3sNb8KsaVZ7oHCX7LF9wUBs0GaEuzc+hlBZI
oAlLThDbrkg9nxZQBpUnDHtlq5iK7SvUvpCq7JYaYTxgH2nkdBWG67mVULyhp9YI
NPDKr9Xg2ETgXWBJzamdGDcRZjlYjKXulYIwfsTDX3cC5+mNGinag6jzxI+QCVm4
N/wIsE5EvirPisGhJUlhbRlvvZ2e/kNCP/pm42AoPXOIJR5s+NsjkaAQva2hBAJP
02pQKklPKt2ZpAhGSKR9o0cnJ3AZAgJ7VozcQ6Y8TfBlHkK0Gqm8hZ4+Mc9E99xk
+PCLwTvUHVr3btNufRx0qEdwlbAG8gW21Iq4GZnexi256282UD3AGddfkzwe5S4s
iGYVYiYfU6GubCPat0ctmEI9+loWwZrbQzQ32cuMhPzdPGxUlkDzGwhXycsALceH
KDs1mya/X77BHC5xb5fAhmb7oeixxdhtqwzC5c8O2KccCCw2mI2tGojYZmHLWgbZ
bguYkOx1pdENJMtSxEecNXPUzpRvdHWX5UNo415TbEqQq9jIzSvJkJFAwHbarooM
Qg5kLS2/JFReYkuEf8RMwklMcRTdi2gP07SAGKAGOfNYamQ3xsROsG8ga6AT3s1+
E36P3RODbYE5D5G7+AZ5YFQd8PV4a5XgqRQxXhbIsjEG8vaZ1A7tv0HbekrM26X6
H11h1/TWL15vFeJZKNOhJ8VWfFBVbaYgrhPX352FTlYx/bPb5PzfPEprm1DIXUtc
IwmWJqxyA/Kf8J9fLl4uvWfQVQ5U8b2xsHfub65TbbsiB7S8atbyzR4ic+znE4bZ
StGwPcJl9L+n5WVUkqZdVHp//q1sn15KPHWuyQYQuY7ipdIi8ACZ63xLXQxbgRpY
8OXhqFAXrgc2UAZoVEIZQhkWfvnz3tjnxprVzDjnUhrdXlsCinH+cQvXAUagRRb5
+EgFpfh+kFvet8tq6ZsqzA6dMNAwNDhR9bACPLkUR4/b2QcwzKtnAxhelbaovKlk
y2CUqUFDhuy8TGj/WEqHegHBvwng0bTRLF2Mr/Fr9h0b/qyGnLWdXFQ7dLrCNY+v
QhV8rSfkMcmN8RbbSv7psz9DwY7M/UQXiWYmDldlZzbfAoYmgDUYCgsfeSP44gpP
FEuDkoKNa49qphesHpjlJJAYQSQ/szd7JarJik/oC1xkTqDN88mlbOzcef3GmGYS
HZYcLvrxsL+OHfofGYiApX1kylK3MPxfAhue6GT9/ycwf2GVxcswi7cANXmdlIsq
QQPhIR/C8u2j4ImQgRYB9TJEZTo85dyqjDQjolLB9kGl7kpeSlKZdlac1U0QVL2c
ea6O6lNvkDSZF8EhG8C7gm+SxX6mDoHkZ+vUhIn/IqjJ6JvBqerzY49DU6DmsWwf
SWUsfrahY5FkVMnbCoed2LH4G+hRYBPT8WC/kZ9FokThT6RuwWyF9YQVtjNHp3Zh
ZGY0rlUO37+Tu1zHhndtB5/11qU9p3PZ+mG0nPcxWfLsWNojwaVeAuZ9nm+N/+OP
lgJdAnhPQ9PPdJ7CNdjO4FX0+AYqQUdGhy2gLXv1nSFJynOUgqtSwpO1uqxSNQDM
+s4o/OXeIdOr2/NKkhE+8TBZ8oMrWtXky1V1Kc/TLDto2Bf8GSzKRZELPI7cqBBX
+GdfnFAWTu8RZm2U21av7SxmghcCEsjrHhmnDJeTZSINYWDOylwQWpYvnfODwP0h
HazRYQJDxEtVc6iU25VhstTkIKIBKCk0GzmQoofmBFW/LK/4CF1AdES1L30Esi8y
MrRNk8fi6Bxj98mzCW05iiGM+tOBxC0XGEgx0BWmF6MNNRmPz2RJKBIH46ur+a5I
mN/lHMTXRwPtQPubHku67uXgKVv2ksdy8ozMIIiMaV9KK4NEEVj4TFMrpQrt6Vgh
hDpah/9qkjMH1FsfYMjAtnWEM6qHxfKPobt+Yfo+o4V4TdW9wTIPeGmMohhF9sIu
yhw+lfZhRSl9YFp/ZmIh47ROCJtCFZvEmSWhJGVaJqGsITKpBc1n1v2DQP2wA8pv
/bsfgFvgKIajO4gX3X3ik8D9MCuRugMUKt8Xdfyjc6j7DALziPBE0SwtoosaJG3i
CKxYf1HpSwJMQTuKd9X/WJ5FO2I0GZ4YHa0WxXIM1897ld0u8iopRo1lYwQvPVjP
qdh3iXquDTd7XRiSiRnddHrulfE+6cuWvV7bTU+p/MZ+yzIExxMmuv41VUjYnVJm
jzFD+9mZGVElFcIayt5R/ow6gHIevt3hGKbpDaPjrMlmNEiH3zXlWmqOJ63NwK1k
LzOo6hSc7GC43tF4xNElhIIH7DPqNSjetRzpA/J5bH1i75bjLuQ0Yh8/wX3zJWtR
rOKFq+VWtqLOhy+yBHRv4QQWRRbMIhEp0/9BFNYGMXqPB9JEuq993/HvrewEaQA5
h2UxRuqqj/knqHMh8WD+oq1vfm1X/p6OmdssSbcwi0qYT0jN7yjrqD17o0DZVSEN
joxcLX73UjVtxy0YbdyhNwZz7nwMXjQn17l+MDNov6yFbLX2HzpWGqNhelaB95Q9
rZYxCr1c5MNEOcuOn+spce78FQedXgyLjK0JdQ2A2/bIHK/Dav/fg5F1sUPO6Z6N
wtd6RVw0XNGkpw3ddNQpqxAnQvOZzvtWUjFAsfRd88Lv3BiA5pUSgZajcb42Arqn
vwIAzZ3ZO5UadGS8Zk2p5nWhwKrArkgQgNbiGX4NDj7FwLUsz0W9acJj6ErfwKgQ
fQGPpbNoOtItqTe+AxAotY8zCb+75gX6OsJ6uIfZrLTDcclpRc2eFBVm/nIZsNz5
BDwx4oIg9MVNQhIKrry4rZWcMaHE1LPkkCf44KHxF+mvomHcRT96V6XI+CKpU+IX
8OMh88Yn+uk6ePnfQVLSvSEWS5oF4aireKDXcI3cfrLKrdU/s1+lYfdGTTwVfByA
K0kIolZvEpZ/6fTLB7QNjw6xwnYugUes2UpX/HLNJcrGCcNCQajCrGOcF3A7BGO5
nBWKJTh5gCW0Rtx8nNTFhsT22VYd8x7USHYifHUGb4mHcbfD7GOzAKyN+3Q8/Jfs
WBuwQnadyVSK64jWUP9/1joLHCzPnid+4/fHx2a2bO0BtOIUINXOqWBFpRVOjPjw
SD9srKZ2Vc9cTvHlj1T0BbjWZIqBUMyLpjJ4C2PLIjDiV8nkBJnLZOot75bSzidK
L9NfGrfTuGM8Cc45M5BzvmCIcIgjRuSA5kda80aiVZq56IVhB4u1f8vlliKV9v4s
IUn9i1uam35G2Jg5rsKKHRF9SCkskL+5cRWK5nE2sF5UZwH+FV5UVvDmJS+y2YwI
lxSCBZE9Dgxkx5JlW7vkHUa/P0oKdGhfGokiGm5y6CcRS+N+uAYNTCKFSFefXXZq
rvklsEorAmsVwD/5l0Kpzsi9d6p0vWU01fN6MeuAbhLJfJUMWimuBoQFmXLFKvUw
hxxhvB6AlLsGLzY4sv5Sb1a73it8JAEi02XM0sIwVSGAzJ+qaQjlGD5ram5W4JbJ
QM+hdBuzjYtbX+qqbS+GZYHJd6KPBVFa61ZIRleJFlFgI62GUllZrJS3XughFH2u
mnTU9L3xNGOM/ac3GAMUFHThVVI1FfEdAowQKp2fXYcvbWqXjWKqKwIYd3qVYe17
W4ekke0NRVYRYYhmzO1Z+oxoPhoLVgO7dvuiQKADGXkiUAxs0uIfxVjM/i5kqU3x
/RtfkVNSm/1BWZeLc0jEd/QvnpOzoJffYj+V77XcRNM20aibbMMUf998ouFkpA4q
suFripPXt+aYYl27ug5Kj4soKYGVulsYuFy4neSNOUsajS0HLZpIVMwkO/Qo8YY/
alUTuBJTfSZA8i6H1X1n+4icF8Kx9x3VUabPOd8rIMhz6+xwQtWkjpjkMIc5nwj7
4jqBDKuAbv45oYiDtADoM/XkodorQTf/6ZLVRB5B1QijD/og/Mp4vaUVk2q2EkkH
CUgGQJXoMuusq0lstjo90wThVO1dVi+y85eXeHxJCnfc1LkAtdeznu8dYDAKEv3G
kB+kY0MSFlP6t0qydzGLgTyMGNolcabgVkAAKMSJ9VFyvQciUkTmbbD9kH3mUURQ
+Am4R6Rrhh8wWKLPlIlQGRiojqZXgJYM62ZRs+KVcvtq87ATXdso25Pl9rAmXSrZ
qhrW1yVO297rh1k3tIYISBsq+cVLFR+OW2v29684/IZ+dMd+tqerhIgOmd43XnFO
HQybnHLzlY4Dbv6EHb22Tzx8M1mNQQFwUMLhdsW/kz3v1HWo1dph6F5+CqkhryzW
PbG1vHnEcIa1sRsDUHpVlT8XEQYW+HuR2Ha4k2NtFvx1rRx9cVX7vOIYaTFr1jPX
jgYPrrr9TnlCvFfrUpinRaQHt/soBGbQCQgZ0HZQx9/KtTiXQe9bx3M5oGbHYmxV
d7DxMJ2kdqR/hy9Alyh99ZjsvoayfBE9rEQXBNSMxKpl4b8k/KoO42ETxK58hNGY
ZgeF3JGpXz9jbD/qS8vd5ay2HlKiHktLcig3cz5Rut75X2VaOfIoMo+Ur/bzvudJ
+W8B2EGUshU7rDS5ZBU5ntD4LJe6wqxve6fWzO4oK9nLF4jpVFPRooIZ7RzCIHvk
/jr8uk8ujoKI6fEKinZV0bBNOPP2OlTjyT298wQr6e6E0mwl1368p6Retma3ifTp
ylBa+GH9jHXlQnNTRIyyYr7WEPwYQhXvSBZIfWhGI6CggXYwQZAWDbnlpi/ASGBf
RTi2geKSe0QQqcvBRJqamT/1CX1CPUGSINjHP6929J9TIzVKym+XXgxdrfREMErk
KgIuioETTz7gRooDa37oCQosEUsHjhLh59VAhGl3RCYFokPqT5oVETv/xqjEc5Ez
gIcoGd0MhuOh9OYPMlO+WxIREJcM78+eH6r+ZGaq7px4rVfmouG58mkA7JOD8ch5
uKgER7ns9HsolivF0grv60Y+ay02zUL9kXtmtAKDAWg442RTlUSvlVrjl6S6tJzJ
P8Kp9HbyxpWl86hnOETX2fdyAitI2Wrc/d6p0nKdaaqNfcQZc/FKUa1K61I1z3pq
+KzyQBCZ0zr5F6gcetYFkgqQZQzp4u+TBElpSqZsyrkDO/DWwkasFDCuOAzusVx/
XGtWBnUnZLeRMBGIpTQunpid6fQgpGzRO/FPj7hgxL4jE/1nhnbRLKdCPu8X2v5u
BFgcwdJfexbutVlJw7/CusNUdi8RGM4hQXhhMporDc70sHwvdVgM3jE538TdK1xr
1hQT9D47dkjuuwFSxOXOmI1M1JpI2MJPVM6OnFcubEAsOn6NDeoFR/+C/RE5a0dm
LVhOeo703a+e+MdjfThY5veMv2qJJDRoSKOpw2dh7uPkj4UYN3XPMlUrNqmsIyFh
HypQWAS1dkkEHVIDIUSuBntxlrLvVYo302trUbYHmPy3XrtfpEZtByVya2u8kUZj
IJWkIAlSbB9/MzX0EOT7djhGsVNXN40ZyvhF3Kq2LuutoSbSwEwOHRCpjJyRIiBo
HCOZ8Lm8YzLSyNj/3qahwxaUMN6jqFYHDyF++XREzVUrTLfT4TUWHBdTr9da6hCO
MQEknL73zSmRUEPuTxXbyl4fWCDxIcjqtDSxREoPJU4soSinJjOiKhKu8kzZD7J1
F27BQJDQKdVEnfBPtOdaD44zwT75gEMIDwgx/IkYpP3GLx9/a/8A2ffE55X+3EFa
ovNrb8QGZl3FFSP1UpHl+/YlqPYcUSZjvCb/ussrxOckmAnb/ngTrkPIvgaT51bH
j0mb8Sp5HpCQBiz2PCamUjxfbnnDvI6Yj3kTIhkonJrhke6eA0oyC3HHEpcrwNSu
u/2sjExwiBljwyLDHtCKc9Maf1YXik3uDTiNpsZ2Qk4fd1bHHS04FSAJt/u2gTD4
jeYzd8NTni9TD/2PFE7xiJJCmmbAzWDlCa+J5onh+CLgOJbY7S9a5QhrPGkUvjvX
XdZxNPHBv32LuYKSW/9xOac2F6Mqt2T9LT4eeZypfJpuFSnqmHb0Krmbp10/6GvI
pbKT07lpnIBV19siUdVE41vMMw83ZMlPsYGDFO0fQbwgt/VTiyE9ixXaAIuxjsXq
FqUzWN4l8hcyfxZo2KgtpUoa13qIKi/eeyKu8ZdUSuXm1qaPIfgv/nPSbQ6151E7
QbkNAUzyZAPybeBOx4RNnX4BszWMJEnLZGXXRsJF7EBidlfHUf/5SGzLgj+qsy8Z
loV3ytro3TxYKARysU6kgxzmvd0gyL/zwhupqGnoRwSQ/iEEGUzuN/uiSYhZDTLi
eBe4LuaDJjNK8yMVNDTzF6xhfXlebSl6eh0n7Fl3e13DF6sRIITnY0GvWPbxbdNh
MK/6QsjXLOhYdX2cpWQq/AfrGmWXC13aT7GRTFB6UeEWlY1jBAZAOyzLmOnvFAyt
1Tu3+13XlvgowHuF+Vtm4PMuts988Q6bTCIvSuEQcBc/vpwjf6oY6iZU602hy2ca
pbx/lhNgeuuTlnXAq8Kl0VN9XPrJ/UgxjMtKeDp1JF0XngI+n3Hmx6Y5TxNvf14e
GWf1srv69lixyLPlaJ6++WwwMbxTcZU5XbrLdIaCSJT7QRJbazmwTe8V9C9/oOu9
FqHsZGcxDHqhOHUPyGSni16gNCJ+b+YOsKndVkpB0x6GWs/Ld4fPFIV4XWVWM97a
sVdSEr0pTidAHIcst159egfhpkSjc2pDgUL5vwqrPsYVyW8w/rGkyGpQ2eyVvtsa
rHwB7/F7PA4WGl59IAOu72JdSAUsUSFv0KobFgw56PqxQcRsYvC03ajeEVlmyq3H
NYOz1r22ji+H2CQxMsqBCGRFLq+eq9WsEMWqw92kAInIkv24VK7iEkkvJuKIldcI
1HglFGUZw7gBmYLPBYf3wX5Ff1CMIR28OeL3TGD+gh9jcJQpN/0D3ztOYJGdMo0L
Gt8mRLaN5eWuHSgz5FQoo3qrQxHMHEQlRhYVw62zZ5gAtQS9d9hydULUce+N+SU7
2Z9mBqtFFPUTWun3HjgFBxBboBtoTetfXlofq6Zdgr1OLS4naE5TSRuCb0DeyUu6
a1PkWL9ZZ+DrVQx9wWTU2kInKJGFcoVA/M+IrqmYiqh5jkIb5+KbJWZL7Sstxscy
qLZW4LNTqSXkPzcvMWYP2KB5bZkO5xgwFZHFmxM3xYz66b14EO3zCc02+RuaeT15
SzR2mqH86Eax2qL9OubSnExgFqQAYwNLfVQJHB5dqDc8qgAs7x02HG9200dy1pO+
oPVoxFUXosT8gG1RAZ9HIKPUtIoCKmgy8ublF3MFFiSDOVMBdaj0TfuJFRnEk7De
iSPG7vDvcd/EPbp2Kl0a5JrhVnLD7o97EgtN5RS5U3v6cnOZXUFu+GvRZ9DkAgz0
YixpyRjPBqz/hBYkLNPFIDAtABakZ3jZ8MNYkKEeVciX3xAZMPQKWfqxpyUhjhrg
cSYbyDvTEMNa185ZOjOnVivT9smHt+TGWuZpeugq7Iwwb+oslCj+XCru4w0p8BNE
Dla9RWYycizATeVClW4zWV/zOyMLucCzURf/p8n0z3MkB/l+RGi/xsIj/AaAu7+n
4FFPW3g8pP6AYwR05mM29KZTbBEarz6eWxtHxH9QpMmQAbttukSAvtiUUhc3LZce
zTPzQoofRa4TKyaNf8u5BL1HwV+eHY1bU2a3EsG1kIcM2c7VheqfXcR/r5LdDhsl
is1HzQkj7BOpJfF3z6ULoRKc/koN3cnYP8zOe+oQe5W+3/Ii76l81fbYZrsyAjh/
2465hh1CGPyEzFcRakoWuilgfoO6AzZ+lApR9XBwhds51CmDPCwe0fIZpl6CmHfE
qnwzYaKOheUdes9uvV1hvMvBO9TFujx3FGdTWq1OXDRIwxKT2DYkOq0lJimGrh+s
ge3iNprVVeoKoUHXfCpISsHoh1OHRPDKhz0FqEZjJAZqc5nyCYbK9U0JmE70LNhQ
vW3YXfGtxSvNP8a0YnH4zd65TfD9CFSoogdRnIYF3p0AJvwG4/CPGZQU67zh/HNU
PQAVKPM50RdvT1KqL3rKAFDSQf7AF27CaNxeH34RBRvMl88xIUL9paKF7RPmIp+C
fPsfkK1QK8W1NLlTUuaKZE/tBGQw4401jZoI2d2eHp/ZFvKmviFVvIc+i7hIihD/
zc+E8tP4bYEaRYbV3UuQGkBhlmFCYRyzRE6dHUZd5Hg3TGXzl6e3IEA0VhOjsULZ
soBGtORLVsJfeF7WTJcryxnoRAwRvEYOlPWmGEyoyxya5RsH0MaLP2z1qbllD8Rl
WIkkYy87Wh8ue23VXI71Pgt1izSeUlkL4fRapo3F36xT+s43c2hgHBUUs4d4BAmU
9XIRfR6iUc5/a2ZX0wA1uBixdQhFajEZ4fiCq74AhqUbroc7xKDCCtwMHvfAY5t1
DMb2wJXiUs5VW0lQrU4HPm6dY1oz4ZVORL/ntsCVh1BKO+IuHNc2uFuZudLWqZFW
sYUtvDJ75MEpe+iRtOAeq8MuQTt11nXDEKIwmUl0O8zigoOwTc7dTv1HhXi2dPej
W0xWKMIPLeQPBrMP5iM2LWC4tbyLQPJTMPKBF8k4rfS6Fa3qwVPc5yAIisqTaCSw
qW2ZBGhXc7gbv6KQo0mLSLA4A8Tl5RKW2rWVGw5Vwco1A0bzDTZ7FdF8n4bNfDUQ
WtnZpT0vQZKx8QwU++Kx9PCkiXN32WBVdzllhX3DUL+lqjMrmaujA/QEbOJk3ild
9n+pAbDe36qa3+FWMKCvtwkDcC7QVrRziO2kJ1oGKJGN9zwCIGqSghZvQCooCjfz
3Cw36QqtgqrJc3OFbASQ0t73xGW5o1/kevsw+F6DUtsWXJ0+i/K2QfJ2Vwawo+LA
rDFoY9ijS4/e33Aoin/lClV+zFTiO++Y5I4EpAJRdOwXic+iPFUTpV92XmmlWiNO
WhzqIVCLOxKdQKaRkI7BYzK4Nh+PZbQ1YC23k2QGj8bO9RjHHKUMFEkO6lulqb/g
ly8G3YzovDwoVmwRngBQnslbQ3QS4bo6G4RD6x8Sy9MYkIFQAN8rmF+1qzZTa9cq
0OiN/XqddrgkQwiJU9Vi5zHUoVm5Tb+8USCDj2mjOORzsmab3GPJk81hNdiZjLK+
tsuw5IfbxJNTKDUZU7fKqtdfgqpVuP1al33rQa7flu9lieSIoobt21jBHa3V5zZT
jK8d+kptp9xXT3lvynbhNP1PrKPrc6AanaeHZGw0VB/c6NPyAsJzgZ16TPzjV6ER
I9TmTx3xgKwkWTxHXyGw2+27ooOkNs04wwObXz44OPXTCmyrQGgM+1DRI+RHdE1T
9wj9veyRG4/O9fsKoCpV8Eo2FnVmD7I6K4yOof+BPf588P0sNMtjUm8G3ynAtg1S
K5S2XE50VE2ywHZX+wClRqhyHhkohXhlB4C0gGHTsM0T6/z+CT9zhNSc18VB8YtK
LUUVtk2F5c9uHUCIj+GHVTdGELShDUHDbeFADe1pndEzKEmslajlgNj7+6pnD8DZ
IMc6cup0IdLUCN40hJujsbLGCWqptDJuyvwK7UIogKcjU6F9XYrhfrGC2sW7tGLR
/Rs/poZJWCPxn5x2Qg4GyDjkK50kBOzVWHp9rvgQLSrcdBaV7RpiM5VhOm3IyYoe
51GbTs6Bg/1gRJufHyaeDOQo6bKYV4fEqvSLuucYqBwxj773Kvd2wzixD54QT8S9
U20t2JisKhnzJYhqRxqRg1lWQDpldIbpkFkDOrIqBI6B4Hje4Djs/gTbrcDtLtE4
YqZGyP6c00LHRuW+hKID1FrNds74hh7EP6pVqRKFRNU3K4TEgujsW3AcNQB2h27j
6B2VJoaBctgsZN20iujDKOk4Gb6vo4oVbzaVw1A/ICpUw9M8Fut2q+tM/fQAOLg8
OY+iKrgYJIQBXZCx4PAsaDvrpFznmYLk2nq0+AZyzlug7OX21EOjzw5VXdWpzA/J
mEuefdtwozQKPUGR5XXJuyUZVbH1Zoo6C9v3YWyPZCgq/nGDkeWoLlxdDBbfvkrp
E8SYt5fRRRos7D2vcOoGVuW83Dbzako7IJ+p1u4YtjAvU6K7HWxzLq/Zde0Bh1tP
lE5RflUeaywDgeKWf/TDoC23ARlRwuDNgkMogg/g0vA/9CMqYdzvvg4P6c1RtIDO
YLA9DYDeCicHEk1MpZQMGBkN1DGYAVTCX+jQQgi8jyzJUq408JVQhag+DrefLslF
kOc72HCpCT3TiIRgse+xTtAyJ82y4bM5OyRE20F4VUWzsoPi9AcxMJGYmGNWnQZz
vfXWF2hWXkKVdJmTurBoLiOcNHgPfEgVBWl/7EAmhGoFX8O50o0Da7a6hHusZv1N
fFl0kFtS76qzI7zPAYh3J5WuLoTBujV65u/Nn8K8f/AR1oA7UVcNxKjaw1YsbHHn
q6cmEKS9CWKAvZZBHdQFDYbIkh+VoH5UXcpMHht2AYtkMZYsuwuatqdF/m+juPVy
tNtClYYKQ71aVsrCZK1x24XwYc9vOVCOou7eCzYwAN/xiO5NPQq60HQxWxkFoEGB
I2YFnq231WikVmOHgMUZNUl7aDacFE1fZWPtxag109u5xVpfuoW0dRmBVi8ZmAZP
3+j1b+7beZbvp4LRCuj3U8oN21253sS3FAeP6uOokiiRyN6lRbITTBf5N9we6fAI
qEBXrklJ5NCLothpIXCreLtrGM41LuOqrC2SCM6q0/JsfmKRp01exk/yqsGrvK6K
w21GwOd0wFU3GEJNPYi6LoprFkjTuvcyAdmC+ZCVt9twwilGECkQakShH02WyY/H
TeAz/6UqJ/7k59DO6Sjvdt7BMOgZ8jiOWuz+NnCHpjcvpYsjHYP2fsjMYMsldNuV
wgMHqK/i0qTPSS+SseYk3daRyklvathQ8SBnvK5AuGgwQUatY22GlQ7BN5odyXem
tChcbecYmZ1RjGnL1Em7jVqWXNJNKkWjK7v+D5zHU8ZXq/IVJQBsuvqyKrHSyrq1
1UMv9pQII7wgu98Xa23h8cq6BpK68eBK+FvE45NdG3vRHTxOl5NnTw9lqplcEPhb
ipb9KTHk+fdZ8amPS6zRxOVUe+Ghkb/SGKavaUImaNNUNEpZGsCJTwQSAP964si3
1h/O0GttUEY+pQjxMTafa7Y2WW3DcNlOuDR+qucc8wYSk4x1ZNB/rtfbG/BeUsHT
8k0qalOmfcQQo1JdQA7gUvy/THXOGxEkLmafdvzmb0ek2prb+nmT5Yvu5J0XA924
wSTzAyPMKKnTaYd6TGd0UTRXISi4Y9KbQOdi6j3j8BFZftOvFOcuJtAOCW73KkT0
ElUe9eTARx7XUeth2fnUtvxIGQDGiQ5/rT7/dZCWuzLCytTyi9FhGqij6hI6hC/A
542nWMfrUWBxybwZs8+R57y9X4Nt1csYQruj+xhebx8rEke9d2WTQGzosTTQ5fuJ
s6x4k2whlIPh1g1rEU6vW1hhVoxigSIh4BY8ECqEKL2IC0n+Gr0v7ISoRFu23mVP
GwlszX4bHcWwOQSuXPms1fZnTZjE4WzOlL6p59ebUMLmkU3lfKP/dgxfGBCPDUJU
tGjtNCKZCZXwGtiVjsVy7K8EGuILdlWPVix1DefIzYBh0gT4xPrD4iLY1MuNiWcp
4XPiz0QKh/gLFmeM28eV1WEBf34kWfCcr7Ht4ipAJ+OTTr5WHHIoX1iA5I5//pkW
zHOr9d85rq4ERHsAcpQwBlKEd/T58NSJTlXOztP9dVPww4QhqJjIOyM4ZKFG/xD/
MybBBkveQOjGK2yi8EvofYXMBsD6xL+QamDQZLWsDpN80Dg3BffRICSFEWHaHJsf
lfrMLt+QA8cZSAPh/w/oZ1LZ+SqYLoiNiQTVwBkd9JmzAR5vWfKrOjfnyJpDEVnD
2lXRTkUWJIe8QBWSRS/SkJb4z1Gk8lSY1KFUYhtM5eWZ6fzfCiWHIpttGvQuTQym
0r+p6ik3Gsnguck3221Gxu5wmXS2kFvsK6nJbL5yWO90EmIfaPaIGPNUT03JCusn
mjtMIOMHssa97fN2f1376pdOOSA42b2LwdaQHAhTePngSjPBn5iIo7fGkZYuxfq0
OUebjVo4F9/9CiLeU5JvcMsodWTIPcCIH0myESQ6oeegIPp6wkTtJo5hm2c+jnmN
fBgflWEc+qjVBwDnP0UBkzOQ8IJe2mqsS1+ACTNw35ysisDd0DcCZPsIgS7qkn1p
AsIdX3e/eep1fIMkKqRcS2QRW8sbuD/2ZYSDR7ScVbdBY31Z3nmNZfYHFdR5Q4da
9jZVJZ/11U9ah9GAzuSjTLstIyfrhxy/xoylsLdFIlyffhoR2ZnIqPpbwk8y/z7A
c2pSYBRIkO8zaMyUS47UBNGtu5XTYOvpuDxZTRtx4UWV53j834U9ogsy09rQG+yI
40CX6otxIl3QTmitqJYlxpgQv/DxiBtSnqqPTFeh2tAFYZdQv2edt4BJGOWy92cj
FQeqqHbXoNy9lrBpKyoIFN/GbbJkwHaEvhJ93ZkW5Irf/XEloqeeI0z3nUs/dLje
sKnpvVunRRMdBbEDO8x07ynZtJWDid7I3srmGkYyYvn9zYMUKNCUlCozXEApGJgL
/75qX/RQILrDTjPXZUk2OEZpioqhyHv6w2BwKcev32orea6pWBFcpKnqgSNqjxba
oJLtyLrkh2cv1mdc5oE8v8eM95PPZgZJ70IVlbCh9sn08jQhEuVAG6iuGf9cG1FP
ITn3b/UThmTXFK0fVXLI1HIAAAZaCgOKwdAdS3jugwuGTelPET/hIcGrCntpCzqi
Ta9VQHv2SpbbhbdQ3bQrGW2Tu0jrJLTiuT4davpwyDOdHRaycndlq9qBFjhzkXEV
/qmbrn7XayrdIOuvPADoz6RU8LXHfTTEBMN/MD+5hpwGtpexQUC9cBe5Fin+/l3W
CoA8j+Mo7HL5YPbwZmZJzWCBfxcJdhim9a1jtmSyEIpnM9rqveeyNjzb6U+fQSzu
xEp9UMsLRvjIFK1AmaquacHUa0NAl4Yid/J04x2KNAZSvkN+OdocqKP+wmiui4jf
W2KtKKzuVyqd1KFuJm4cWCYIcDvJzrJbvOWUUekN4GmdtZ5teoNp84t8rAuJ8FjV
T1ObsDYArUWkYluIcb3oxtRnXXi/DtuU/ksopQK3VdLQ1BU1zP1CcmgAPsS4OUxb
v8xnfo9vXFOfNcOL27X6oCPAJox5tIBU7hfgiYEUX+9r98cQ0KZFZCARJS30A9ft
m3Ggvgapb3S5pJzd9TXm070AVJpuw0KpJoLc4s83+LzuXDhdFfyxGAVcn3Yf0hwp
rcn3GjpaRpT8FrJPBRMgMYViNkDwwUA2rUhWFhqXKnKCdygWy7gJMuUne5GFp4p7
jqWQ2JUEAC8HrQy6JwSNZJgp6697w10cod/NR6lsZGj4qDZtIQDWBbx9zrlIsXp9
y0C6ziOOlGsfhg3biwX6w320SvgICl7LXJG9aitKOL+/wVUIZR90cGS9BK7jL0CP
W1zbLagMQqfUgAXL+Dqj9TvoMGpfc4fISokEc7an/fgP/FyPzVomt+zB276VBpXd
/f9/gCYYLm47sArEPtE9p2x5XSn6cz4KsaHHqZ2a3S9FWVOZU3vk8Y5hzAH+k2XZ
RBsUN3AO4ypLMkMZsNE92HZtCvOCoHSWUMDc/zDSvUD4/KVcgXhYvrv4WhU6GXiG
QDHOU6IgrnxEMnYR2mBbikhKLw6kjT5MBPf07UCHwLESMnXE77WYQhIoKSX2W6GR
XqxXxUeQ9MZfmTkwq2x1oXpsVnl1B4GBw80stAVv7luEVCpNKsdqy2qcEaOEoC7r
+wTXLzVI4N25OWEB5SYlj4WoAGEm2yoc3EgaTCYsbNMURHn7T4h1BACDmkQjmtkm
/fTsg6ecUGfYjv5Jx+4Oe/oEHj1JczkH1a8GaH3XPRnCyRKY3xlJFETkm8qY4DFZ
rlWroAlez+WzxTgDtJkhg/uQCJILhP4v07vQ31KA3c4cFsZxDUZ/xEOI0jQMzhBu
oB1uZ42EEN3HATeH8YzfOQ1NLr+/ZocBM2czbkOmpnKO3B3TBG4cnhCUadzy3dRd
KCUalC8SFMcymECrg6RMWKl4299jjgfnhFJJFxFAfgfcaKQdOV3Jyqc4uI0tTXbV
7Pyf22FGVc8kqzvntvhKIst9+wMfOdzmUSAzfzfnxUrEOMHclAYKlapQG3GLP9Cf
8lh6Y6dR72o6oR19PFQL3l6B6Fz+lejFg5rjCZvkrEaMvm5xkoeNAeNasMV6UugK
NhmhYzThhLVeP5USHzkQY/rXSWDSLZMKaUKHCymXCwN4QcWg/aCZk6myaQW6vYeD
ZbH872N3DU5QFifngrl2UKkLbARpbfChF8HlBYT7UQVi0zTnnXXcBnfqw7bRivjb
sHWRSFgMzdgMG6mfx5cBLin58l9QBb62E+w/ujeoQq259uPMnH9pYT5uzppVEy6l
HfsJbJb+RTBT1Ga7p4pN0tJ5Pq3Qs6eJAZBsJQmeZGLcVTE7DbCqTTzJQ4wvZeJ5
ss2Xje9u7rKNIet2espzLhzcRCDoo4BiHwkXPtarmnxbrsvi26fC8tSW/w687mEJ
mrd2a/3MKQK9aZrAjmrsGF9vJ9u7OKTyPCFKRNb3IT5h4bS1jMzrf2T3MvJlMnqH
K+Wf6MeCJ7+agncbXEQotVSkyEdJIn1QDLrYNXl30ffuLpxQBABXYd1hQt03MAsI
UX7GJQteMh3vOeClt1Cf2UeWaGC/cVHvDdzk//wKY25oTjlmWRwewvunBTdInLqj
6vPymgtD5uej6ji1P9rfFaqlzLuH5BfL/PtMKiHmbThx0mUXgeyPCVYNRu4Yi5wM
RDTqD8qaoEK584tYCiBdfWxLmfhrodANPYY7z7xntX9HEFJYpoDPFza8Rr7x5Zt6
lCc6cbuBgXaXbB6vwfdduyb4tX80o8abz4/Wa8ARx5+J2nWbLOI91dw8OoDgekTk
CjQ2LEvFy0eGus0mWXIgaLxYJX4tNpCDFJCvPlY2ZqP9jeiwS+WiG4+Cy74WxwoJ
E2rCv+e6pkKh0gSkBytvUFKuNX2Q8+XZUgvoIjdTZTPFRGhaYJK/7bnkMTlmtgyg
VggWhur57/O1PS1qGyXOQOfN2GdUgjabf42BA4qXYEWh2xAqHRETofq34LMbDdyA
NZnMbZ/8CUdMRl0o7S+d+kHANPitWYbt6vF0UQwhyuG9MvTKhzrGK/Nb4N3rQdng
tCoe/fYc4bV53euetUo4ZpKp9DmQEqN1U/Ef48epuiLHGAMhgqYU6LM4s28syt9Y
t/1LUp0MOhDqpaToosUGRkZafZ6Z/xpuuUZjgCpmYyiKD19VN4ueONYC5cOR+bsU
Zn3U9O9ZFUJhF0BvNln6q0okMHiIoVBkneTVeFdqTsRv8X+IEPLXhr8Jzh2Q0Mb4
99jNnqRRUAP45oAVAOzmVrqy+2C+Hs6zU9av/66Nu1c8rk7duKstcQBOqGO5c8eA
Js3C39KJzzb5P7BUhCB68iR5jO+jU8fgdPjUKkVGCRIL+6ZTJPBPirZkUfbAwgnQ
SsVGWDdqYssxZjZ4AOEdMUEFAOSR9uRbYyXF2MEupdc88hCrFwXroWYWCQsSfRJi
yEFw2N1Uh3LNHPMt3y3TqPze1CKXYIcNeLqekGDmIzVs+OcqbqyN9y3RXE88n/d8
Wqa5aSUo3O1d+3CHL26SBFqn+7CpoIf8B5qHBQ2wwfShVtmE8830rWwXXV1ri+TV
GRvUSZayKWpt1Nw62EiMb50cWnHLhtK5POabQ1Pp4sa2h4chvOdYEmzG82yvZmFH
JOmKkvXA89oNgneb4a6uu+j+dphSIUIHFXDD7S7jdD/9hzs6PFZd2d5QcmX1FXvE
sBuReW2g7o0u6M0r1T5Xu93yn2YWVCfyjtuf65iLIg71WR5R7gqGqnCJMXOCx+iU
CeUIuWR7MmmIl0d2CLZyGggQPZ6ti5If8hZrPOgp7GAZqGKZxhuuJTyqO8jpwUhJ
UYEx4XmgbrF64lY2IeaJBUNiKGWoKmqZqO1eamwjETG+VNwEs9p41FmwuLrVKCCW
EGnshLV0By9FCHM4yTnM5bvTUzly71ICeXuplMFALf3QGP7IjWlt+Qy1oIvp1u7q
PjnyAscTh4bmf0gluPlxd8/3Ebj6xJV/8Un3DQaOVQRSa5FVu/FfDQzyYY1X0/YT
vRuWUdwneYL9+n2KeOMgZKc6ppUBMR0x/olHf36iRWMvjMZHFKE2QhdfjKuc9xfM
qzAMtSayDtKB0X0AlDPA0KWYejagm617IhB/SIjEYOiBhcX3zpmj+2UA62fJieKJ
TDg2NYE5eiuR/Yqa8dK8ez3cRWFfSIXbFFmLbgflgIoEFqTl3sBBvOPbQBLLLRKx
8OITZPZ75/4iMddz81HGjG2hwdGnQHn9ET2ug7X7nDtYa1PTMoHH2aRSwrLxLMUI
p86oOL5pVJN0sCgQ31eIzsV+U/zA7gYk5YjaHYvJmjLKN7AqKVzhun7Oz3EcFOhU
Tftma7is3JwhJvRAfilzMuxdVjetx0/Xnfx2X3lTZd5uz6yKXrLscHPlsQ+THjNR
oSpOk5KNCVzNn4UfPnUtodxr5hZrGH4xmvXP4n1n2lloju93qBWd2D9nPN71cQV+
L71msuSQjUaVDgsvSTM77xYYk7wbQlWqatc3SrvpKQXpk9Lvat3A3D2HlFk3q+ND
+DTYCWfTKaTVruHXTwnyDLKMnO5nSuyCS6DJTsjd5fAsg3pY3bl8FSjuXdqDaydC
AN36BJ/pMzVUzbot/ssvTVMH1KFubvtEIFtelw2qYITBVNy3vbfNHsjILu8vSdTV
zGm57GPHiz3zXhsaVa1PWQiyKZUZAR5C6Q3VQJbA5ACY8R8XwTh2RwRGGFXrd4Ph
inRnWR033EWW6qnAo1RY9ZZIR5PnBgMSkOHnlelPFb714BOGwP7OwCifOgi41EHg
TPolM8rpShpLZv1h4eLPkQDQj9shD3GltBpjTvJ0v/3wEqwh75xdcoVoaX3zI6ka
V4rPvxtIJB+ENkrjxlfpKLH2jraeswJM9l9NaISkdzFynnWkRdNz1MYVMJs8OE17
b7j0BrxVfCjXqAWrRB2trRIBNBKRavGrbFVsK3mdT4mf+CdZniIwEPPUZZsh+ABF
KsY/k57kdWTWOoB7KnpKxxNbMdY3s1z3a/KTiFcVy3CxOu2ASmvFRFQ0ZfF68Wge
ppzMuDacLt9lYsEgeNd6fkDKVCnEUEZUciVupUkY1/MKIlqwIbAhoLUEP/WFKKSf
ptHYiybhgEG9TTBNgoFtJfSs1FYfONE9yCTpg9Kgcf/87UIx6ZFuls+pgSXZ3P9U
GJ9D5BKZztWJIWoYsbLhXRppI8Kn3ozuaVxyZSZhgJEYXA9DYTW4wpAw5wKMYRmP
ozIA96aZmvEl4NeNorJJtqbOiqIxjMzRAFZZTk1UIxq3eWpi0w/uDEOE6wx0r2s9
X3bOWeMVNkqhgY122lmvQPgBlU/YWPi5rCxxQf1u9r2bXpYXAgpRMLuz7CoMCS2K
0RUQx2boW53ZBUz+9X+lCV7rnPsm7vLuLacY5ZkGkHcjHXXSfDIr3qyqFGlBUUNv
3WWpimBYjNtKTmwwtmthCmuH8M16JIkZLzQFaBPxFPy+hHIwfmEfe2KSI+xhHQcd
b88DnSGMHScrbysUyDr+ZcS5+hzw/3ltd3O2QSLXKfV+UbRXQwoUDu7HFMaAT9RT
S4x1hn8bXDndr/YKCiVaf1TK2Zj0x7kmGHM1U7tZ05KLjrnFiEtbOhwoaLq32j5V
D04WQ2mEn6JpH9yZiS6qWYA2UPOS2zGGLIZDwY2NDk+jcggpmgIbHhpnzl6/TYv3
cs2lPkH+/sV1shLKX+W9hlKtGmUc91/nP0zT+aiC92DDQ9kg53x7MRKJERwwbGML
aAb3KDwkAQk/l8/TbicAjmZ74MRJkanyhZDrsL2JwjV9t1kjpE1vfuIqFsmb89WG
o9LBm8YGYdW3mdyf/QVTx5DKJ6eqDSV15rWpv+RCKEQPwG0N/Hmqtm3IqHM2h1qa
jQM65DlFnWlpICjhBLvszYL4Zco6soaPNeZnHRTLkdJfFfblkpnc+dW5uwHAFXq/
PY+Ltpt7QM+0pd2Pn79XtE0UmaK6UKcbzmQnYIjF1Hjq72b1NRRJiuCgPCdWmv4z
Ra+MW5V4kFf1P1gUsVJpajB4LvLEm8XLdQgoS3BSTkcfNIy/IUX6VsZYFHBa5tYF
HTJaXyg+FN54q50gTOIuvn3AQSEswPGfutaB86+g0R53JQSXhoBJARqAfL5OwDAh
Sh+vIvvjxfQbcNHQ/EOuPJTUfQMiar0UgJchWtYkP47EhGwHhep3NMQdm2PNT2Rv
4SB2DcZPQf/e2orrwa1cteNg1Ny5Lrd4V5Xo44Xr0bnRpecXBSn/JZv4Hd1xQVMi
lpvU35UiUIMbRpQcpRp9fX+Jp/tGzNYmc3eWI/qDt5Q/Jse4cvgjI1DaEa3vFdjT
AsSYNZsw5k3DR3kNJxmGviDGgvhDqK9pt4UZHOjyQaKMA1v1BaIuB/MwWOqI7bfu
w66b59U/34XmPtLkcmUEJerjg6IBXzh6hUybQjZFpo6SlmMczifovANDlaBFa8S1
ZRiiqEMX2tCVKP0bWrPsQkeQnpV5GEmCYd8eUKjufpf7Wv9CsqH/vOCEPsaiRhXL
peZi/n6hy2w0sWMvuLrfIYTlJQP0VjHhC2a7Vv43YwKRFhCuUybu6NOuP2T+eBOy
yPYUkzCfOGo/F4y6bPCJiYrTLGd3gnYJxjMG8BuhIg0sUdSDFLISn8tuhvOZ05vr
bB4YtHRLI5l8syisAz/2Pbwh+9WDLO56vnvIZUFyanYV5XPNMyyFuBSbR8YHUWAG
c/doYYizwkrsk1xLJlK9rx2+q19PdBE0Kdjv189X5BmWuOqakNp1GPrGi7k0UTXb
GQHUjnO6C94IjciYpgHf/28NubnBO3Sem3JTrRoEmZYkZJuJBHRL0fqJhG6IyJqt
xYpqWUhtQ4ehLPtb+t2z4ronPeXmoKdGQINuSIbF/LWJxMvgtqgfs9+1dSULShqQ
zoMMveZ6/RIILzqcgBt76Gqf6f6yUQKT47rNOoX71wPcs2Q1RCi/HWRpHpj68fNf
q5rMuwL3k/XyKzITwopZ4O5twNhfvQHSj3FBsjdC/M8dhL1CWxzAA37uNZzHtd07
W7SnM3Xw42nQw8a473lOgCQdHmHZvWWiv/+NtvcZJHGEZl0ISBKvulcbtuTa5MTa
Ssi0rgLZAjlKToM9QjaR7JBUlCTSNWIa6+njOrVQ7XEj85I6pY5+aTjH+JfzevZL
8mTFyoFQd/OPpXeeV0LaJ1gjfho+U/UAGAG4au4ivcJLipNWNbk1FKC0x7NVFo18
6Ivb+fx2g3bR7Zr5tIidK9KaukTaZSFBWOEb8ihIjZ9HmYf+sfT5T/lw7zuwd6e/
snJFK/arzkdavFma/0rbL5htqX9d2KZrCJhTV1wOrclYbnnqfo504GXUlAe3MBtT
7bRAKUKVSyq3A6sOAmQLFCG28GQm2vjwAwqngKmF5AomZPhfKVJ5MJQ1ii/i64iv
ypzU/ysx2MYecFolSVE7knc0vrcHq8LEj5z1JcEMJscOXQHfZS1xj+wKrAPmQhye
j8hDmsYGy4ZdmlPvG7j+NinHAh0d49TyB24b3Ll5dZjiv+ANTbPwNGTKhI/Q8hBR
rt5w6VL08qgLa7NFYN9A9DHrKnv3o5nNafbFCsRVBwxc0MckgUjZcuoMv1XqYRul
l78wMSkuRQDA1ZyHi5i34T6zRbL8ZKsurNskFogVaADTkDBWzHqspDmQaemuzUl6
sE9eqH3fnAaP+6VeI1Y4SJD5Fyzk337Gahv5+WWVjnESkIaKoPuLS98KSFMA3+qO
Irju116+YsM03/nDKtNKRHAzhNc1MAoTrbhZsJ+kA3CDJHcirzZSZBfq55C22De5
F8VsxgMtnYX2SW1d/ZJUvK9rSlZNpF2bdViWSX8BNc17hAZS/4mgcH5BtCFLgYK/
eJKwNQBPQRODHVyL2uiL7DAd30XQFT4xNEmCCjFRKlkLcyq3yQGmMK3Qlp3klZYp
XV8qfr0qjEi1W5CPWXEfDwFwgKPGMBHoUq2iXTZTBb0GPCGcDEo814nAkV4Hy8n6
W8y84iW2n5FGGahK3LdBK38TCRrsYkj130cgmxffCAHDzg+60TclRC8xCP5ED37E
6L04f3lGLaDkMTGKKwkUUuWVBB29nH+AaROddQJ0DEafU7Q3wxLsq3UDxoQwBxm9
4Gw+KQMxjRN7t91i9K1lb6Z260BXJMXSq+R4YZUWZX61D5l91iHXx2EMqVTQ8swq
1tvOOK9vHS8c+iteUxUASSQvAs7u9pcKJQQO1y3BTEdLzLB5c/Z51IHxxcL4dplr
dhxLBplnuGjPMi9fGZ0D2Nj96Mfaq25Gd5LP84wET9WeSVXuztSU5hTiaLvololh
fXYXvuM8liaGzS/dbnVvtPjQ4gDKOQ0t9Qn3cs2zM0vdPk346DS5oaK2GZIOGrti
I35iIp/+Xi7sAapzXXb4HQ/atqf2M0sngi16oT21F+CwCchn00/59GXMihyogLz/
Ypuw/KcHkMugvhRHHmi9qPcMd6wxP7BnHHEQY1y+EUF8L1AGun7nYcDnXpfRRO/g
5YCFLyrSPz0qgRrGbT4z3GKi8FBa71ctvjTbDx1wIR250kKCKSJwR1/PAd0FKkrA
qAG5xVQ1EmGiwXM4OOI0fiCSA7tX0zqdQao3uZydyxMV+LzQJQNW7g7A0uZ4ZzJH
2RtvRWFU+9u5n3a/+3OjrIll+OWdDP1HWzTF/n3/KmpqoEbo+Bg1dmfpimAUk2/f
e5cgm0oC0xDH3YxfueJ7iktLLUd89NAm/SwxVyUWUM3egjIiIsZLU59IwGqeDPo3
lOUN3o6up4SU6xYn9oSyhmAPsHM095v5drlUsMW1a2GnOZOOLmuvW88rl91fLAH0
Vuv1U3eZja+id4mm1TLWfQ8sCL95Q7w3BXR9bqHBzvthZaYv4mPXmvWGBPJqSt5y
sUCVpRetR9XbyX+duPT2hvPt0j3dly80xzSfeU9sGdilAByIcr/f/nIj96gY/Zz3
TzlGOs2mD4PlUd+UPBqIcS70rgRqmSa5u8i6DVxMT4CXrtgYmO7YAHNB+ileuzyL
+N6zSVGNYqpPI0R+Qh6AvEtjEVUIcdg4+AdQFWe5WiLqNdN0KxAacSAXsQqhFXt7
E3FxyDBDJMFMr42oVyKJTeI57dgGPvD5w6hPwscywwlhK2OQC+L0A6W/nX6y151m
7VVe0Ko5qOWM2GUTzUdEPdDeP0+aOil/QnddOogDmWrAKme23i1TcboIF2SQlcmz
rpYqin1qXRcdm36f5Rg20kCPWL0W3oK4GM2LX5HsGQFYOjdF1i7TIOPFIOh0klOh
1I09b2L2/BYVKU5TT/7ORIgeBo+CXjkq1Q8IccOO3GcS1QepykB4x4x3QSXg9r5Z
WGQlIOfP9XkDtCJEvw/S6+ctZBNEIFCBUwK4ckOEpD2KkwNLoGqao3xTb//LLaQD
9vQ6kit6VD7obGNEXMx5CL1MpW58kj0jZPsliAKDwEgJF/FOigE4+KsMc0gg288U
q3GJgRg+//9S8ThP/dLB1jXqUCCJWwpLzDp3tJ6TtrF6deH8US7x37KmQtnvX9L7
4xrn8kMPSyzauAet69A7/aiAaq9eBQRgXlri2ppp2Qndw7qGJKMsKlk4VrSC4h81
+bCnNAalDexA7eThFmtc7/eLyQ5HVA8dB69nbU2jrLTI7C9CtkpKzh4dKjnR6rwt
3iUBAPAKDY6J8DP5iTebuPUEoNZkqlBCKTh/iH8hQraY9AGPD+ddbT1l61MjLiKk
5wWFHcRBeqUj2lE8NxXZJCN5tm1AV254S7bH+EdZpIQlDM9SI/qpOoJV9SupNCxi
G8QhypPaO/swna9dEXCXvEtHOYMQ/KulgkMK+roX0okmfxntrO2Rydb0RXgR/xTK
WkOY41fVwco40arfttsqiLpY3znmB3NNPx8BFlbItbcEW1vSDdZlGFCRQyiDwZUm
PgD14jH2ZpridFcWmlBIQlaFTfG/9Nex7iA9IYZckFHBD9wConzNWMR9tf5RD6ah
nLFjjVNuv93S3o+kOBFugwoou55MKO/Pj2UMKAJUDr8uvHqgsipvrpantAP5jJNr
MT44xc1ZvD6qcL4YaNwdtWtWrskJ0c4UdfPdsji42lx1wKAs2V3YHF6ZIH0pwww1
nYdxNqQJ3qd3nuI0n+fH/wRpM3P0dwwbvrv9jV6/sIbnH3Qf1SQLn8Neq3N6B7xL
ugx6LUm554m2tY9ZDydqKfcysXx/EVquT/31vQyMaAGKyZOe9TcG8bnVIhmKIpXT
csbze91Y3uOK1j8ddECI4Afbrs4rMwaw9bGxVyARE7nO1F0WcsKfE7gxGZs1VoP8
q7cTjW2cZ71vPDqTfG5s9SZ2tV41uUcutNgQ8L+rZCq11ZohA7nQD8vDrx1rlGCM
NDvQ1DoaTDqi9BahECNMFO6kiqSD+gzUfEMOs0w+sVrbqr6tUIkz+6BTVrSx9Iol
01LYXMyEfiT6w6j06YlHpiYu3zf3/wraMRujJRNX43hJ4TYHNxtJD29eyfab2oFZ
OaDKu04kv1vDDvniZjyTesWyy+qM1Om5M78rYsRB2CbkyFVkqzqxAqY4IKf+xF9i
G3ZrVcWeZ4gDHSSLJseuXhzwJiyAx1OXRSxMNvww7JoLnEh8OoTziKKPfSEXjy5z
J9ZO6eYPBLt13najWzizQNP4fE+wBAvfljkidIKOD1R8d8sG4bxqRpPUErmbKr4F
a6f5cyTz8BkFcWp0xD5jVXpsGPy9m5ayaNGxzXO95CyQtwtSvJEXW8xeQlG/Ktmy
EgdoJiODqnpF2gxeMpyY4SPn++Yp5em+P4vgqWGkNwZk3tEIeYx7fNBpT/Bytk5+
d4gsCKQ4IjOFTdlkkqhiQ6Uio93AL7klmbngoDkY9xe5fkKXITU1pm2cVrAPORRx
PNXXGBRrTloax9sAUznWnW7hI8P+i5BTq7A33oJ5jUyDPgD7JckGw9lXBfF81crC
l1UB/a5D6JndTAVLvD6bJiSn68JxaljZOLJJ8wGegfjeMihUPpIbHi/GFqvFmXZH
p3oUq2PPnbPndqhsBMYMuhxwkFrP59HZZXO8YBvi2j4mKmXh9S/ansf0ybbTbRMt
I1PwZI8PjQXasFRG0M4m5K/JCisU7QBMBNrIM5HAO2tnQcYa3CP5iuasVHHAXp6s
SiDPwoaIETxsjj0nGMIJZoSKtAyVsZ8rcE051jUnjLXJhwrTY4uySBMLVijPqe7z
WqClvBR0kvKDmztRkd8Qywe6tUj/bgTGLjy5QS6w0XilVAhpY6dWNEOsJzLVcK9y
yzLfn1PCBvtv0ArDdQBqeHx5y8DWRrKeIJ4f8m4bKg9AHRyyFgzTKAPI4yp/6VeO
IwlHoqoYEbxYnpFI4IGu6/IWqGbkw1m4oIXJl6YMGkW9f2YSUAVI5hiwTqDC4lqj
ClCR/Dp4XLAHyIDnf8uEMf+R0gOG2f5sX3I2XIrW+DEyDCetApLfDgpDZuCrO+Sx
vbbajyIE8rUFjuZPPy/r0+sKAvoQxjkIWaIuBMEwp7gWoPSPQj4Ci9UboVm3rN+m
2NbbLGGnndWC+S6zXIiPqu1pYtn0PhA+CXn/7nfe5aFVSukfYLbYMo1viwC+Y7ig
JlcgfWeNVnaVuJpVkRlLSXeT/ztBsD4K5KfS0HYWelZDfHuMxqbR7gkQDWV8ZpHv
ieKevN6vEzw/gDKovx1tX/Ac0cvRdszURLsD7QQOPzkNpr/Jn9/mRwdaq75ykDBC
YvQTSFY2Byr4YeUt+wAA51vdcmfNMyPFPPh+da/adsjHs7Y2Bu1z+9PNsTtpKynF
0OPbpM2vzSsX1E4f9zOc1sBnPnEQgY0TJtIFAbvUlMG9fge9ZUwonbv58/EUMhaO
nEKfJajmzb/BliP85rwfsCToUTHh4SA3pul+egp9bg5sLp4jwBZpHBXyqEugcvP+
1fNpbzEpMunXfp3l9p9Kh4w5ISKeQmJuAtdr+tAG5P3KTL4Yq9gKydiubg60Kl8R
XG3p0TW8HPuL5SmOvMwpazGzGWe0mfkEVt53f24zmdSlnH2Lh1wGcTMM2MCzSoj1
GhaZAbwKSqcetUONyHoVaUvSwMG+ZGKRs0Pz9tVWqtP8EEdUi4+UNwwZzE5sR/fV
IF4WU5nlo50ZiQb00UHgHwN9CtQhjvKfB6lKN5IOBgZrzlzWoUOw8wccX0Zz7eZL
3TVZAWjd327IpT/CIA7tV/ngicEULX0xcKVNXLZ6FZHf1VqUE5AIjRH8ZUvRahWp
+AWAu9rHmtpG1tw2HKAkGch3/5tXeGHHyXEM4PcRQYZK6jvRkm7I8X5t6TayGzz8
AnqK4SF3XInjlFqszbnkug==
`pragma protect end_protected
