��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��CN�M��rY���k�d��%�����]1�d	a?���u�P�e�q{�;&nĲR�OL�D��M��:O!����߸���:�6���R���{=I�9`�DW��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�I��U���B��<s���f\�-d�o꜓��
5����u�9���_=�����C8���M'�py�tT���)9���q��V4T$��G�CW���5�` Ă־�7�}L�P��$�����8��
&����w÷��AXR������3t�c#��@>���:Ј=1� ��|���U#t�
ည����du���y�h}"���뤳>���r�gz��ir~���ظ����r�K�%�����y[�~n�7�=��떒����K	N��.����~�����v�ρ!��-��>j�p���MZn[I�.��\�8]�?I�+��ˀ?�(��53|U�.�>}쬤"pof�q��t<�|�U{�|�!�rDl���9��*��x�&_������1WsW ���o�'�D���Gl6�̧=�d����^F0=u`d����1��Wh�[w���`)��sUP�ǩ���#F��=��}tjKp�����U����]qV6�[� !��Ș1'2?�B��Q���N�'wͯ��̏�-�<L5q<�^�ֳJ�y?:�scBv�D�H����>[7�8V��N�V��{h#WVe�z��I��rR��]�ڡ^4�U�D���m$��׷
���-���x�]���[�a��՘q�;LM��A�V�D�cͺ�?�nnS����w�0y)�R|:>���e/]�N���\�ޥ��H�@�'Hu��T�p��P'�K;�2���A�#���H�l�>)�a9�^:TW�	c�$"��o �E�������N�K�&��kj��R��&]��������BihF/d�N"�w&��b�+�i�a������E&y���=��=��zDG�\�\}ܧ/	�B����r�Zp�廞;�.���R��ߨ2���(O�T���/�s��]M��=yV�g��6{�:5�m��_�ʩ!Q{
�:�>�`p����8gkۿu��`gi1�����( 揻d���t�8kI~� �m����ַ� �����{_�c�-3��@���L��X�¢��2�|�I^�Oj��>&�gW���H�:��_:���ܮ,����`�.�}abn�>3�z\e.q"ό?�-�2��x�x%�=�T��-���t�/w�w�m����3���3|cc�z�O��C�����L�[�!4�
�P>搙k����@:�[f��C��_{va�b����~�� �W ���qV���m-��ڃ4��"�G%Q�D�-��Sɰ99P�	�6�>�ޜ�z�=Qƿ��`I���eܒ�D ���v��K��M�=	�t+���9s��[cjD��plȸ[�^��ɸGQF~��J�8�q���4���V�,l���7�%�QXK`��6�Z%���sR�L���%� Ё�	�k8V�w #&q�|q�qE�\��J�->m���ꔼh��j���%��ʩ	���;���%6�rS��Xq���6z��ۣ�%��r��w���.S��"�"�"����M:�^�q��I��1oZ����ݙ&�y�Bn���w�������ͧ��1�;�R�Ig�1U��L��g�ӕ.�V�
3�r~7��ڃ�h�$��8ƙ��Y�w����`W��#nҸ����>��UɄ��0(��
X�Q �.;7%������b���Ky�����bY��q�E8��,�������=
�ث���jr��P�����p�B��^Uz���� f�/���-sr3���{:5
t�+%Ě���G X��Q�}Oq��B�9�r��/�DSS�~�E��8��(i4��۫�mY�c|z�{���������P�=]�Xqljl� ����\��Ж��b�VچO���1��책 M�1&�lA��A�Rb�/:�������.>�t7����7rN(��\y0�~1Cn��v��0�Zo�^���Vf�s�P�z��h���5�H���Cd�����*:Ψy(�]1	���<;��x�����ߘ!���QZ�9m�T��m�����B���<3?�J̤�}�ޢ��<�
���P#�lb�2������"|�ۀ�mB���X�;��DK��)c-�p]���Y0�[?�t[�%�GyX�}I2�;!���&��i�9�~�a�N�G�ܦ���T�N�{�'�e��k�Qhҧ��0�/+�R{0����~��o3�)ȝ�]�Z�ba��*�$j����N���(+Ĕ_	������c���#��j=���R�f��'�g�6ī�~�O�j���y��6=G����FdhH`t�۔y>�*a�[��;���C�<?�D��}rh�.Y�������]�D4u7#�t=�,8���ĳ9�L��(ڋӼ�,*%�+u
�'|��՜�j�FCG�,B1��f�/��3a�"_��$i�t[�����Lrh	E>5?w~�����>p�JW�?C�(^�%ĀV�#�Z� +�h�ʿ�J#�nz����<�Õ���A3��w�=�>s�u��|��.Ÿm��:�tX��8��c@cRJ��n�ҝ�"��ө��,��"�yPK�vI���S$Uh�X�¦�W$�4�Ơ�6��%}�]7�����K[����1�	������b�X�S���=)���(OV�i%�K���)�d��j��-��壳���r-/݂[�z�~��S)���O�KF:]_�������xo٩�{r؂U�}i:̭}�F/�����aM¯gdr��0�qy�lW�iÏ\$|�b�h�s�QU'˲/U_w'�J�	���4K���أv❉QR1R�΢����쀕�֯��u���|�G@��w��H+?���o��nݸ%˃��+���(x�# @s9���N�w��h������/0-�ck�ꢶJ_'����*���r�|;6��8�#�P��w��~$�a�i��Lpd�JTȦ�_��k�]-���4q9̧<�=6&��T��~���=�T1)�SxpYj�2g�V~�\��ER"Z�~>K�w
a��������T"�Ѵ�6L���}�������v��k+n�|��Ȓ�7Y6��:&��	$#T��(����i�u_�.����O��k�H�����K��95�\ $�� L~,�fȽ�,p>J��0*N]0<�E��g^���o�F1�)��YwɄ&O�l��й#�����}c_��c�����6a�V�ID�����,��
�W�p<"��/9D;�#0Wo4I]�̐܌m���Ho��� �,&=�eGdX����^6 3c�����R��fWU���#��@�"-ZKE�x.cI��
�9��a��1b|��D�aYȐz�^u����X'iO���Bwڂ���a���z�V�YCp#�T�d�o�ȗ���@C$l�Ll�R+2˗�@O��'�����>vK�q;>�]/����aR���A�@�fR�k��ź%�H��+e��m���Sm	�Ҏ�,:�m�[~��]�>wHP����MV3Ó�M��4�Ǹ�{(�3

����y)��uM+��� ��gqf������6e< ���?:#<i��Ӣ�=�e~
8�kᚰSQ^����?wn!W�KU&����ߒ�;�Ų�s��M����c����O�_K�.zb���� c1|:��y(EDT���j��4�xfXv��O���	���g����l�Y�ٱ)�C6?��4����D@��XK�/�m���`��7h�*��YD�W��s!��}��Ɗ�"� �ڼԐ��5�R! JG�y�	gRS@Y����67S���ÛM��v6��皟"P�;:������`��츍ȫ��q��:�E��ć(Q	�S��ek$@����â8VH��wK+t�\�>�"�|��%�@}��^��Q8���ܝ�5r��O�o��*�<�"ӑ��7�q0VhXt�C1�k����`UF5;���#�5�
��Hj�H;�1mF��2��P�u9cxL}�jֹ�.���R$Z+�]�B��?f�\7��j�|M? �|���hٵn���B���9�a`�2A��U�M�Ԩ���2��j�,	ȹ��a+ǐ2?���J�X��yU�-�A��ʨ:�t��V�v��P�h@;��~#��߄ȵGІK۫��'�R��u���||����u'�6��Lq�a|��\� H1z��ֿ���f%-,`����_R�(� �O�4r���W$�dǌ�G��p�?�y���3��k�N�z���l�ۤi�+�LnɆ ���zv�ȑ���Hg�0a��[����I��Y%Ѕ�qd������od�~���*9�AU5�#��w��W΄,5�督��5�,Ca��O����LKy����<md�;u�,��
D�s�}��杍�84�n�sΩ���p�N��X/$f��+�XC�}&V�[�߁>�}s"4d>�1�/R]N� ݧ�p�aY{���P��4�1���y�PC� ^ھ�ݼM=�	����լ]v���e%�DV`(�I�B��t`����=�Q��m�Û2_�4�i-FD�Ni���"��һT�4yQ-�g��122�MI� ��N���b���B�	� ^�ɐ���WJ�m_� �(ݱW�D]S�Y?�P_����1���M�G!��iŸq,���JX���˱;e݃a&%�{ޏDl�7�Y$XN�<e����:�2������q��Kq���Y�V=+�����R	�&�7<��쟈��l=�g�w��Eg^Q���Ug�QPi�9�м�i\�Z�`p���sM����kqV�z�J���VI�h���MYhEpq����#��%.=�)��[�5�OOr�n�g�2D�HH��h����:�q�9F(��ݵ��a����|qX�:�5���^������(ҐA8�4��L��+���J���.��d J_WB�[i��Q���8?�v�N��/�A� A���QK;_U��Hc��h���f��'���?��#�W!��6�~� V�PY]�̰������|�^�GW��.��*?좹d���"���/)�Ÿ�3!I�ЯI�#�%{�;L�K���;����2:1BAEI�N���ba�X|�C:���X�FB1���K��	�T7d%�+�;��$Q�Z�A�qL�ɇl�e��F�LUNQ�Vٞ���Ž�YX���xX�'2o2���"�4E���?"�_Sj��5�rL��~��/=z��5�=*O�0�����C�@eKnjX��-xW�$�8��2��\�k���FP�f�C���wo��]�&+"<�����'���1ե�s�ƐD�3��­M�����v�|n��������]Je7TeX�@G��t,P3B<k�3C��I���Y^�:��$�\�y9Dx���L���쟚]��f��U���O���O�o��&@Y��s�	s�¥�{HVu*�c}��Q1�
Y�M����䁼�N���n�N�R�GRh��W��r��?�'[��b���lo��sS�8�;��q�����P�(�z:l�=W�7
��j�\[P�Q64�����٣
�Q �i쌜uUh��amr׹҄��l%���Zҕv䋃%{G����*�s|gCkh6�UqF���N�d�c[���Ei�vP��Y~�WG/ec;�2����'���,7�F�$���׻u>�li��8]܆����;O�E4xS�y�5Zb�P�A�IV�)�g:q�mB�s'��l�Q1^d	(�)�0ȑ��Ƚ`
����䂅�����8��oco(�Hq�\~�[4ٯ�� �؋zQ��:��[��-u'i��f�^]�;����l߽�:�q�/��{���C��+��+��r\�`��y)(Zy�6��N�������S�!�C�U&>�m'��F�:�m~q�a&Ș[`*��a,w�{:Y��1u��e�_Cѹ�W��z�8fJ��W��*���0*fja)]<\��r�Og�8e��V���B[uƫ�8[I%�DV�ZO����y���$���7�/0wg��han��\�B��^5���_E`5��=��-����f��:T���/[A�<1	�O,��F\�n���7�9B�ƑSm�����_ar�tC�+�q�P.�(4O�\/��t4�sY����;�O�>�f�b25閶6������yUbkD��(<��Y�}�+iB_��uJ�c�A8̫�����\2���sV�<p��"`�И�9�v�C�$[�?�>#+U�� ��G����,:LQ�C�v��;4�׼,j��Ɲ�D:B�5��y��voG����� xA|IJ�##)5�5}��uڈ�ҿ���cD{:���=�G����-�]��0��34�V�Ҋ�ًx6O%:�!����5�t8���"�bi��X_�+f��'��S�I
@�Yfhef����8n���m$/�P� ���:
Ӳݙ=$��@��~�c��!/Vp�'mJ|O?����IDy���֝����pC����Hx�� L���Vq}��u>�49��r���
d�ľMg-�T|� ��ۡ�{]r��|�K�����,�����=� u҆xf�����������1�[6=�(e\K0a �'�]��i(�F%�U?�z����ï)�1����3��JƋ�����^;���/P|�����z���[�~�竸���G�����������2� ���v���̤~�?F��!�$�iu�	LFbt�dR56t����소��s
��V�SɄ��<�����U���۷��P�s��|S]�E��&z,|f�hRE�9���rH��gsݶ�JܳB��7H�J(I��RR-�3�"�����u5�k���م�y�+A�b�o���8I��i��-�����#�VH��]��e�wx��� %P���)+���Y�
�������$xL��n��PJ��U�Լ@��q���_f~R*@W�.L��!��A{*�v��=�K�o���^����J��"�[��'벝�s-Q�"]�z�F�iF@L;>�Yq�:��}�9!�	�}��wT��A�5
*ۻ�JG����M��u3b�#��'k�곏�Z��ܢԽ��ɜm�ǲ�D�i�+��_�C�A��E$"R?�1�����s2!E�A������'7���N���I�kG� ���5u�O:�/�i�Skىh  -�^�ƃ���� q��N��\�sI`���ŲVI7��Oh��3{���[!=�# &x�����]�ɘ���L��MH�M<�E�N������T$eyH�ނ& &j�w�F�E}�kZ�:�f�Aƈ ҙ�p� KH�߂��ٕEざ
ز�*$F�:0�'��"۩�#Zd�Ck�FbM�;D�B����8%}�"2���=2�|(>)��#.�xK5���#�=p ��e��F\���zn
�:쾄�x)6��<��1����������P*]�������Sڱ��/�}�<���[�@eU8W�-����_��߯t~������<�����ĺ�m�+�/=��!
�/�t�w9Sj�1���� n7@�������37x�#�\������,���))o��iH�0��U�Ғ��D��Z�x�
�*`�(�2����������(ۭj��P��+�� ~��~�5��G4zvXT=���+Z%U|�1�ev��i� �E�4޽���x���H����f��D���ș�꺹~2�׮tl�_\`�+���W�����=�׏�Cs�(�l��9���P�n�{"B �p��V�qV�QTeP�t<���l�(��$�@�{@1��W!RXQH?^�5�����j@��[d�2�Z#q��^�uy:�E3<�V�2�-���@?B�������9J�K�r����M�rֈ�&'��ka岛c��h�rd	��>B�q�f3z�*�%�Y$���`\q�0��w�MpR3�g��Z8��>��X�g�?�^�;�4�V� $���Ų��l���h��,�u=�~�ߠ��m0U��,*(�w�b�Y��u&9I߲Q�*����w�ώ �s�X�~`�l_&���r�d7�X~F��@5�>��K�E���5D�Vi���2"�Bt��[+��&ޅ�S@�1�� uEpM"����Q��C�ל�\bA8�@oc�v/�$<��JQLuv/(|�/�_�k�}��衘�Y܏ݨ��	B��چ� a_�����̀XZf�'���B��mJT�ވ��*��V+��~��N �*C��[!<)J?��멊{.)�X�%z#�D!q����оif��ajvR]w�̀�;��>�b�����U;��o�����+��MԡB��d��=;LT��%G!n���#��2��񪃻a�����E,(*=9<hc`m�"K�"P!G��1`�_��u���~EN������<�3���2�Ԃ��{�����,.��&�%Sp���Y;m1|��c�펟rb;Ms�`�ۑ���)����d��y����)���ŭ�4-V����*��ʵ\	�� �B
t����[�8 �k�d�c���5�+�>]`�|R��4���n�LXQ��b 8�U��9ⱂ���&��T�Y�dU)�	Ia�:�;n۰�	b>�&�Ǎ�Z^�1�4�/6��Q�:�O���#E.V6n����U{&�He�u�Q^F�������B�E
��NB@�_j�V���b��̆�j2�Ŋ[
���n����U$,H�K��7��9�-p�0��~L�x�6�U�"��6H\�d��_Q}"&�H�U����� r�-��.��VdH����(��e�Z��A���`�\��1F�c�L�X�%���{����6�$����-|%�6���
���D�Bg�����2�'��+�����uKx���gΖ�.����\r	b���Ϧ]�a=���Ɯ��bT�d��)#B�����CϬY\$ﳂ�8�D��-�3���P�U�����	�_�U/��C�!~h�a��H}>�"���?&�4��w>*&F�57P��]��t9Zn��|������Y����D�QZ�kS�HaȚE��Ĕ�J&
�8���;I��u&�2�����lȔ��77=	��E$���g�3v\�������������GS��4�ti�7(Du:�Bg�s9J!�{�)���.�ȭ��)ʥ���H���χ��Mv�Z6kG����#W�b��B��Z�a1��%l ����Ս�R��]xd���Z����Z]�`rBm��G�$j�v�@�5wm��\�֍�ME��@
��b㏼�5�vk�����!��#"��ƺ<2�i���@x���"��b��y(/��O>��E�MOx"T�u�"��LGr��gkT���:g$yyL��F�� ʪӵгx�����cg�Y���̂i��G7��k?<�	8Dce3�V�k����w�d]58�va�9"�塡7mo��i�m�F��κ`�o�>��R��$�i��$U/$*/繺�w57$]��Z�v��0{�z�5'�W�.V8�5�$Bq!�Q���/1�tYq=p�N�����%@Pȧ��4���z&�X:v��]�m��H��e�I�數)�3�?����,����{����*H_G�fN-n���ڦQ^W�0�K R��{�Ki8�'V�'�ݱ��@�!�����c�Ǻ:�ƝF�"���,@
���Eԑ��+RAO�QKk����,�tP"�gt��K'0��~Q,^��h/��2R��h?�KG��Pʎ��G׺A�j���,���j�Z�7��E�Q���2����o��	8����$��m�R�X�H��)Y���l�N:��@���r@`K>	'b�*nO7o'��-�M#��	�\z�� ~�\�s\�TduD��(wh�|�;xP#iu��>�{�{�'oXs���6��s�4 �{�џ�*ȃ�x.�Oáb�E�b+��E� �`ug�ո��=P�GtW�G��kT�o5$!�����{:| ")]�-'1�B�zv����u�~�T/��d	ը�Vg��8��o�-���)�=�����h�뽧�L%�rPF����-�h40�]g�a������;@$��EA�,f��q |�]YoA�h�N�Z�2DDb/4Ly �Ә��ru�*��BxT������쬰Là%ueH�X�6�NAҒ����hSʢ��#0�,��.���n���)D����+g���R���*���|Kj�&�7��N+���	�1Y�2+����{Jv��?�	$�>����v��+!|������DlH��rT��q{�eD�-��0����w�Ou$��`�Yu��d��
�YiIyQ	�Y.I��4�fcƩ�F5�Ǖ��VCۅk�j�����[�5�I����I_��B7gU�_�_!�@!�s��"HI��_���A(����X���t��Q����Dq}���P>"ݿXs5��!V�[�T��n67<���Z��8���!i�����j�č�d�_ -������~��᱇���6D �rjk>�밟�i�ԀI XX�F�+�oWpMA�s�&�P-˽�[D��	V��h��&�x�rn��L9w��+��iY3\z��X�4�í��������$��uZ<O���(:S�q��ߊ��sI徰h���1���W��Գ���pQ/
�֝7���>���m"#Y�SL�E*��e���l�F8 �
�|d�M����|OR�v�_�J�ɢ
�� 8lT[˖O���m��F�,Y��� �5�8��[�X��3�oe�տ�$Մ�*�[����tE0���J5�%0">V_e�\ǔ�Hcsj~|Ro._	_Z��i�z�ǵ�_����S&�Q��liP��:y� �W��L&.�1z���}�yUEJ���G�z�k˔IE�Q�zt�� <��!8\d����ݨ=ͅ�dUI���/@����Y�vo:��˦��fK<��,'�vs)E�S�3���i7�!yh�l�mc{����L�;�vLͅ7��зb2&��.���GG����;l>X��<AkW6Ö�R=.��ب�-���|~(�J1��;�%�ƀ r$�ː�N���hW	�n-M&AB��F��Q6��Ҡ�]��:�d�2�7����?4op	��zj��cA®�wמ����A7+ 8 Z�5[��^��s��'�j�{ �q���s��ܨ����b�}�G["�[1�F:���x�6E�mI�X��:3J�C�ʋp��`t�#ϼT%���GCc�5�
�����rU�S�Eqʖ�����|w�p�^��-M�o؆�u?pn��v��h�L���B����I˒m$�o4;|��J�� �O�����Ҧ�;0P��U�ݬ�F��!s���5c�yrk���j޶���Te@c�R�㿑F��9��C�ہ�&v���_#�m��t��.(��*j�9�O�,v�&2�d�vvQdI?�\��|oqk�]<8�����5�DGt���?1��K��3	����G���BFF�����U����<��ŌEZE�!�ʑN5����p�7)S"t|W�og,�]5OZ���xX�F�ht���G���%��a��K��r�S2�N��*��#�ə�+�-@(k�6�
��6�w����} U*���4�w��5rl2�z�
T�XLf�5�	{�r�D����p)I=��N��xY��*����"y��ɇ͞�V�n���Bld��.��E����z͔�P�5���q��u����T`ݝSB�׊f�i�\�;��/?j�{伾C}��!q76�a�Z�uWYrZ.�U����l�nd�:֋�U:=�LU�y���gq�Sأ|��5��I����V�Hڧ}G�A��{����hsF�w)�2V�t�2��
�[|f��#P�8��m�J��D�� ����V��Ho��E��o�&�utش-]����T#���[n�#��J�[:��� � ��jg�
.˚�[��VY*�n򡹛���#�N�ƿt�bzy��c�8F�m:|#��ӭ�"�91��WM�9d�-
Ha��\��t������Yc��z�y�{��='񀻓�}��q��(䍷��奚�v:��q��?긡5��̃@Zgk���Ǫ�J�F��ʐ��n���1sP� Z���KS��M��V&79i�bw���e��	��a��X��J��Z���yEn� %�&K`������A����OU��{CP�RT��Bqlv��l�����[Ƿ�Ј�Z6�H���B���Eh�9|��\����!��=�q�v���9��v�����D@�E:1��y!1+�ߌ� �Cɖ���a[����4���3R���_����\���P��@�<�������S�#D&�,jH�a�����g���S����%]�����Hg,
�
3��|�{(���LbBO�%ʖ7�{_I�Q>�Ψ��iФǅW9b��]�LB�1hK�K�.�|
�J����_ ����b�ϰp40�E!ߍ�]n����T+A"9�f�;�U�#�j�Nj�F;�u����
�>��j�W˛��M�^NK6Z�'�����o��i��u_vst���h����jD���p�밡N.��яi���Թ��S�Xm�.��S-1�CM�O�#^=����ն-Q��ͤQ<�AD]#oYˎ� ��mK|x���K=����`�L_M~ڹ]m�'΅VP`C	MtSm͛z͑���=�
>��cU5�$�����B�Ԓu�=��}��6�">S�}**�'Λ��#��a�D�y�K��I���ԣ8W6󣒛�38������b&qZ������+���LW���N����H8��l��X�<�X2�V�g��v-�;���e���~ݍo�c��(�����S�P)m��D{e?-��^;+�"5L*�<��Jf���|�����t�n�%��]��޷O٬	t�ȥwlWm"��@̺e������X�W�jG���`���&,Plh1	'	\Ҭ��:�D'&B��R�ɪi�7e�-U�&	�x������Qh�ʹ?���B�2:"���1�?$�[�д)�#�ٶ@��*���zF}���w:7)�7w�!v^�D����]-���l�*wqu@d98f��Ʃ�m��	�GE�����	�A���LZ���)[}6��m*�<� �ꌅy�HiLS���Mh��n�Kb�bǘ����Z�'�s:8���������|�f�o:-]���e�tB����˅�Ϳ�t���eZ�#���/��:]c�w\���Ҟ��8L�21�������s�zp}�Ru�7�i����[6D�;7v5vڐ}�.>p{�M��JD��{��P�ً7A�2ކ�&7/{�F7~�e���Ƌ�$L[[;&ɕT�y�=y`��,r������^fϼ?�Yr���ܦt
��w�i��>H���f��4
��K|7Rc��!�r����6Gb���	'2R��/L�Ũ�'Z������)c�~��1�Y0 ���d�m��������u)t�S4!v�}W�;>�p��x�hى��%�'?N������u�X޴�.�=a&~�"4Xt��ͮ����	Z���Apf�F�u)��e\�
ƺ���/��D���B�Q]0�9�O,��l7J�E;&�a֑��R��9��?��2��tXtda�.g�e��ME�1����K��w�	�����e�I�f���;�R��%�ɒS	�= h�3���#(�lX9��L/^&�A &R�����yP�{-$_1~)�.B/qd��s�κC�)��7+k�<U�rC̫�LW��zhX�(ֈ]���%�]R�?�����^5��\CI������$�^������,��V_��MI�O�a�E��k7|Az�ׂ3t�J��V���������_9Ԟ��7�p���STL��4���]�H���]��.v���gd����O5t�*y[m�Gx���摿}�r=��������8U��˙���L]�!#�A@2��K�:4�����~ĩ/t��<C8Iٺ�����ڿ�f���[�{Αv[��#T�V<(�Oqp��O��/?�?8
z���vu�x�i;����,J\B'p|�K�B�"���g.��-��՟䒡C[�L!
Bǲ�����؇�b���U� ���&��-�[�p�6s��OF��OsTk4Gw[���b�쥶��"S2f*�W�`��|�[���2�Gp�4����"J� ���Ћ 2Sڋ�l�kb��!�+��=$���q����3�|�7w&�M���I~n�Y2G@bp�z"ǯ��q��7�t���L5���k����aZ!��nGB6�����i��,��b-f>���}�Jx"��'���U�9�m�b�u��W�������ˀ��z�N��n�o #�)�Č0�/�e��/|w���������˃I|�,���Ǯd���.A��h��U�Ι8����g ʢM`�@҅�r�wHÔ{�|^i�3+o����]��JW�֐�V����a���f�cֈ�:Y� ��d�b��]=]�V����N)V*4��x0or#�G!z.t�3�S^����{���Q>���M*����-Ŀ>ٌ2!�(��QJVE�yzG�mTȽ�b�ո>
� ԩz:tU!kx��_��d���PxZ�������ݤD�f�X�@��]������ڥ@�;V���C1���`h�0����x��ƒm�L�$=�O%���v_���㇛_]��=���]��f�
H�������:�8k�.^ݔ""'b��hO��2eG�+����``�{,��/��A昗��	�iK��)`q�]�
j�z~d��v�n��R�m�1�Z�~q[�!C�o�
UR�$
ȝ�^��)t#�ᏣH�ז�9���Ӫ	*��-��?t���O]�p{�"\k�?�G�/_v��Z���$�y�5��!�xOƹ�+��W�	�y��Z��İ�
�c/��dK�(�IZ�;��{6�	Mp&Db#�6�L���CbݍċC��E���h����?�b����`�z��P���%1jm�G���ރ��=X�o�Ï���uX�H!_O���d��h>m��G�Q��{#/a�:Oy�m�'0�
H"��1Q���3W�����aZbT�Ƿz�飴�G��l���������O٘Bxyb�z��苟��G�hA	+�Zz)���w�� ����_i���Y��Â���	n�?=<�"x>�C��#��M@�\�儂�F?�x<<Uz�>������ >�%�C���:���:�K�-ܑ�}���04������#+�������f� {6ؽ�ˬA�K��)2q���㥠g�s$��%/li!�8i��t=��HY7��v�2K$2٫�C'i���9��>��{n}.ޱ�)��j}B�X��W5��K�[ (��6�f,8$aBV��Xs�u�3�.�'��݉ۊpyf(p]q����XޙN��)��.#}�� #Qm��K��'��-�~t�*�/����d��vW�Ԧp�Q�J�����$��l�L�:�"�o��*�o��YZ���zC8C�B�9\����wkh
o3��(SJ�Y9fy��o��HX�V��JX�8<�c
�PX�}I	�<=T?�k>�vӳ�@�B��|���B�Ye�ī�`_<�=�����{�uD(y�m,� �WG�b�i�|�@��O�I����}������On<v��4ܵ�-��� ��o��꨼��s�;��4���C\A�iy1^�'��5�E����RJ�!Z���DA�`~F6�+>GJȒMz�ُ��1��-i?(@�R�2�c�Gi�>��D��*���/��t�T����AJ�z��@���ư��������s\:����!�>��p荊����9��$٥P�O���w��K�ek>><U���]���<iV��$�:�j,zdܺ�'V/cK�/�#��M� ��3(G��Rs�T�r�N�)V�x�s�I�҆|R�|�������Ĭ�X��j�Gd�"q�Lx2F��O����Sg~CJS~ �/�}sTz4�ٯ�$9�����uJϩ�UN/vׄ�1�ip��uי
Z��1�վ�X)M9"v�����Z
�j���BZ�E�D2 e�g�;��?�6�:^r,b��,��,V2��#�<�߷�I�ߚ��,�Շ�u�����	��������^�;aw� ���n��Xa����d�����$#�h����Ȣ6��-���:����dۣ#8��珴��*�'�.��6ōW{�x-���6^�Luf���ֱR]p&2�x�&6��3�<��cPĮ�	o���GP�b�5�YA���6yVDk��^Ci7��6�o�|@�hj�R2ڳ������{�����i���/�f>�7�-(��W-L:�g(J^E�[j�/�oG�qI��.O���Z#�CI����Y��}��h��aͦ5�HUH�|���f�a����]{�W�=�� �={�J�j �p�Ju��<T.����Zv�c�� hxhES�	l�ރ�p]���
s%#��c#��?:I����}��d�FQ�O��j��2|U/�UY�57S9пz&�G��'*QvH��r�L�M���A��aǇ�M���a�ZH%�<A5%���ϚY������4+���)E�n=�m'g�ԉ�C�3��"a��g�f�������)�����S_�|��{y�a2!��cxQŔ(9��o�6����� �#�t����L��*[k�|�lEnxT.P��"���x^`NI"�A�"P:E��g�kZ�6Ӟ�U�k�E�}r�t���L{I�~���ԇ���nDe�edK�l�(3(����Ĳ9N�l�f��G74���gm:#����Բ�m,Q1H��i!�S(��t�0��e�|��L�p��
��ȍ$Mr�U,������oqܫ�o�����ʅkڗ#-p���0�6r���i�ي�Jذ���Z]ٚ�>P}�m��u�ݳ��(#��	~��e4yj���BeV�+@�D=4�ٗ��1�
�\��2=?���J����{kz2j����ч#��[Ӱ�"�u�E/g��$M�������-�QuZ&�3'Ztz6Y��vOB�Ϸ���:OH��D�7�'����1b�4~��#򣫃+���*r_���V��f*g#��3g��B&d��3�uow��o˘��㼰w�����e)�4��=��x�&C-���Cw��O�H;�6_�� �8�(���hӄ���*<_�a��8��[HQ���A8P�=�B �%�� D������~��o�H�d\��K�8�o���6߶_�l�O�$z�}.��ʩӬ��ʺ�.����WET$J�ْ�:��I���Ԁ�1Fy7�ߏ�s���߃uم�L���@�l�#Dփ�c����h7�N��"~��ܩk���-�B�f_���2�/����U[�TJ�T���e��e��l_�|-ō�euG%���I�Lėmn"A�T6�TN�'4���m;���ݪOa�)2q��������$k��(m%M�(z�_���`�<�-��T�-(����(4��p��<1���:թك`�T�0q#����]ΐ���
n��0?1^'�p𶥛G}+C��?5�7�Q���"#�����#�\��,�l��G����<ڥ:KM0P��T�B7<�y�e��>�@�9���K����v�y�!��޵�|p��M/�m|����l�QO�o/ح;ht�Kn3^�]�G�W%T5�bA6tr]�ݎ�S�-
0?�Ѿ��I����'��-�#�4�[��W��n	���:YУgOYC	�+|y0dԱ����m�h+���;r�ɐ�Y��?�� ��&�����'k�I��Y~!`�})��g)v�PT�|���),�Pss���`Q��i�)Lh���3�:@J�������u�����fA;q�����)���ւ�B�f��Q�է�q�{6p#�OH8�]ݥaW^�8�+a9T�׆q�E'�#�|U��hr�?�}�:�5��'�E��ǲ6�^�;�1���͎_g��7�J�BI��e���a�|d�جktTB��V������SO�5�����7�t_��=�9��J��S����e�M�&�
RߍD��wU��1�+�E*�=�X��2lL��֬� mB]6���m�*p�?�����7(!� �8�7Vz"e���8�+��9Y�oj˼焾�"�0�k�2K�/��W�C��,ǪP�d�b�hs��Ϛ�R3�
a0A8Nr��_�f��-��G%���p���Z{�_�-�W���Cc����ƪ�D,�(K]�	
�qC7?
I���di����	�8���4�5��h��n�;�Zr��y���e�ZTV�zP��r��P�@r?��������B�X�Ӓ��c��]���ɬ4�� �Wcg�_G���i�~��i���᳂�ř����
M�'Wr�Ƨ�
K	�B���W@:��	V�l��2�f���������r���3l�6���'C�q��p>�7���L��͓��J[���Ĺ�])��6����KB%�7;n[9B�d��ivM��;�ziԄ]�������~��CL�f��u��W���tt|*��C�?#��qV�i\/�U�Ǖu�Q���e&p_\�)�}�X���	;�E�v�Rk4�t(,����Mb{DH�������=��� �~ve��D�J�i�'_ێ�����Ķ�lV۞�^a�˝.��H�����}������T���Y�W�mCr��*�b�M�̥�&�9:i^tJ�~,2�)@��	���sIYM�Z�;�R�@��v����L@y�����tN�[��)���X	w �"T��?�ԉΝ������{^R��Y�ЍvE���P���08��m�~c5xg�{b���2Z��}z߿���V+��;����b���8QN	ew�W@)�b\c���J1�L>bL�9,�Ȃ���{e0D�:si
�naL0AnAY,� `�yX6qm�-A1�@�k1f6TP�V_"�Ύ��*����z�;�8���i�5Ʃ�zs�h#Z!W�_|o!VA����y����B>�6�x�!�42���?C�e��A:A�E;�I4X�'��3�OA�"�/�oQ����:���,t�
i�QyicX�8�����4�3eU�U>��?(<S�w���O3V����$���ɲm���w�n9vU�z TB��ǿ ~E�a���Q����ī�,�l���"Ӳ�
�3Uu��1��9�T���>�b��tJ�["lI���ܼ�U��M�V�ʉq�3dԙ�Q�;��{�o���x��J���4&�]'��g;�����H�'NX��)����f0-�\8[
a����Ե/��7A�-.v���H�p���#H�P-�����b\��'�sR��3�fNl�-��kȕq�o�"|�9���w1k1[6��N%�l�ö�~4~�7�TҤJ�58S㩘Ն�tج<yЂ\8�/o>)���n�:4�C��#}>z�p���r)��_�����)�bX�&�-���lC0�f0�붗�[B�&�g��M�YD��	�������E�3?dO�����YB�Ch��{��qT��`{D��g���._'����P��ţ��L�⭞\M���e�Z�~��9�J�2ܠ�!��r�$�p��͕d�]�U���V	26(�@,�����$p�%����!�NPAU�BQY���M-�=�I�&&�4�d�ֆM�i�8���Ar��>y��-�}H�)(��XO�����=���NiWը"�!� Y �r�H�����3B��ŉG��O��.M��mbQ�z*I�
 ��+D/���<�L��<�D^.i����Vk��A��:+p�!,�ib��R�GP�tq�@�A��tk5V������h�C֠�k���.�]o��/��o�S$)vPQpi�������M���C�����T|� �AT��r�;�a1���z�,!B�j~�ؓ�T����už�б������j9jE_nv3��e�a�Q}��_��C|xп��5��,�0��A�<�$t�� �N]"J������y�&wo��K�wh��$\�N�f���5�L(��Di���A{���<ƥ��𲡸�u��"�B����,�y�.g��S�\�wj1C)f��[�+��\k�y𳧋 _$��[��*'��HT��+X�uW�M�j��f˽�j�������~�Õ�g���y���d��!{�u�����]^�W��;�ߓ+Ơ��`N�n����qo�F�іq)�w�����݃�,��"������|j�ݻKߠ������:h%�B.
8�K����!����~�`��yʇ�r@�[e�cF��2.q��y�0S���}�|��T��)P��j��0�#Ը/�]RUr��b��tm�:�" d#X��>���i�
W��z:&�,h`1����p��L���n��(��.<I�1�P����ɯq[���/0P��Bk)9g&��V����_���͍�	��ZhKs�U;�Θ�q�"�	��9�L�Ő�v�B74�n.HX��0%C�
���ΚN/���5O�QW~��} ˎ�:���c�H�<8��\�7�+p��L�1���D�"U�L��:�e�gTG�.��Vp[�6���b�6ځT�Ө(ۊ#�ҲX�
�3�@����z2�t�M:18ӹ��v��M�wK�eԳ��#� �a��������}����\M62u��x�!����D^��Wן7�Hђ��eM�9�:kt uZ%,T��?=;\�x2|C_Q�Y]�����
`�Z0��߾a��֦��I�ʠ�B�Ъ-D9���~x_X~��y�P;�,k�H��uHI]�]������3��^�Nu�\�6��|ע��B�{��
�ų_��:����w�*t�`�0z9�m�0Q��H�e�n��������pM���U⟷x�K~�K����<�O�r��'�p���%�!Ϙ�����i����oF�h�#��[ʰ��-��uzɛ7ьD�������S@vD�X7���}��:n,�Ŏđ���3�J��2Ф�F	�!*���c���4*,�fGD���6�Į>�0�D(C��9�n)++d:�Ӌ�d��]K�w-���eN���:$,]�x�nWM�~�+����@̠���O"���c�a+fb	���s�\V�ԙ=��v���`���\GP��]"Q�[l�+��)��a���ld-u=�i�\�^H��ݻ_Fc�vBB�W�����8� ���8D~�Bϊt�W�Z.�R� �;�x[��d4���j�n��S;Q<��� g.����J���ZM����\�Z�j;C�C�J� v�u���kM�������Jqg2 ���8�͓��{@&�eq�����u"L����xB
w��Aj��p�{m���cƯ�@����%ص��[�B�8����^�n�m�-ݹ��^S�T0J@����`2����
��t��1Tk�%����)rLJ��꠺ca�[&y�2��Cw(@�S�1��m4/b��w�:if������@íN�O�B����H���?j�~{'ڹ�8��MFp�ѧ^�W+��.����d�=�ݰ�Y��PS��k�Ȓ�����CV�Lk$��SX%P��b%5z��z�e��,�Q����T[b�+�ȩ���3�M9��&R�,�@	0�l��4b�8&�P�eH���N�w�`��~��G��,y:�K���r���#l뚞4>�6��`ѳ�xz�jQ�>3o����:��2����Yȓ�^��e؎u[�����{��[�?�������<d"ӽ��k=�#����5�������ԼF�ءʩr��.<Ik��Vc�L�����4��ϲ�s��R��ZPp7�9���K�n�lr�倷G�-īH�P��m�3V��k��u��E/�rQ�*P���. �ѣ>�>5Ұ0���ez�Ou����6�����$햢d����!�n��b��NO�dxK6�#�zF��\M�aU����v���_l�<��'�� �w~AUXC��"qԧJD��#�K�xS��\M�T�*�_�9�f��a�B���]��9�T��\Ժ��3��8T��L0,����z�s�?�Z�ت��a��;xlhʹ(OvU�=��۷,}�����;D���0Li���7���:y�3��^��aZ9{X��KT���/�~�}��*��]{�O��T�~l���Xu��1{w�g"+Uj1�
P��ǪmG޹�B�����A�|O��Rp� r!�n��P�Jߣ���M@{u�Z�x��p��z�[q���~[�&{��G��K5��h�6��������=;HⒾ�J������)��������^~>���a_2��,�ў0�5��P��j�,�o̪��W����O�@(��-���ZR�W�?D�s���+-�AtF	 �1�-@l�S�Է�	沵�5m�B�&9O(7̻�/��j���z�����t�[� ���|tKz����,{���w޾9Z%���gXv�*�=W���QM�U�/,�@�Fl�z�xW��E�})��.�.�H%>���5\��N�_�(י��6�)B�ɛ�0aP��^��e2؄0��E��h��Z�uei�c/�����y�*[%i��ӥ�~�Y���;�-W�l�<�s�K~�rg�;QP�4͜��-���;��gM@�<�����0r��p�K��B���o��w=~֞&��d3�� ��-K��';���b��	=����2~=� �d�o�ط��q*��-۷IWh�`����cWo�����%��r=�ؙ����W$�h�|�e6���;�W�1_38;<��P��D�I;�dE�<w�_�^!�!=�E�$r'\VC��\�c�e���%#p����qJq�O4�����̕0��<몋兰c�pnA���q.F��&���Z���J���!����9��1K~L��]�GAqw�w������3D~�CK��H�G��������;W�i�����y�����>5�"��,������g
��HD��	���iX.�rI��3-�_)�W���v��� 뙾�Xg�E����\�y�__8�W0���ܢ��yZGs���P����S���o���P����*��U$�?j�� �΅���␲�yw��Ǒ�+Ow�d�Ґ��o��g&qQ�R�pq��U "XUQ���`��!,�4Kb~2ϳ�M@����T�N�|�s�i߹��׳ծ�f����q(�4���j��%D�27)^`6{�.�ίq28~� �4�>�\�Mni�[��si�Ǜ�U<���b��Xt�Ak�X�RT�ES^lЫ�(8<��5�qiʳ�2�����a�+���|�fg/�_�IR�.J�)KX�B��ˌ��X/�-wK�9uux�X��x�(G\�w1(6��i!6�<΁;J�N
gT��m���!��F0���<�3����3C�(s�H�1UL���	ö
��ߙ]�,��k�gp�r*#�P<>�g��_ҳ�`��S�^"�Qδ���G%z?��6�璧��ͭ}��KU	�G�1�̛�`��kL�\�}C��0�+H���֧���$F�~�DQ��~���8-��)k��,��,bB�L�}���lQ-I����Rc&a�a\%�����o��,7Ir���,�(�Q +�&F�y����<��6��*�]�	���{wf.���,_�̐Z[��B��Yґݙ*���j�$1��c����yES�Y���Z��;��#��z-�+�mZ�G1�R�4}�!$q��G�S�ԃ˽�Ѡ��sLePSr�V��y2e�N�f������'S�Γ�b����o�i�#�u,t�=�n�~��?��rQ�o
x��zN�.�Ǆ�}�EA�;�`s��7�#^���\S|E�M`K�g���L�����1��Y�ub gl�LT|��(���W["�5�Z�?{̜u��A	��⃔����#�R �Lk�է�ÚS��c |v�>�g��H]�QW�S��l6�/�M]�0ؗ��t�2��i u<�<;�U��ʆD����<�?36�a��@���}k��j�ܔ4]�g_>kʮ�}R��2֍��z)�ԙ�3$s�
�&p9�C��HШ7�o����^�����](}��BcvR�=�F�F�K'ژu��l/[��
p�JdN��iqgۺ�ow��w��7-���;���1��3�M j|��1�c�gNq��~mwn���,Ѳd��`3�)Ƙ(��T�K����-�#LQq1��k�B��ǎ@n*��2av�ڦ}�mTn��c��f��%�*6Ս�"� ��FƸTQ}��.�Jt|�5�V��"�	�Ņz����T�	@�Ǌ=���*�qف�o��ܒ^�$ǂ����>��g̯*���?�m�<.�R�"�$Y¼��p�R�'�wV�s���E^l_:�9�cϳ�5�`V2P���`0�)�Q�@.�xHbhnJ��IRQ;~�����b�y�IB�煄8�%c���"�s�}퇝2;H�'�Ւ�֭�[\�����p��|�Pl��y1���4��or��0�ɜO*�g�7����V��G��z������;��W����mu)0L���U�eq�ȕ�~��ȝ�g���AC=5=�`j���)n�Y�2�W�K��~�7B����� Gh��;P�G�/kdH�M/^�1�g�6��$?���g��7}��p.~�� ��	���%�߫�.7���{�����U�`t���Zb�!g˧��H�<(����vʻ嶮n�\B��ߓ��I� ��h�`��u�$N\��g�n�����6�嬏����?�E����ص���%��q�mx��  c�E�M�c��g��nE;���C!�:�h�J0Uc���=�&��_՝*A���ܯ�Şh�@.���cС8�.Ι;T��|9/t>��������T`��Ea+�EAjꢖH��~�Ժ*Ʀ���gN*�r��ݻ�&����"u[ች4�����������fK�w��a�q��0Q`8%A�pzy�KQ���%u�Q�G�����z|'A�|�O��݈[��w����"�]eԤ�����j=@[Π|P�ej�Hݯ�@��f8̐�O�ӿs�0T/;%W�1 ����<�K9�LM����C���m�ɓe��K�È
�5�%nq��m��Rj�v�)��b���M����B,$�ǭ��S� L�M�Y�H�a;r59��h�}|6�@C7���W;��:��{�rn��֌
���҆~��0��j��K��z�@8�翖Tṫ��Nc���L�@�>�~j�����{oW�萮�E�+�4�(����Hܞr��l�y�
�cE�x�f�ѠU��T�?�w�#og~9��r�5\�D$H�AM�vNd弛1�c����1՜����q�Ĺɐ~x�H�"#�R�
4ǲ�(A��j�&�x��Øz.P)�Ŏ���7��.�L�y1*�'l�pW�:U��*�eȩ�	_d}�R&+���'�0���]�j�ޡ��N� J���Sn�����[�9�W�~��aB;�_�𡚜}  �f��t �Z~=�e��*|G�;��.*�ʯ"8�+���Ќ�����e�AfO���@���@���H�t@��q�Y��6�=�-�װ�k�H�a�ȥZl�uVZ��z"b���v��t@��#SϦ�):�V �`��Uq#�"Z��n[�2jl�_��~�c=!��`'��l��$.��@�@���F`meWZ �*��R�0�gq��b8U�*��*����A;�@� �[ٮ2�����N��[F�f�K�V4�����0Z�C�d�e��X�{������u��'|���/;$;R��@E#�{L�K�|���@n����V�\�$�����q���}S�� U���a�6�wˇǀ/z9w 6���i�2�z%�4�'���$9ff���Cv�饳. ,g��2Q�����Ap��|vKU����F*O]@JEv9�fj�t_����&L�<M��%E��Rf�f!Ӆ�#jĦ��r�q��%�/����b%�u�	̕i����*C�S[	5D?cf
��h0��{��%�~�iaxI�4��U�N;�S�p�+�B.�f:@��g�<u	6Ij�Tt8��]��;��m~�$c�Zl7!�uJa�^Գ�����7�������g7��ݭt=n���v���B�͆UO��;��-��SM�a���C+G�sX�����w����h�7�NTH��ٟ�ӈ��4�r�ym&~�Y�u�_P\g���@X��ܟ(bu?8o������I-L�L��t�J����(���+�uѪ3�=mkEή��K�b�!rAc횪�DgJ�okl�q @Ba�ʥ�z�� ���9�V�Mb����v����N+1w	�%�6�7��/�cÁ����}%�Ŝ���l�a�Ezg����y��� |��!�mm���Nt�B��R�^" �ɠ��%�h�A������Mv~i��#u�4��p��6��<$�/]Nw#�&'1������3|�.�-?����
���V��ms�`{͖�=�p~�	au!�_��!����k�Cf��&�D�ec�,�v�H�@��?t�	X���5]�g"��=
����^'�Q�Y�t`~F	��im��g�w�Z��-56_�����[�wȖ�*��M�+y���ЄM���<8CBY\�\�4~6)��#�^�SM����3~����1������-)	`r�����䴱��������q~͹�Q��؈l_��!�Y��Vo7�'s���>�~�+�P~�kY�_`��w����)�8�ٵ\*��$@y��}���������ʑ�R6a��L��-����G��׉xj&i�q��'���f��&V�7�H�\s� ,7)�lr/�M������3�����/���v��n�w�	�.��g�!#Y,��rQ�Z;1�r�Zɍ����C�)ܿ��jm��X�_/�`�3z/�e%���@Ȗ���x}ayU���"��pI����w��=��^�|���,��P&�`{^O�O����K*� R��5�W�W�g���Lb��Q2���A7��j\(�*�Uf|AS�sχ*����|lYE|8	Q��{�1B
�G����o3bڽ/�p������8��~�mlL4XK;���܃k~����S	�W������+e�������}�͝_�QJY	Di��� Dꡆ��ĎT{u*��ǒ�����7�'�����@��+3��;6�e�(y`ཡt��#Z�����<d�����62�uI�Ŧ��	�G3u�k��2��t���9|�yX���~��@����m�p����}4.s4��]�|
K��{z�K��{�5�����"y)��:��q�7%�c������t��%6��(!y;��dKq��"HH�`�+�|�>%���$!a,��9N
S�|�3�5��:�6�N`[��b��=U��w��Ni�c��E�)���E�X�s\�7-kh�S?vE�>�3�c�=�?�zشqh�Jp��M�Yf
�0����8���F�+���.�Z��t��3GÅP?�jN�7��V��C��W,s���Cc�S�q��E ��K�m �3��2.�{����G�5@id��Ax��qt�K���c��7�E��+F�P��C�A]#�s�zz��?�W%��	�����8w^�Zb�82#�s`����7a9Ű�veY�A�fʤ��F�����i.;��F��91TH[�r�I�_nh�fi~Z���.Yؑ�D)�P�h|g/sܘ�H�շ���-�<4����R� V���	�g����)��+�����}�Q�(6ŉ�öV�1E��	D��җvQ�me�,�3:�}? ��O�~)�âx���/v��C&��W;�r�YZ-���<���ђ��=���u/2�P]&;���(�[����J�qK�y������>��Rԙy�K0���6=�:���>s���6�	�K;��g-#���,U/:���jS5'?�-a,�V����V#q4�	����o����|=��H���c���L�+*_���+���}]]�,�����h%��.�ko��ox�e(1������*��8�,�K&Ò��n���ζ���v��/��ٗ�8�U=���|>=I����'��+��f��b>B\�ԛ��쯏�Hn�-��Z��bj�έZh�ɯ�1*$r�u�,mN�����.p�����$O�/C�x�ְ�0V�P���]
�EE#}����Ύ�����A<c���̣Ҟ�t۩�[���BȂ��{��j�V���>���̬�f�;T"8�:�a�����<���i.�0�q�
�������V/(;�A��{1E+_=T+mG��+����p�頠sЩ::jJ_�@3�*
3�ۯ	��Ӝ�`����$�j��xȞfG���;1�hn�O�'^b��|�>�R�SM?��I�����	Ĭ�;t�%��������3��,`g �^Y�=<�7��ZZE��Z\7�b��=�f45��h�8۞��m ��,^�o����}�+XK|Y�9N�\@�|k*{�OM<�7����Aw[+ޤvc��H�Um���R�~��.��D�����,䷐Ƒ�k���=i��Z��m\��H�EK0��y�����r��d��SQ�P+:��=���1����:�r�e��3��z��g�6,E��#wrQ(�h��=���0!��z�Q寅J����� a�@�5>��7�6L��k5;�],��/��n�Nn�nr�fm�f<I	��ڒ �=w���{��J�A����q�# �P�`��L]FH$������E���`$T�XQr���ҟeݞ�0x�4�g8M|�5�h��ф��69Xb�Y�+����B���!Pe �#�z{}�l�j�����#<��w݅�*V��P��\�Hq���/企�E����p'G�;'�/����l�ݺT���΍�=.���2�/x6Ng5��""����?�������cB�����З��s��p&f�`��e��
��}�S�h�s����g�K�z !F�`��M6`��;�F�� 8�}R���ߠ�-����6��2��2(���ѝ���Ҁ-�Q4a��;c��i�UlĀƷqP��.��6+��=���~���d�䯃�s��5�uL������ڏ�I2տ?�h��1�}0�$y �2�d^^�1(�f�X'��?�'+�Xt⠔���i%J��قE�yM� ԁ+
ˢvן1k��d��Xx[�9䃪V,Yw��&z���,��{��]vWi�����,G�۬Q�L0�ER�1:H�Z`O�ad^Q���/B%��dD���,�[��)�3���Se�p���ċ R#"�����d�i�?8�W�S쨵�"_Ǥph�QMD�Y��,L�Z�����2�	�iJ
i(㒡^����pӶ<���#ú#w��x/���dH��.G�p��w]qF�e���F����b�<
��o��y����3U(r��yQ]���}򠡏�����
�x��^dIhQ�-�ʁ�̉{:]8�Jd��WUq�2 Fq <xqS�gɵ��t�?*繸�rＲ�,�����������@#���Zް�謲����4ҵ��q{�1�) ��+�{�TZi%�ʆa�\e�#n4��(�>�n��i��X�A�'�KϞo1Q%��[޴mA���JM��\;���;����&�r7��BSR͍�&=�����ӑ��vk�Rk��D�¼zK�i��x�bYbD$����C��x��� ڪЬ�d�Y1����w�=�#�gW�"r�7��������y�2�wj@��U��<��!蓤�zL�1�lcJ���Nj�6Mx���v�!!���qǻ���H�&383�~c�5������� �~��.�-�C�.1^��J$8�D���w�^Jg���cGΈ�?���S3�����d�chP�3�P���}+a)��\EaC��QK�}�s�#oz�+7Q�%��=+H��� +�t��T�n��b�9��D�!]9����ԥ����|@*��RJ�mm������3E7ԝhv�y����	�-ƤN0Cī쬊jH�a�X��D�&u���'��BS}q��ߞ"E�Y���eI�Aҳ�U�!"9��� �}(j��z)���R5LD2Fo�?�Zo�j��
�*QBa�d��G�пZ8�3(�^���vdv���-	�mC9^b�!$�ͨ���܄b\VH�S�b�`�<�vS��@$-�%�l���T׈�V����L�	�n���;|�^��pG��"/���[qb)/���x���L1�j�A�B"楑ꪷ��2F�A�n���� t7_�现�ø�%�[9�A?I�ì�@X�����[^m�P.l����?L���f�xm��Q�2��N�0_R{�zʫ���߫�h��Kl8-^�.q���HD�ւ���pƣݹ3$�Ţ�r�L�$аa��1��� �����ߔ���Q�������~)���'Y�xw8�uW��w=U�
�%�Y�X�+hf�]����a��Nߡ_y�YX#}{�ܴ�
�D��bz�}7�����=�5�
1E��Ast��+��W��N�/%pT�E�ޖ�gy��yp��'7CРIlL`��_���(��J�TQ퓏��|w�}�]!`R��	�Μ('���ss������+(���n��X�<����>;���z#\a�m���D���qZw��z��Ѽ�z���Zpxd�����QN��2�^f	�Tع�f��!��iL]vף`�q]hZ��)�T��
?��Z�P�j��z�Iٌ�_���Gf���2d2yS⁽���)Ͷ���T�5�|L@����9�h/�xD�!��9�I�
�%�Nt�Z���dM圕�W��5l��r�O��l���K'�c����6�T�Og�%�G���2RdPNq�ݥ�T޾ylj�������RB4�,�
�݊+��5۱�;�T����i4z�G����/F��X]���O;�U��R�p�/�&P��vvw�s}���j��řt_�m�`�B���D�@ּ�h�`�2D�2��)}�!\qx��Tp_�P����&9D35FN裄cF�x�f�pE��@x��0�b|��vS �{:��FV���]��J�b6e� 2�O8�-��X�F����9r�Of!6���<gp�x+$���r�xO�AwtʤN5o���G�d��f��ґ��\(�RT���E��	a]�<���rr��Yc~�_��;1s���7h�bIR�%���R�3�d%6�t 6ˑX�{��`9_*t����q�	�<����>$���^cߥ�bz����@,�6���,MU-�p
�����'@fﯚ�B��6��=�dh��l�)$Tx^�uw�K珸�:K��۔��6p�9�O�Qh�52xF�}�s`��t�͏��o4ϊh���&��޻�_�yu}�<��h��CŔΜ^߷��h��mW
t�xԽx"v�QI٠�����yF2���,R��(�]Ee�ڬ�M31���g���]��/ɨ�q\����%�X@���݋�V�n=��:u�$�d���詨`��7ۇGݹ! z���!����e�|��u�]�IY��`�ցd��"����ٮ#7�H���
�mwݫF�lQ�-QO���h�=�8��T�g&ʵ؄)��^?�0�tP��l���/Q���/��6�{A�������'�F?��|����Ӑ���{�Y��قD�0i�5��z��l�#��ꪃ��? �(�܌�\3���e����9���m�αei�f��a;���r�vz�Y3�P�%Ӆ,��1yq�dF1c��Sݫy�,)�.��N�@����i��9B�E N���nqv(O!g�5��?afT�sL��E�^)
�M���ŴtYP���+4��z�'���offq���3��#[b�TQk��˔<^t�	��C��6�����|hqP�8���B��u�jw��fÉ�����c�ou�񈩒�4��5D^���$�<����#�h������O�7z���YI1��R�E�;q�%rM�,_�Q~��]a�ʐ��@�{��V8�<-�oe}_ ��8�E�,V1��{[�u�L��ƎD)js�>V&��*�`4�*����� �/LlQf�4����l��|�(���a���)�bu񡏝��hh�6��=y�fw��M�P	i\$A�#�z�-���Gs�d�����j!��O����6��W�Lp;����:J��O�B_��R���{��Z�fG.���8���|��빌s`%��fA�M��n��	�$�P|mSY7Ѣ ��|�1T�������U��ʱ�x�U�S<ż]�����1��w���"�DXn��X�s9��&�"�8�$jpk����ZE��Nt��^R;�S<���`�`\˭�"�-D�Y�?��]�\rt�}9��\)���o|E���?X�_����r21�c#�񑳨L<{�Z�E�^d��So&U������ix�����r�h,�ےh�=���(u7D�0�E�,�?�I��r��8�Y�[>�m7xV���wx�y�@��c�H{�\H��N�!�"M]�cm�]�>}	�����/l�KL�Z��C��h�-��艣��� ����ڨ
���}D�=6Z�bUD}�Сt����C��o�,n�������p�#��>r%i{�r����zs�5r,~��L���{ؐ�~:���9�Ѷ��	����ck�'�ezq^B��h�����*Xf�K߅>fG�}��$��d`�`O16�K����^<N~�<d*�ݺ���`�Y�U7�Tt��Lz�0�����RW��}�orꌢL�",����D�O�[
���#Fxг�q�@�	���X(|e�����Xbވ5K�8�R�FN��ILxL�:l@����y�� X~a8�?0��Juۀ���,�A (\�|~p����:d��w����[W7��o�*בmr���P����?$���:y=��t�T��Ս���/�ƿ���%j��:H��w K��^��ѫz>���0b˝ 	���D>�cs��~By����G���؎��x�O��L�2���>�,>H�M�<�3u����1id9�q�v����`yH�P^�����>aa��/��_,����-v1T���mC	�8O����ߐRP_3i��T�QM�aa�
�Ɵ+�d�]��v\��������5��n�j4��h>�3q!�3Xx��p�Ӿ2Ǳ�L0������-�~�y�>��v��HD�%���m�XnV#�?���ڳ�_+�!�7N4�$�G�,ԫ�|��i�Ի���b�5�m4 mB�gf����S��/j呂p��7�ͺ}5���&V���)�G�,g�0=D�c�Ŭ����`����1�1�����o��m�qś��! ���Z�����Y�����Ó�᥵�T���򆖳g��-���E��s˭X�E�Mx��Tu�>w��p�L@@A`�|8�Cj��m/��
��G,�[���@qPQZB���z�T���o�A��H|�2=P�;x�Y�-�\U����5��' *���Ś2������=�1�v�Ȩ<Bn�u*Ԑ|�*�����$�z�Rf�/�,]���\���q�<e��L���fj�����F�Gg���x{H���79l��͊���ֻXEI[KzK���]�b��K/�@�J�uאh{�$����*Z�ILq���)G��@2�����s�n+�r���\�\���C\�o��T�\�Jĭ�q�<ˇ-#��81�B��]\����!5iM$+��	k&33�ҵ��%G��eU���ا#G²&1�WE��Fw2���5�x��yC�k�BL���?���>U]�$ %_Ɨg�t[mo��Ub��5iW�|kN>��ubB�Ak["����L�AI����VL��3�~Zo���R.ݏ�{�Qy���0Y�1�X6 ��w���JW��2��/�)��2zѤR�0�3@��뽑O*�0(է`�t��ꬥ}����Ĥ���7j���!+�U8�\�M�����2'���W|@�_����U��?;7�R�]DS�|�s�i2�t��dP_2;���@����j+�Bq�6</��(}��Ht
Q�A��4lI0�X"U�<�۲/������͜���96kb���&R���m �	~.m�8�r9b� 4}T��L�L5�M�3X~��v�� �=^��Y��+!ni*.'TN�k&��\�J4e�'��t���u�~�1�F��B�����Yl�LKd��R�z~�F��j��"v�g����Aa�bhEq���&b���K�[%���瞷��H�����f߂\���,�a�����m`�@n�t7E�����%yF{GG�|��r؝�^J�H���X���E[JJe�شL�j��{{���R�	 q�L|��^�ڞ�K�-��W�m�)1���T+G	���S��A|zE��,*Y��vO��0>�Fa`� "a(@�p����}���Cõ��%�K�N(#�@�0p�{HO|a�
Q�j�'�fzչ�	�1���E�ʱ�?C�"?2���R"Az�h��Ř����t1��_U.T���r|�K*��bx�;�N`�]�;+�E�C?����Rj��Z�)�|]cR�\/k��[�p�e�cB��f [D�g�El=/��a5�N���*ݼ�/�F���[����\�|4����]�q�}��^�����؁DdF))���Z+��<^�Aw�S�;@C�w�'�ڈ�xT�j|Dl#׷��~SWL�ƱЕ�5n+XX�Fծ4S�윘O���+�E�NM�;�HS�VL��U��	#�Pu"��س��S6�"&ι���w�}f�b��%֨EE�t
~��4��U��/*c�7ڋa��߆�ׅ��n��'Քz�go��Z���l��;��.f���;B�^��a{Y� ��v�H��h
�]x��$�J�m�/��=��r�9<n�p�j7��i�zWkQJzˋP��~s�]��#`��M��_�O��C�5xQL�6d�2�[��=d��>>� }�.������7��׮�8Հ��4�q�=Yk�TG'�����V>L�./��L�2'��G��FHV�� P��]��v}ނ7�ĸ��@�^���sC�?7�V�OC�P�)|��+_�����*;��>����vS��a�ݸ]�+��z��;��1ܔ-l'���i�ne��r���o���/B���ԒT};��i?��չ�\m�!#k�l����:�\ �!��io�4��V�aJ��)>#܀�M�1�M���H�@����2G�'B6�n�\@�to�7mņ�X\����MQ��#-�$_�� *��0<ܴQWK&��n�4m�P�]@	����/�Y�Y#%��4~7گ�SPz��N�&S���Rc�P�bI�A�]C^�N?f�`,���;�{AGX����4=Y
����CI_*�.���au2R��5pjЁ2P��.{�XlL��2-���):�;(��g���F�)F,�s�_|��&�'�.i'D�&��g���"[(���?Pu���7�KfDK���Y�����W�.�=�Ѱڛ���-1��Y���A�^�����+bm4�P������ȍg�p}p����7�s0��B�}n����F��ɟg �P�y����qy�T�t�e�Ef�̝�2ɯ*X���$ �	"ٝ?��*�G�(�v�6�D�z�@�"��4O��H�i4�	���N������ω
��l�(�	��4#Ub�D_�'p֪�mx�%�" ��i���g��G.,��]�A3��=��;��{v�\�
;sg!�W�F+��^���]&R{o�̘��e��S�e���r-���\sd�tqg���Я\񰆧��G He6��	4|�1옟 �Tg�ޟT��N5��H�L,n|�Q�\�����v���q'�Rl'���>��%��Z��~�y#�\���*�R���"��;���Ld��-�}��)��&���Q���%ߘx_FN��6Ux� �M�&�@o�`���+��8�!���+?唗Rpr1 �	+Y+�jy���A%�5-=[/s)�qp�����7���8+�r��H�����OM���]k�0j��ťl��ӹ`nj(�3�ٵ����S;��D5 {�������*z�{tk%X���H����в_o�U���>N����5�~H�ґ���OOyjr�2�'�&֘�Y+�^��cH��T���ٞ�#�8\A��]W�E6�i�m�
�A��|�v(ښ��Ն�|s\�N�9�6b7�ŗ��nH$��宋=� +z
l	B	�1����A�FP�L2�"��ܥS�t#¢��ȋ������}C}]���ج�6�c�J��U�4X�D]���nS���l��
RTm�<�0�p�]p0K��տ{H�3-3:�&�|��������g�JS�q}�8��n>�,}���� ۨoz���>�s�P��R���**��D� W�|�
}�!�A��=&^D$褈
q4b&���|0�>Y~������{FW#��A� �q4J�g�j�k �8�<��r`���'�z$:>���9���3�g73G��7��^4���< �d����e�z�K1�,���������?X��[�(Ț̂��ջ�(�jJ@����WI¬R��J��B�:�0y�}�lқ=��r���|v2��c����k�=�H*�'��:t��1[i�v˔	��T��~3b�!�Ӌ<�gQg�]er�(,s�m>��2�.\��.}�m�j/����4Q2v�QC8u�vEX�sOYt�����H�ABP`��- U�A�U*�L0ՙ.��']�!u���ɯA.ꄃ^I9�]�29��®����vI�V�%G��X���y���T�<����hh��`�r�����5����>��� �s���٢����lo{�ʌ%����Gzk��@�#�KbL��'�Les����o;�w����7�>��5K+C�=@�}�:�A�s���kS�;=����##S� ��ra��BU���}ݬ�;L�V��=|��Ҋ��E�~����6"��q���ֱ��奨M�	g�z�X�#��K�!b�T�mV����}I;�&�m��i�"��K�^��e'�j�	)��5����]:K�ՔA��\�~%��/d�O��~�P./$��P��*_�Z�`���N�y]]��'���;�J�ڠp��!�@�&�D�
�Տ\�0���BU>�D Ӑ�ndU[fMfYX���u͸D'p���.� <(ub�U���xA+\�u�����r5��i�$
�u<��#���bbtK��Z���m�
��%ү&2|�����s}�T���R�ٞ�ԃ�W���@��j�zB����Tٵe�y�7?��dQ��:�S���5�U�������1���B\/��UQ�M]B~l�>M��{��G�gZ��؀�LzZ�����mz����f�O�Ay��S�RS�_�֍�n�D��u��ة�Y�K�K��h��Q����,���g���2fB�����\Z�yl��hm�@����{�E )f��XU$���q:7��-�&ѫ�= �� ���L�1�F
�w���C"R�#�/r�b"��]��^�S�u�g�d��@5���"bR�<�%�	���s)��g�|{;��h��;ח�+�y&�`jmF����j���{�U"�p:�ԒM�K�sx�� �At�N��R�1���i�m>����c��9��ک �=�S.p����n�p�����k�������v����X�gB=��/n[}?����	�ԄY�벫�y�(������
��x����[>�ѡGY�s��'�OWu�I�`f[�I���V�8�Ş3�1�Kf7cM�Rm�s�y�9wbk�Q �t�O(�V�&��u^*���$�ңr��9 ֆ�R�����C i�n��Ts�s�ݳ����M%#�硪D�Lq�>y✷W^�H!+��t(g^�Ӭѻ��S3��D���|�#+՗���c8Y��s_`��؁��cm���uvs�
���r��!�j��^aJ�� ��j:֩��C��&Հ�N�Ai�]��t��#K�Xt���g��X�4�B�R�`6��J��i��A�O�S���}ޙ�L��7�Xع�*��L˭��̡M�����y���9��y���h	�v;d+��3P	l�ܛO�����,�
��I�ʑm̐07�B���[�# ��+�GGz���)�d�0Q�\��>�$)��5Z�E��+���p�߯Zy�T�k'�rAGT4�����a��ǛK%�#ڽ݂`-s&ڻD��y�p�1 dK��nc�GY��iS��]Y9��pT,���iB�'��"%2��2ʤ]$� �)t��JE���od�����woF�ƀ��g��0���3?�5�3n��g���Q�>e	�c�/w'���Ei��#���a q�ꅻ�v�YiC����DݓH,�\��xq�����l4�CXd�+��+�Y���f|�D�'���v�VC}t�z��
�
�67߈A;�旼&|�\I���@�1��>�P��XiN	E#�_���lF��YT�|��̭�M̊ظ��V7��z�R��q�}�C���H�3�rK�AL�g���7N-̙����uȳ��21G����Xl��G���0(*�!*gٌ���ܲ�&$
�j,�o.PO�� kH�^�G�����Ձ��l@�Z��+��*�d>l��>�Nl@Z����$���r����HT��`�����vO���=�A��a:*�Z��y�Z�P p2P̆sI�%�Ғ��_[�lg��Ѭ-z�6�)��\��I~������'3�$yϋݙ��``e"�N��,z0�Q��~!3p�\����i�u�ǿ��wTs
Vԛ�Q�c���]v|���"g�lvO�71(�o�E+��+���6�^���^��� YGp��՘�=�	/�!'�lUC6�a[�f��L�-V�ow���.�Ds��m�J�4\�����\1���'&�iL���;8����b��17T+�7r����YbF�:	������m���%Ɔws`R��gKm��O'�<ډ�������REn�f4�	)?Ĥ���aЦ=�Za�p�V��K1Q|Ke|�P]G�d�[��֧\��*"N8��*{ 6���A�����G]*�R��Ru'�m����i`�c��U��FZ��i��)98��y�������zj�V����Iջlu���^9o�/�7�c�s�`WkK�|�i/ʙ��})�I� 	���K�s������j��T^�a-�zr����7c�!�qMd΁΅l��$9���LD�N�<�t�~�Ld��� �4�����'���=ٹ%UXl{�ƒ�.� �d�A{���%~�@�Q��[z�#���r畺�%P���+�b�h�y�$���^	/��Kps�M�\{f6�	�q0��T�=:��-�<�Q���hŇ�ғR����i�t�j���a���*�ܗp�k$��%�.�M
6�k>�B��W�z+ ��.>l#�"�j�r81�b���<?1��cb�U����Z(��f/��/ɪ	M���n>�*�Vc$�<��T��љ�.�(̀'����#W�3G4ޛ�>�q�>n��*kiq�\�1 ������BI������蹩�2��0򽬦��a�� �=��l�Ģn*�u��e�n
��_?c:��' uN�呱[R�7����Rþ^G�;�8ا�&cL�v��<�q ���#(uV,j]��7���1�� �B�, ��QWp�BH��H������C��>����J\��Dp�\��M�C��#8�@�[5Iծ��\�X�u�dV����D����m��;խI�wٷ&aS�1���(:�L�ȹǢ�bp�E�k�m�᱀��o O�����z�A���/��� 4~���R�.�䈚���f(n�pL���U�Ƕ�)5f��������|"���]�_`�<�2�!�4�|%I�̪6T����5wߥ��L�&|�j\��A����Z�<��/�J�r�����M:Z��H���nd>}�t������(uO����!����V�%K�4D;�ݒ����p�Ȋ��jw�3�2����hfrA&�J}��<�ʸ�acQ��4��A�pS�C�:��b� ��E��x�L$Rkm_����;M��Es���ϟ���]�7�[Q5��u��!/�m���h ��C�Q{ !�>X��w�L6d��ܛ�W�a����T^R�h��d����I��8��C^v��`�q�ހ��}+8��-�F��e�f�D'�&�2�����R��G�c��H��L�������Q��B��.��(�r{��P6�?� H�T���r�L�M��۶j���R�~z�ϖ��D!R1�����t��R̘�ۋĪx�hĂaÿ����F?�?��	S#��%��h���[��w�N�޳����$d��@$��Z��R��
�lyb�Q�?Kl�i�bo=����-Ky$9Q�+y��u��&��~��?{>���aaƁ;��	�e3��_�]�(������@���~�1��&ښ��F9I���Ѽ�	�i�fAC�K��xe�$͒p ��I�����꜐���~p�d�uia�+��3�K�{],1�\�*�(�:�kh�(�I>�~����g� 2I�ǆ��s�"��ch~�kdS6!�fp�g�٫��$��X^̗�ؤǃq{㎓�|�9@LP�h�q���M\�Ǉ��~{o���5�y[���ə�Z���� �(*��P��FݣH@��QDDH��-0�ú7�%�ڕ�w���d��9���i��)�<C��j���b
M&��d@���74��j�}I�~�D�&���M�{��
���������[�x���+NZ+���Q����wqg�t��ó����h��-ӛ��f�^�Ka���v����Dmjl�����n�|�/��c�ǿI8LO=f��o��.߂)ة���X<�Py{�ݬ���f �l�0�@�\�=x��E|N��Zy����ȸ�{���S����6��q�s���p�Wɕ#�23�CP�L �%�<q�ٮ�����ghF��T��W�hR:�	-��<}I/�"���������� �^�␲09�I4�lc��~[�1��d�p�O�o�W +�:��2[�A���`1����n��v�]���a��!(����~�n�8'n�p��q��@SaI�y��SR�u��
�0�+im��+�*�CXԽ���S��e��;�1_��q<�-�:X�DP!^9�^-!e���� ��b���\l��ę�Zy��&O�e�����ӷkhk���P;�.��8�`��HM�p��2K�x'�3�:��:΀��
PӸҊ�'�z���4~8K�9y6�4�P�J���#/0s1�lI_�Al��.� C��\G�	&Hz�˚���TL|31�ZK���j��5ۑ�lԴ�D�1�͐V�R�^W��zZU׆�J�q�tr+�wӊ�$�ҫ�;zq<wܱ(����Z��]M���Š��b?�{�z-��|
-*�����HԈ) ��A�NU��z�s/:c�/��Kv��#+�`Ƃ"��c*2A:��y �>��u��1ĺ(O�f���a�������+0�𭾜�[D����+JJaļ��PqZ�]�����S	�s���ӯT�U��~}�O��LR(�r��y�_7;����������k%N�!D���vB?�+`��m(L�jP~3���S�?/��eJEV'��q�k^ud�A*�o�0�#�0���Rf⣆��1Lj��
t$Eo�QG���P�yR�@v��I�WI�B��e�A^\��;����8��p4�6�o�N�bT��Ю�M����Ip���qGړ�C�ꌄ�dС@��>�9�����U�8^.$Ւ�zyR�zv�2Kl���o���>
?1��u�$�G
�ݨq��j�$��_/�Aͥ͋��S#��ؓ��l��{�{�i�:be�KV}�;�̑�21��$?Ȍ5�\�$j���A�3�ޠ�t�*�V�~7��J���(�^��~��/s�2���E�x9����h��~�ƅ_���b��	?��N�0W����x���n0��^=﹉A�T�@��.偳�T7;� �M�Љ��>���T/W�l��ÀՏ  ��(�/��|�!=�9��{ ���v9�{���%��P��ǳO��<�67���/���bQM�{At6���{�G���o"��6Jwp2+$S��uK+���"�A*e:OW�-G�m��R����/��@��`ژkv$�e�lSҖP0���ib���Cf��`�s���繖x�SiTf�H��`�ֺo��S+dzq X �QY�Z�{v��˚�@} �����=�$�M�[+a�-n\P�^d���<2:��E!G��u������ q��$���A}frl�wF	�9�K�p��{(���ig��h�F����]�e*v��L8�#�� }\���;&�ٻ ܯ�_ۗf����B�e�U�&���`�u�c>����w�Q���oׅ9^�{����VB~��ţ�j�������5 7Gu�ѻ���.:�̰2�Sy��Z�Y���ԑ�#�� .	d�^����݇��oGP$�pOYx}�x��e�Wk�໴�`R�^o�FS͇
`���<c,�`>���(ݙ�4.\��~�A��Jol���&`�]Տɜ�U�fz�4О��F�[��85��F�{�Q��3/���$H���!W���H�/�&N��4���/���E� ������5��s��!�9�.\Z�~�4�N��>�������$��6%��V�rD�5զ+�GK=]��6���-�@�G����0�і	��~�����a�Q8�a7�ժ�;l��P5�3��9���e����.~��dH�е~N�Pu4�~�����cYߴD��3�E翿�Gm@����J ��N�,�������H���˱��$p�B�/��=��SVzNh�]���B�N L�*͇@$1�'����Y�Y�|�gJ�;5s^�r�h�
f��-BB�d���;��yȫ�Lʁʓ���#�G��
���@>�	�����ۼ�G� �)%���%��x6ܨ�.
�+����}���g(�Uf�՜Ƙ������3�U@��;���B35����W<�#��/��ga+k3a�=���|�}�:�k"�Jц4!�lܚK2L�d փ2�H��͠��%���˺w$RP���5gGyfe�ૼ&�l�	����U��Wa���7B:�abGP�KZ*[d��s[E�䬸̟���:��-چ�呧(H���>B=RF�)l����`x���!v�b���� ^s���Ҏ2�g�~��>oek>|H�@-�oqWju��u�rM�4/z-���Vˢ�ź��� �PV�96����m�*����1��3��e���-TakDbm3e�8���N8�}�G���[���yY�ZiɐKc/T�����'Q�Gݶ�S�tj>�0��������;im�����1٥�T�0�����8��טk��W,Дވ�	���XKZpm��u�@kS� ,�9똏�X4C$���hA�ߪS��m(p�xR�0苐u\��pn�?��c-���g����&�8o�GC������A+��Y���D��|�c!�	��4D��և����cWg n�|蒤��s������Ѐ;�u�c����J���cU����#�كpYRj���3(��0�-�ʙ(C��?H>��̴E���'�`#y�%<�i7/`�ǔ
��\S���M�����+H7vG�a��Wn��2�BS�ŵ*���i(ߞ�o���E��r�>!�<��AK�qE�	�qpg�r�D\ �d��
!��չ��kuHYj!�@1��eǄJ�)�� b�f,��~]�����ȳ�?���Lޔ���9�O�?���M�BMU�2���� n��Or_���렾Ζ�{�����ӟ�����%�ia;�p�1Ƅ��n)$Di���fRp��t�GNt��H�[�܉�zɿ�Y��#*Y���OP��	R>�`�K��	�5#,��)�%���JG��mS�~��z�V�7A��ʞc|a�;����g�dp�(XV�n�ǵ���
�_�!�nX�l��[SS;cFy�y�����^/ ��t;_����#$��X�"����5CnJ�����sr�0���=Ku�3�n�R���V�����	��z�*�Q�9}M���i!����3�1/��{:�Y��?g��i?�/��gY>�������s}�K�z��&���qLFW��X�0�g�K���e�އ*����C�;��
��z9ݓG������`TB����'��V���]�\u��(W�=�;��5�:i HGg�o�+].���8����|�cR�� 'G��*�d;!��U|�E�4�g�IE�]	`�3�G֏4c H��0 �l�d�c0�L���T�m?��`n�� ��)����,�\���I� � �c����%��U.5~� l�عןwZK�Y�8�nVo4]�(6dEe!�y�h̴%�PHnc�2My��rN ���z��Ns�	a�K�P6�H�_o��V�j��� Vmы^�"���Z'Рu�뉀�g;�Q��2��A0��itV݉>������!�����eb0Jբ��o|<�~~SR�h���~��wդ(�8).��T��R_zz����?���MpD�&�>	D�=�\�ḏ5m�:�~�{���L���ࠖ"��Ao83���K�/`rH��ƣy�x��%�S0��s���MHn�-��g+QhSpls B��!��	��o���\4_!f�:m��1{��tk���i!�8�T)莩�"[����Z:���� g�S{�c^��xm�|��fK�ҵ���%�1��\��-�K��c�yc��Z�9A[��|��L��g���Zs���'ԃ�������l���C��(ރ缣��Q������p`�TD���?������yn�?V���?&5��}��r�NB��ݍd͠�>�0�/D�\�5���0�#�)��*{ٯ412�6�!��Y���^t1S@4݉ä� y.֭F7b�G��8�I���Q:"^h��]H��D宵v$���v�#�1�}^��(lU�H?C'�V)H�B���ɒ��Kne?��L;��wHC�e��(�uk5�;ri�����e��&PSN1�����n���od? ĐbU\�ڊ~�O��fZ����c+�i��Q��g@��I�~�gn��Eg��G`�����\V&y�t�j�;�J�U���v���ۅ�³�Plf�Y��=k6�U��q�q0�qg/l�d��_�S��S���ю}��� �B��ћa�en������;>��d�x��M]�
 ���j��$ٌ�GU4z)����:q���T:���c��$y��wt�q>3������]�|�:�PLIN�wB	 W9�o���oF���a�"��^;%�P廯�(�+J�y]��c6�-�R�g����Nt���[�mF���@��S<bzs%��e��"����`�	Amx�FDT
���f�si��h�K|	�
�W�_d�t&Z��Ϸ2ٺ'�-x{�̗�X�BSr^M��pG����_��B�z�(��&�����pͷ��&ف�QT�����Q���Z-�Ƶ�,Y�Rb(�����Q����bz��뱸�ES�4�wJ�2��i�B	�
�8 QC�M^�P�B�B.�;�1��@�(���04^��"@{�3��@/ؗ�u��:�_f��u#��c��3m�A���
��T�J�T��^��&�i�b�vc�ud��9EϾ	%;� ��L�V��|O|��\��Bb���e���pV�tQm�����1qu���{؂Ќ���#
 dW9������є�$x�
�;�`G��w��.��^;�u8+�o���ـ8'~43�9v�{�V{���J���Qeғ%Jf	�9�O�5�����b�-Z7�go(��s�0��{�W�zA8�x�=[��Y�}��k���O��2���v�N��J1�å���`�V֪��}�����,:7C��	�H�^�S�`�����θ��������QCF�rh) 
a���Y$����y�,ؑ/ǲ��p���#���5Lt�Y_�����i�����Bq���x8���êL�J�sE�}3�D�N�i�;r�O��ӣ>rB�t;��<D�Q2�K#э �����`���D�\�9�J��l%��\u�����`\9�i��'�֙�_��֞我��s���P6I���[~F��I�}ք��9������*�	H�[�m�98���S��,"�����N�j�����=��s�=9H�ok����h����p��y��`F%� %�+m��ڠ�کpvyA����\��z��}���\iK�8�Yj���������_r6��ȝ]�Bu���E@_At��#&P�3b�9^�I�(���=*
�@����r�-���5�hHM:ݒ,�v�|�އb��N͚�qS���űٺ>\����i`:@�AO���N�~�VX]Z8��a��fP�\<�����D���k���T�5O7����n����+EM�1ϺZ���y�Ӑ)3���H⒘r	���	�EbA��rP����������B�L�\�+�Y�ϔ�eI���Ք�v�`�,7��N��$/���D�v�?�Q��D��w��Y�����������)����'�����b�j��&`��*��h<��6)l�RLޚq��-�5��0��$6K�� �h�x�$�i������!��1��i��Iʥu<fI����Ea�a��IH�	/RP��<w+�sg�N��ɖ����S�W_��""b�6�(�1zc"�/�Ē�Y'��	BD򉜆-�g`�_5��o_U*�����@OD�~����Ae��n:w�c/�4b@��2���̋�����п�IN2�+h�oyoYmu@�[a-\�M�b��Ǭ��aR8����z�T�^�ܕ��*�͑Y�~�Of �]�~Ľ>�'nj`�����:[N����kg��WH$zզ���+)�#ä�!=��&h-$G8�-��
�@����Qʍ����_X��me"�(�$$����y��]~�U�-*e�y�P.A�|��)s ��q��?�\��WR�zP'2���'-j��(�9)�i	�|"��)і��Pj��$��pc9���$Zy����^|eW?�F��Y�q�f#�J�!!�N:�[0�l���珍��0/�-���>��>v���jP����E'�
O����J\Ő���)�0�lW7��;m}װ-ξP���[�iEw��'F��$��
4����$�����	pD���9��o�p��)���d�Hт�����ƒ ��,Ru��Sjҗ� k�^�so�TW�L�>�M&"f��TY�V4�']RF��z�̹i��5��̣ -��8���~�1ca�82�aVR1K�ú����Q��͋�7�m�p��Aw�Y�&�p�=�	��Ҝ1�
���mĈ�=%$6�&��1��In2����,���I�����i~l��|�,�o7�<��X�K	{@�JP
''�o��	�6+$��lK����!A�{@�0z7tbz�c���ƀEW5aA����e��nu=yl�Gcn.#�H�~�L(�v5�W��{�1����6e��ڞ">����,+8~�����2:�����ˌ�o�S��6�:��Pr��B�Òal�Krn8q�]̯��YTE6�UHu�
��x!��C��t4��*���	��a2���)Db彅�>�����&����i/]�5�o��S'��ޠM�:��3�4~�9�b�f��X�@�X�����'#��U��@50�����f��]�l���j����VF)/�,R�5k��7��Q���� �YT�*�{�ۚ�K��P@m� es�{��o�*s��G[�y_���j��q��7H�wfw����+�g�7���f{��=�jK0��Fϒ�R����	�t��ӅoZ������B<��
�H]#��~	����8�����ϋ)����W������7(� �C$�d}��U��w�C-� $5�,��� ��K��&�B�;_���	�+�
�Ȣ�#��kyG�>"�+��j��� ����0��4�������m���`ⶊ�J�ɠ�����$6}���]��Б[��~��坡�ա��hD���o��>�<sQ���k<��.M�CbE�J*Q�F?�mo&'�6���w��
�8��a�,n�`EY�:x
364�nA��f:V ���ʉ-�i��΁�=�ܩ�4'���ś���ܵ�|��,�u\��f36oj�w�?k�틦����e���E��Qv����#5�_�b�@���_���2��F�94�\k�ee���C%p˴����3:]W`r�{��<�0H���P��p�u����k����A��<.7?%��.���@Ms�x$���`jvs%	�����O������@�X�"G���%8��pQ(��x�k�K��Fc'G�J詹lUY)u��9�-�5�9��jM��=*Ѧl4�S�B�P��I��(����蹢Zp��*J4������W�_ ����V˃Ԛ��SJ�의 �P����AգP߉)���Rt#��o*���T?������z��_Q���SI_.L
�No`�LI��n��<`Q��6ʕlU5��75g�B����]���i��L�g�K[���UPv,U[��\��R�2x�/�t��@N��x��K����t����J=_5Y�EDx�d�b}A}6�qm}�&+h���l����$�>Y#O��b���*��(%f)y��̎*mQR��}xϵ�\�1i�T�D����i�p�,��f{R���=c��6l`J�"��^�~/D#�Њ=հ*PX������!�V�eP��R��c�����E�z��.y�=\L�1HNf��ъ5wZ��!a���2O�*�
�^? �$
J�AA��EnǟΜ�p�$I�Q��R`�A�Le�*��1XSD'��.�?��7�B��n��ܢ^8�;�;�b�{m�jr �L\o�f5k}4}�
Z#}�ݮo,?�;�Ĵ��]�f�|�3q�'��u}6ŏ��5,��o8f�Հ�^u~����WS~���K��)�����i}a�3��V���Ps��c�.���^� �_]T�?�����a�{Yh�����Td��Kz\>����y�u����M�#ԋĺjhU쌁3{b���q&Gqc����� /yN�iF��'I��
]θ
@)���H���eWJ���//z�Ў�Dз�g����C�-�n�B)�&K�n�UJ�[4���ŭ�b�
���ظ>:���n8�>���E�@;����ӾqyX�|�)���Y{�X38�]�����;]��C��R}��[�1���B��yZ]���;��L�	k] "�Hk{L��r�y~����:�˧�ޏHÁ#���קr�BtA���?��P����Ƌ�fP�!׀fD2��!\._#���n�V�V"	��iJw�	nۖ/��Q����uqA��p����bbyŊ��W�C��'b����ls%I��r~�i4�f�,�T-Yx)�b�6S��FD��#F��4�:$�Ɏ޴05���
uH܁7n�x^��C�6�BR:���|F�.J���)��W�67c��"ӒO<�hq����
���d��}�p�/��G>��ZT<ZT���C��a�1_a�SML�����p� ����B?W�F�Rn�?ƌh�U]�������X��¡�����j���fIȈA+R��[����D�alZ�FK����#G�����(�@.�"�'�`G�ys¢�XЁ�It=�Q�{:ϖC��]I@l�n:MąR�	��k$>�t0={&K��t��%�"�n6�@O[���������[y�@s/Ĕ�)(�U��M!�Ecj��H�-��^	�^��է��5�r۠�J��'V�W���Q%CC9�{�Hu;Z L�f��j���~q�{��e��>Swsk��x��8mL,5*y�D�^Ξ�/Z���J��4�Y�M]zCN��)s���;׻af�?Y��CPB����ۍ/U�z`v��_PMA��PE�:2{������l�/Y����t��
=�B�R��e���K�0@���J`�
to�L�kn�Uۡ��B��J��̍O7��nIp��������aBA����@�2dd$�!L�1 б�L��\Ҕx�7���㌞tXFIX�8�e�A�h�ܭ[�F��5��,C� m�J�ʟ���q����$r,��Ǩj�����|�S,����A�^�^ZG�|�>P�_Ô��,hzIL7�#���K��o��~��+�*��E���l�1����f�M�ˮP�0'ٖ�[��LJD����5�8������Mp���iх�����d��,��J�rځ By3F��y5u�nPB���w��m��p��!mA�_EЙVI��Vʬ.���¬(J�4�s�e�
�K�]j���	*ԞB��ej�:=|�خ�
n��u�~Pu`d:��Eٺr�\(��06��y�{��_�%�<pl�a����|Qd���E���6<j _��.�NF�
T�Jގ�O˖l;l�yԬ^@��Xl,1R�"R�P��i� ����Ig�&��q��H�T?՛*�_#��;ЩgdGY=@����׌q[مK�����~�:7�����q(7CH�J6�v3��,j���J1;�K�XV��.�G��uLC �|�^$���k� M�@;�&����z��)�2@:�����crBJ6B�dM�u�X�1°��E��rV���6��obkw�E��+��!�"`#�
\�,`F�R���(�J�D?dd���tg�#�=�H��e@���Q'I綤$�3JA�;���;��ǻ}�w��P=H3>�F�'��Ȕ���f����i����Ar�B"Q4��TH�
Ɵ�.�X%7�TFUҪ��8W��M��5��b`+Y����C��C�m�J߆��^��t�?��=��@@�qD����xm���������x_��;Rg���i����E	\bm��� ��}���:�Q��&�{>��2p3��
<9�}K2��B������������͎ѝ{Ð�Rf�Z�B�8C존Gfk����Laj?�y&*�* ͯ�m��*nF.���
�c�¦���_�EL���l-��DH�n��!D��hGf�$j�Km�"�]�Ip:���^ͺ�٤��%�R�5��]�W|���z5gH��Et҅X���Р�zt����c⣡���$�9ݴy���޵�eK�aٻ1�7�t�!,����\�S.��4���@"�m�@��Ɏ˩��N�=�4�dvD��"��"�%��ӊ[���X���ߘ �|ڟ��Q��iQY�g�,��&h'$���Z��B��Y ���y~�b�h{^Q�*�+$� �'t�{���^��V�Ɋ��jZŮ�Nd��ٞ�Eg(�8w�����.-��y�Ji<2�����B_�� ܣG�!6��4w�$J3��
h!�N��e��׃�Pp��$=t��\����/���Qy��r	�97�>+�1-��=5y�d���W�5@��c#4��(=PV&���'o�w��W��Á��5}��AB�����dK��� ½��'���Q:B:2�is�k|���@k����[�x��^� L�ԄgW�8�߿�z�y"ʑyu�,�;="�£J�-Չ�ל�S�daT�=�gm�kyv<�}a��%���B���=�q�HiF�j���E���%�)��K�<��Q��P��/��2�QG�h��p8*iX�XN�Z:��1X�g�P"[Oe4I�ud'Zo�$�a@o�ސ�YOS���>0� a���+7Ll�f���,��~�!��\+����C���Ue���T�8�Tm�\/*U'�A�XR��gf�]>�l�Kp���#&�^��[��	_@�dd9�.��q�b���!�Rӻ/�)�f���:�/�ģJZ�;�j�A{�Ne��:�/ȇ�����E(Bő����~m IĲ˫s��u�zZXQ4�':D���׸�56�i�`�7ՙ~>�P������b���ȕ�eY���,�܏m.C��05k<N���A�R�c��z��������vtW1�i3V��8%�F�(�Yݑ�2��y�X]8`�~����v�H�5h�
���_�._����o ��!n��ZI��ٌ�W�ɋ"q�]x��^z/�i��*�������45��)���Zp�`�-paR'A��V�p�z%m&�Oξ9xZ�r6 L����WT�8d�C�3��NoМ N��|�?S��Z�K�Ha���p���Ծw�
�U@��s�X-�G��?h��N/g�K�G�˭4��s� w�1�K�[(��a1ԫ?��v��T�"*2��t?S��qU�|���XC������uy�7�U��r�,Z�df%�^J�T`HFt�<Ä	����(v�4�M���u/Yr[�Φ�ڽ�$Q��sH��&9)���V��l4mN�K$�&��
-�X����(Y��U��0���$߻"̬|.�����Q���F_�'*�}���:�t�D�c��C��3�������4\,��5������'�;�v<z�y߳^5H[���u�]L'h-���e䘵���$P��?:�^+������F�7~+N�j�Ϭ��^���L1]OP����^��^O7�j�߳*��Q���oU:�{���!���#��
�b �؇abb��*-��o��Rr[����Q�IH���x���28U�s ��vWgO�˔� S�$��Щ�Y�mI���,���lR��.&G��ӟ�{M�w7c�9��H��/�JK�,}b&9M��-�8>h5�y}utց_Z@%����(��	7?\e���m����x�7���J�}X,��ߞ2d�oѧ�2����0��A�[Ɓۚ�{4XA}P7������)�v,��=!j�~�RD�
�kA6[4��x	�1��
��kqb�D���b-䥋r�c����~�q���D�"w�YXn���>�ɔ�A#���T�[��ut�8���:��{�8���O	�L��D���fδ1H_Х�OR�� 6���ӟPiJ	��s�[��� sD�q?*����	��u�?:2'�TB����&I���00L���w��Mx�N���'z
���z���)|��V��޸����l�E�#(Vr�bө:���X������jOq)�$�:�CLW%�(S�{�]&z��P�V����J~�ۄ�ߣU
vB�X�1��G�C��P'=L��C�缁�%���|ޜ��D�O��O1n�eF@a�W_�2{J�u�ې�5���x��h�a������V��J?��C���ua
�A��`:�h`�H8T�)�ؽܕ�� �
�v�����lP܀TrF'��ƺ����k9�Pd7y��4�zq)6p�
Rf�,�.^��ӄm!�1Z8��J\�vu��R�.ź��Q`lh!��5ل7e��s�Se����JGYr�ٛ���u�5م�'sdr��=�&�c2~)��_Z��qœ�~�ȺpN��(�n����ԛ�`��-AV�|RJ.\�45<�:�} 9�T��nk�w�P���kp0j�B�vV�yS�I+eG���0&�ak�k�K�t������w¶�j��=CM���W��zF�܏EZ�'$lN�ot0&##9@Պo�S�8��� �=hO�Ҙ�H|�Α8IG���Y�Q��M?6?����>��~��I�֘R2�L�fw�aH1�3ݣq��	�����L>.I���.�B��׊���Ƅ�R�K��KT&W����^����=�x��uI�j���ʛ��ۚ�2Ў��*]DuM�k��GQ{��9�a.�φZ�'�m`3����Qe��8��S���V�x����K1H�&�Z�&({��[(+�^J7|�S3�L���(S��u�4�1y���p�Ĉf�)ËT_�;C�/	��о�8���	�,ꮒ�W����ě�8hDy�POobd�a�����P{ҫ|7�\���4���u�|�Y dfT��֟��-�<h\�����O���I���c����+��J߶�n���U���s$q#M���������¬�}�b/�\z�K���I'Xf�ʌћ��OF�z:��W�&��ް�A��ly_�*�<���`��~C���HL�͢��<��t?ϹJ7=�e��] g��N��\�]��*@p@�GR������B$?�Y���� �@Z�o���W��a�m�u(�G<K�|@\vga��a�d{,����[y4���·�X�a��:���р>?����FC/�L�"�~?�;4�/�u�8��
%�ڱ��C��=�H�z���s۽�G�`��:�e8:�@�W� ~�)+���r\-�l�{:�
�x�{��N%Ԏʠ4�%��@�iw�p8�ޏ:q��-O��x�>�Q?������da�F�|�YE�~�{P�3)�|�%+\B����ѧ�#��[��PD=��)D�Vl'�;呍�� 1�*U�rÏ%�^Q�,�Ě2���h��љ&�B�̩��_��J�g���M'���1�]j�̠
�o�25U�L���#�H��3mp��$&��-ml���Gz��5}�km����%hl1�%���s�;J��N�CU�/l�TO,`b��l߰w�r`��|룐X]�0O���\[A��-�g%�L��� �o3oM�F����2��5i��l	��}袞��d?��c�{��Q�xӬ����=}�r��۱!g��=�C��ռj��˳��G���m���h��۹ʀQ3Y2�\&��Z����J�*�d�\	��-3�}�]t�6ܞ��ö��?vj���E�ad�qȡ���Ԍ�d}��gc|p统M"��$�Ǿ ѣ0�:��nw���,a"_7�-J������)VWz�0�*y��p
�
���}*��%��̌3Y5�����8�{4DΟ��vp�rG���z"����������%�
y�_F�y.�G ��}t�'�6�%��:k�Td�
ob^���!��Iv7'6����)�w��(cn�#�|&�I��$ſtc�L�Y?��3�K,�<Ysf�ץf�j�,��SH�^^>�t@���S\�/�*�?<Nћ��I�$e����xN�ݣj�:�[۔X7=�����`�u	���]HV!��U�> V��̚�H8��� ��m��UÜJ�a���mo֑�� ��W�*���%�W��'^W�<r�&
ώ��C߫7��k]�y�8��[��&N$[�&	��pU��^��f���\�=�.^�j�����ɲf��C.�H�3O�����A��Y��d�I���K�Z���A��8���&;�1��[����K���[|1�'�M.J�r�8>�ў� "텤����&B�_��24�� )!�%�"֠E-<�5�~�:_Kn�φXG7d�{�0�
=�մ�������k��yIy� �SpT�x`�~��~r��d�v:�
�'R1h�K؊iכ�PU�O�z�O]���$�K5�ZX9��X���c�!'��w�~�'���	Q�W����^{����?�6-rf��V.�T��T�A=Vs
�2��8b��`�h���V���\Ag"0(��T�E�+�3�8�?V�ڙ����V '.��ESV'ROA����v�����_����%U��5r��Ӟ( �u����7������h秧�-W�!�f*�
�%��)3��kB�.�_�f?}��jx��% �l�"~'��E�译�wItlҡ��J+�
�`CZ)Þ!��Tz�#���<�M\�[��R�r�X�燬B#n �tf�J�`*3���ΰu{-�:���F�r����C�}[b�Oj���_P�<��KZ�E�L�Þ�$�[C�օ������?�>7��f�g�,s����>��:���^��"�F�E�o�R)�]���	�>bvv������w7� ���#�X��q~�wyr|�@��_�>(bв�����1$���-l)�90��D'���0���vD���v߼C�m]�n���w��n#A��	qL��W[U�Ӏob��9��a�Rs�,kI|�X
�y&��_�E�7t�(<HV���2�y����=�@�umS�L$��h�����7�)���BcQ�AC�����4�Rr��4�Y,M_�ci�:j0���~�S��vH�Цt�=���x�	��'Ƌ�E&��7��ɖ��;a�I΁�ZU��p��;��t��1y��rZ�пK�C���m0?,~E����qqV(m�Y(�P&tH�_���=����m�Ř51���=�s�m#����'�S[�1�T���au�gҔ��&\zeS�ۡ-C����_-���R��ه�$���s,U�Tk�9&���-��qy�h�r�R�G���`�$ڌh�<3�qpjؽ��gb���"��$�+��x+1�m?� ��
@�ǥ�OLU���-is��ƁKr6TMZe�S�e�k���5ĩޡ�/'Lڻ����+��*���;/� Ԕ`��[�&���j�VS�YP��7~�¤n^Ë5C��(οC��qa���j�/ �a OyvP��F�y^f��,�Ӧ��Լu���:��-�RL���n#tk<�AҦ؋�}�v�{��½��+��OPW���͓T
�k���k�r�n��3ce�b1���q�r��c�#Z։c ��\��z��~�a��,��o��ȌZ1*�I�w<Z^�ІD���v1�:���J��ߌ�n��odJ�Y����ʡ�v�ל,gB��m�B�G�1��Q������;9�
�G"4�:�s����^���\�˗���h�]z!�V�-���c���#�䮪���hl\���=�Kg���6� ��l5b��L��'�jRؾ�p�2"�c���W� �\��W��BU�=PQ�g�@ir30BsX�t��U�6K�[�ȣA�-�?�����.�f�E��ɔ�g���Hp��v��ò}��?��_t�xy�
�/�W�z�W_�������1F9|��_D0uc&S,Qt�J�@�l S�wt��b��<�����d���j�ib14 �o:�������z���8`�,�f�A��w
�Bc}��>�E$��&N�vm�}��
1Wp-��u�e�g���?���A`��2��5^�Ȟm�c}Dţ��L\]J�ީ��nk�y�[yq� ux���-	i�a���)����oHP�������o�`?�V���~^�p�9��FCpt;�[M�Q�Ξ��L��&ݮ�',�)��ށ�O����l�wW��:|�f�k�:��.X\���?ԛ/U޷M7QR�:���$�j��rZ��
i�.`G�Ж3���.� :N��=�U��6�,F�"��%� i2;�k)3�רg�ʃ��p:����� �#���T���?Z�/�|e]d����^ ۸�rT ��?>m�MU�T�g�N����<�%�t���0�s`7�3?P绲��8;:N��p�uO�GP �)�X�.O���H��r!��<����3���E���#��
3C����+��u����t��s�!��i��#R�D��ɦ���������;h��Y��>e��88��1{"k�E]��4
F��������3��{��托��9y�\L������+��%���Oqdف��������N,>�U�e���qB����K?�F�����xt���"�c�T/��2�cQ�*Xa��<�A��V�%���}YT�D6���K��<�)�u��CZ��;�LHBN�.
IN�XFG��BW����X�3E �C�֯W]���miQMsx�M�õ��r�.�=�s��n^��{�U��%.ʄ���ZgѨ��+���K{�� �*�q�'�,$%�'���>L?I�
��/�xOv����#�{�eZ]�m>F�g��Ha��c:��I�l��k����00!G+�ͨ.ੀ6��^��j�vI�C�aо��ת�,h�֔��2v��:L�-�����$��0���=�2\�3.��'�'��V��r�Q{��U*��u��_����Y��(�zQ�'"^紭w�oѤM�E��H�͠*�H�|J�/'��rX�(��9�Eֿ���?�%��_��\��쁂��q�C���IǧG5_��D`��X�O/[��O�^4�#�]Y�� Z�[F��~�9��I�?8��Б4��7�C�?�,y���T`�=���Q׹�~�L�Q���I9	���*�T�}��6c����:�S�>�@��;�O�S��אTJӑ��?VN���_O�ec֬��c��Ԏ����EH����2�5�y�1�P[���.C@�Glk�rSgy�%���I<�Z�����T��Mh�m=���@$[s�
Q�O��_]`��?P5�vQ��*����H7�`]eUPQ$�lR���޽��Iygm��4��b��m�6�y�~�SC�T����'K�+t�/OIoaªw��l�g�x�K���[T�&��'���.mBkNh� �G��W��TVf�\��̽2}^����-�9C8�b����t*��S!�Y���1���~�>�nɿ�EW�\��'-�8p�x[v�eg�Wa�1m�M�dE�Q�B�%;��UӇ���,�v�����0�p6v�|Ki���4��X�P�#����p:=/��[I�?�Xe;7�e�ta���Q�	BXnP���>*wE/p�?{���j7���v�!	�1�v�QL�A17I��d�7,)�i���V�q�FX<�;�~]�S�خ��=��yⲲ�gda�ӥ��>�S�����y��!z�]�A�B���u.e)��&��~�6�q�JGq�0sC����xu��<1BI2�ҥ<�6���p�����OBm8!�jth�gy��8�o�X�2���x~��-`����iZ��PIf�&����m���݂⩣�O�|j�HҀ��]��wٮ��;��M���������fJ�;ɻe��34T§O���3��}�|H�����9�Ŝu���"�5����U��-F��÷{���R~G�a^��M��D�U���a�aܦu6Rh�:Ri�R�u�,��X���B���,���o6���O�D	34=�7�X�,��1(h]gf�|��=\+���^���+ї��%�O!+V��j&X1��_沜'��2�>�m�~6��|�q� ޹]�X��������ڞR1w����?a/*���Y-�v�����q�@������or ������T´��y����n�@�-�'�ڍ��pɄ"�B߈_�`z�*�����#��l��=#�ñ��P��T����M�V�8<�I����+�\⻇�kfßBj��!�{��T:�]C��MJǑ$b�"jx>����N(Ml����H:'��~����;/}����C�w�^�HxY�s��f�PB�r:S�&�ok��x�Q5��V_�g�GNơ]�z��]t���<�؎b����cݒ�>(5c6��dr;�a�$����w�'Oy��iF�:���5+��'�Ų�)��#�_Q	��6d&u��W.��}]JQ��u&W��7+��9�ϔ%��b�Ðr��$a^��M�|��Y�D��~���+�l"�BF��8\ۓa���Z5��ӌQs�/(��p�`ZG�R?y<1mJ�P�m�l�F�[XCa��V�(��<�w
�K������Ӽ�XL���҅8U�ִ�C�n[��5��l�t��� iIm�������P������ŕ�¦[�1�0� �UI��L�<3���9�֬��ϰ��tٚ�%�\Ņn����/��q* ��{�/ҡ�h�I��q�B;�f�-ĜVz���:���(%A������3��ݝ��n8o�è.�ܝ�y>F�⩝o�J�I<��ؒ4S�O=���+H�L ���ڬ.�W#�����pi�`	�?C�*4��5�9����U�;V����i2#�l$��UBq�*���n��7 ��Z���xx�:�&��I�N�n��i��er���m�Td�hOS�� h�T1��xF�*�tf ӂ5�����^i�f�2c�A$/b���,|;�d��L1k��LqS��֫�C��C`�46n���n=���];l��4,�ƨU�iq��7h'�@�����B���-f`Oҳe?3��i��c<�-s���4I�2����.w��[e#~f<|>�z
c�1l�jP]'��4M��_�1�{�r��.)4U��m��,Z��\��γ,�C��=?�p�2��<��PGN >�s�^aQIT���0�q3������v*7Y��!�#n�����ɛA2-|��LM��~G�	�!EN�r `	�w�
$�l�ȝ�!����2����(@oz�i��xH;0��"�WSI��ͷm�����v~���F�_>:����u�ռZ�M�_�>�ng�rtw|sr����gzϋ�����Zq�-N1�&X�0������rX���դwX�����V>��>E���ia$\�Yy�̺j_�	�i�Z�Q�{}������߉�Le��jT�Xe�C��IOj� ��%��b�1�A� ����]b#i�Y4�	���c"Oy%�0X�F��S]�\lE�d�.T%������Vn&�X�����7q�[���ጀ�_�ϸ�>ۀ����`�����qTh?r-�	�)kzS&�#����c�6�9��z���K�^�G'�nw�>)zI<t��t��>���Q��
���r�M���(J�r��}�*O�&�Xu)Y�H����UQ�t`�c�Q�"�{>�X�R�F�Wcvڢd�Z�i���!�?Q�͗cT�S��C����ޯ�@p�ȜIGV��ǿ�#Ĺ���v�>��c�ڻ�'��U�dݸS˸�/G�c2�z��ʖN#a��f���"�Icv#��An��R��:��:�\E�md̎����/�y�2��8�ʱ2��*���v�������4�E�wIa4� *U�����k�Ȫ��'ے)�"��O�NrW3n(������d�K���Z�r����Zڰ���Zm�4��}���h�b�&��ʛ?I�.���潇p��ľ.4MM ٷ�>D}1�X��aNT�"5^�O���l�X�p�v;����+��0*�H�Xq>�R��V� �E;] ��Ӛo��+�3������a ��+/gB��������&�5>R+Y�Ъ��m��,�z��T����@�V}�w��a�B�n�w(P-�����G�ec����1蜁+/}8��A���ڝ����Ֆ�ײ&�nǭ�"YW�����(�,���ZfCm��L���dx��.�ӥ�����u�s{���+oȊ���j�w��9�2�g�R'@��fs>7������$�'ه����N��@�M��؛��8��r3�dU��A�1TP�jA�qWt�T�~�m���e�zT�mV#R-�\Lt�[�dZ�����5��e'��W�6�~:���g>�L��nML'�ƹ>�bu%[#i&�~���%����?P��K8���ޢ�0_��u<h��Q��x�.��Ye�b����"�c����	c��u3�*V���%z,�y2�Kͨ_�f����	��s
�LI��^ZUF�]�%p�@�3F 0
��A������K������o�Q�/L`���Tx�-��d��O �`׆!�^����n,S��\�%v!sZv��"�I�u,��w��;�{<��Θ�P�>̋Ԟ=V9���P���6�c\S,��^^�튚�8~l�D>�;�z��}����u�� ��3�)�������c#4���D^��%�u��X�+]fs=��<@� J�
ц���
sڶ~�?~҉[��l^��͟RKe10�bg���av���ܦ���-�)���.�[o�N��Q��%��� $Y<��s��F"�G�c&�O���W�z������J�p�[�24�����/�t>���Omq��f��o�eM�a��̕G������
�z^�[�p;ln?��`���OvK̼��CQ�ɇ�h���G����ń��Y��+A&`V�Fv�lh��t�m��=)��t��s�%���C���U��������JR����$�m·X�q�+���{�8�Ԉ�啕B��~��ݣ��[	ZPf�h��,�$d~ӄnV.�Y���q�n����:��4���om�
��(h=�X1Ԁ��\�����?�u�Wt���OZ�
��ߓ��u�V{X�#��?V�!#9(��y�ܣS}����V�b9�����;� #�UQ�)W^�����"��F��]��Ɉ�ed��������v*�w]�H!�F�k�P���pܡ당EHghJz��^n��Cmp�����ܜv񣝨ZP��������:�QaC��2{jfo�w�3S����l�{o]��yJ� _$j��뜓�1�SX���Z�f$�I�a�o�-����>'���~j��~ƹhé�m�u�b����$�(S�%�5���@a�I�������VD��4� Ag�GƠl�\Û����F@Ȍ,�Aw8����!��`�<�[#�����w$wt!m@S�k�ms�n;ߝw��|�/9�̕v�T�K�.�9��e�J
aWp���F�����[`�4�I���X{ޥ횊4��8̾V�c|}ڂ����,�]m�˴�4��'�RbRY^f������&��S_;�*��a�Y��!��qL�y��̶���+-$h�~�I_nM�R�۱8���ԙ��`�0� Q4�]ɷ�SGC� _8g��H*�I{L�;�4�6�d���m��O���X�W�œA�)��#��uK��#��2B�z� >�\�yTQf��=P�7?����&�c�3�!_J����*�x}�@�v!�����v`��#Ը��J����)�s����jU�#��m�P8�i�U$��j(U���VE`����`���.��.�s�gz�{���]�iL�����dOD����Dm��������Ĵj��h��>x�`��ǩ�@"�Y�d�⅓,��4Mx���� �$0�Ly@Z?�($㟎W�jϤd�9ل�s�b�i�B$���ٗa2��Y_Â�-���x����l����8㕓[g�B+ku�ũV�3E5[!��!�/����� W�Z[�#�-3.,�9�F� $�*&e�Ty�m��[�Ph7[��H*yFHš6�Hv����b��VڤfOp��ٓ2��~)w�K,��"�h��	�s�Z�Ci�����߫�����Y�h����d��*�N)�I�"�_Y�9q-�X� ���G;�9v��屣��5�����,��h;���|���n��g��
06C���}���`�A�l�_S"C�0J�Θn��,D��:ocQJ��gd1�0�(/zO?��>
�;���W,wP"n򫚵���	���đ�>��f|֜�:ʢΊ��lSuh�8��x+�Dޔ;�)��%��iS�.��Zm�/%���y���mr_+��`RE��w�o���3�X�����v&}(>����[B���}��M�C/�%���o��Km}z4B�?�����(�9[�#L&�z ��Rx�5��Y�_�	-�,�!��%kQ|��.�Z1��W�����������a������^�l�=58qSB����
1E���'��EF�Xae�E�{|�6(,�>@V���<�GPб��[��~��w�k~�S�� �^�������k)��*���4\S��T�]!�(��7���(�����f����۰�+�Ƭ�\�Z���G��P&�Y�įч�d�|I�͊8�p���N_�)s�i���=v@:O��UI�*���B"�wP�ۜ��8�v1'#M;n�	V%H�m�~f)�t���0k1�������"�]�D�&�	Mb�M�`U��3ʑ�jG��Ud_�-�g�0���m�]���C�,֕{>Q�~�w���LM��YFS�F,i�/�6��S��8�욫��;��Z�LHSƽj�����֬w���#y"�n!���:}=4�O�����ᶀZ3;:���G���UJ;2p���.���V�m��K��nO����;�p���^
��_��N�¡}��P�`}�xƖ��։ZW�����P#�\�u���oE�l�I)��(��š�NqI���}Y�Ң�6�8y4���\��7&l8,~���C� �6]P���]���	��1{�־�t��n,9� 2�ݶ��!�͆���4-�0'>/̷�\L1��$N�g�}$h�T�!�F;��q��
I��~5,�R�7_D� �(�a���(E`K�5��`m}���9�2E*O�w͘�yPs^�l��|��pk�V�i5��ϴ۹�3)ntW��@.-h�Ǫ N�=�YW���VP~�����o}��&J6�Pi߶)%�Eē��k�b3�6�n�����J ����
����^�D���Q+OJX������ңjT���p���4���*k)�	pG����w[#�f2Om1$���!������C����b�6���*h܀�ҵw'���T�~������$+Y&kг�N����*^�	jb�MbE_�I�6s*ؤ��ǆ�H��5�&�/�vm���k!�����0h̟O�^�b������<O]�ѭo��Ҥȓ��ue����~�`�h�Ԧ�\�if\c*��Z=$��){U��|}z�D���Ӭ1X����b��⡮�B�~-�0���$�s����9�-~x�2�#ui��KA�^�Tj��ؿ���q����]�������ŀ�v��+���:�����SAT��_�����yj�GZ��Y��b[����J�s$�`h�B�y@O�Y�)O�5#�'�#!(��,�|R=P�ϰ����D�U�����>�jwP�c	HW�!� BJ>$!��)�D�6�(U%��M�M��}�\2�5�3�wU��!ि���*uC�n��	���*u���V�e�W�Z�A����_�n�|y�'���*��R+���!��$H�&�˓gթc��$`���<D�	�>�@�<�N҈����ܹY�=�X�o�x��l��v�(�"Ү�p���T���w��7%Ő�q�A���W)�xn��*k
��FZM�]����] ⫦%:��	+)��4�\mQ�NS��uG��d�=]�1o��6yP���m��& IpC�5�?;��0'�����X+�js�N9�,�=�O{-5�,]2�
�͢�u�e��_���ɫ2F~t��΋n�AE�;�����4b�U��pHr2��^��۳�'�9K�\�LԵ�d�Av��+Ll��;�<D�X_h��z���2*�d�����A�䪈������7/l�����h�z �E[�87Q�v�����2_�3��<�{[b�-��2$]�G"���!ʪ��#�VD��oE�#�D
<�0����|��y0ӥP����/�U+�r��1��t�<��|Դ�Җ�৭{�p� !_��nR�O`��{U^�x�}�л6��YV� l���܀�'@�<��f���1��+�P|��Z+so^v��#�s�T�rk�	�GoE ���P6^ŵb_�t]'�sW(1e6aw��lU�'��.�x&;�!��%HL�+�ۆ��������i������	�Zf�e6����W���y�MMmz�8�A&?7���r�n��8�����>K��G�q페��ߪ��5���ݨ��I�^����p���m�A;?[Qj��e�B�k�.���/W}_��_4��a�/C�b��/�6`C}�}R 0M���{�*�!rW$]�H.��P��yG�.+��'L��q7��E��]��)��-I�E���}�ဌ�浍u��5>��h*�TA��u�\���<I�u��k��M�l�o0�.D��0��
?���V�Ƭ�}HdS����N�;�h2�bĹ��F�2�Q���M�Y�������8\�%�<N#'��v�7)^@3�Y@�;K�����vDV.�UA	���V�C�U	F�d �b����?���'��*����kC�c��d���ni&��y
I@��\ϔ��?P̸g~�RF[*&�E�$Ѷ=�sX������5�UE� �Z�u��P���sh�����'�yܿ�A�À���� #���i�!��S�A�ZI䨦+b��	�&5���Iewp8!�9�R�i/1?�*\+y�MVCB{@��D����t�-��Up��Ŧ7K��kh���]��� �R$�3�:E��c�u������˙�𳖯G���&���?�� K�k��!y%l99JY$e��e&�`����ڰ��}���n;�~S.Is�&�;�����o �����`8�����`� #�V�?�k�p	���I'�<��4��J�\!⫒S���pHp��.� ��u�q2�H�K`�,�8H�AX~ԳUL~^����$5Jޝ�y<r��SpE�ĩ�?� ��PH����븃9�/<(�ՠ�n�tā���r�e��"�uJ�F���Q	3�4�	�fX�Iz4�IT�h�LER�r�^�l�	�"+�wď^�yB�u+�<�F�dC[��'�[����.nJM� O1�v��+ba�I�$L��B�+���H+�G�L??]��V�H��.�Ś��Xn}��H�b����U ���FA��p?�>����!���	�'�J�$vB��R~m�W�u��r	�w���s@h�b�ʹ]T{1i����]R`�~:�
����F�]�F�c�2Fw�;Ȗ�m����j���3R�o�΁2$�X��;���C�	i�_����o��˩hO�9��>ri�Ԛ�A�b�!Ҝ ��?�y�?_S����DM!̱�����|���p�Q6�Q�L4���k*~����ߺ���sC�x�v!u�4Y�'s
딁uj�����*�]Ʋ�C���e�.�=u���;P2��AV���Y����rW�/_��c�u�U��V����:��;�r�H�SDiI�Y���,�~2�$�[֏Sy 	�J� qj}\P�F�<ߙE����TV��"�r�dH&ې��U��=D�]E��_�8I��ƕ��t�8��Ker��#������.�܉��Pd7��ܵg���PI1��]�X+(��A�����[n/����<$��m��@o�Vnn���c��SX��M���P_���/��>'7%�!�w�O0�֬Gɦ��|�1����z�R��X�>���C��J��*�c��bO7O$ ���H�Qأ�H؃<�p?��6�3��`.w�����`�fn��D�5`��	��-J�C�'�J�����CYw]�鲸.��	Y���3R�v���+�Ւ�Q΍)r��{��Kܖ��ё��`韌mշ���w�?�-6��U�P�c���ߖ`>4/�͊Љ�a��˷�4�� 1)A9L[��^���Ypi��,�CK������T���eޡ��zlr�7";��*���'�;��k��Ho��^�[�Č�S$�nH�;N,�(ʹFf���&o��82)�yrx\L�����Q#N�-Ys�6��;��;.�s�b�T����s�~���ɂ:"ک��(��&��_<1�{��F�s�gí4]އ�"`d�]z���	����w�8�O%�bى��hV���W P������-��Ŕ���FG<��&"l�tG��՗/bq�f9�鲆˚$���J4�V�e<�� �A�lK�_�RuZvU׵E^\�7�(gx�պ�y���qh�HҴ�<�����>~]��5�qϺOܥ�4]���	M촷�$�e�8~=���Ay��pz�16<~3�W�U�k��Ǡ�G��厅ё�T�Ahç�E�F��]4{D`RRԏ�w$�C��ֻq���bk��G�O39`�W����Š��*�|?l}��Ū��o=�z�T4�!��� ^�~	;���}gm}�r�D����$M4?+�x+C>�7c<�M�>���v�g����_b��ٱ#���NO�;f�3"�$�&@��n#����R��D�=4}��c�P��-vx�XDTp��L�4!'e����.���\5�+	(-��9�r�(氚n�.��W�l��/M��1���'�:ţK��T�>�j�n�ϊ���LBN�,(��B$����Z��t�=	�<\���#^V9Ø�݋��j�֍�}`d�*���#��8�2�L���pp�n8�=6��d]
�ĉb�ox2Ö$���2��^�{�D��/R&n�W�Q��A%�-���?R�6�ˉCd�%��+�D�5���˙a������U"�/�n8�t!�zE� T������V�@�:�o�b�Y�#J-��ڗ��t��JV�����:�� m{6pK�<C�����t�?����*����Ǐ3r�d���̿�N)uSA����'��}yZ'ׅ�	�
K�M��Vw��ku�ǿH�{�������G��z�6���l��Ӳ|g6&)��"��";'oHw=�܀�i|po����]�.,e����څ� �º���'o��^J���7����1���I��׶+�����mqH|o��I�����l(�;ӸAx�f_0�C� ���A'����v{�Mf�\���"�����A7�BD:����
%֗���V߫���\Ι$?ƹ�}��Huָ����
� "E����,:�T�S��s�1N�%��傞��[y��%r,w�l�X�|4��f��n�ϸ����U\��	������5"�@��)��S)':([�����ǫ]�ڨ2#X��q�g"E��$�7�� ��|bp�݇�9BE�!Z��$,��:fM_�̕10��\��0w���v��O���EwJEN6��	՝�R�\�������P��������Z���P�m� hy�[�7T7��|�oY������Y �2E��o��M�"l{t6,:w���E�9��Q��ʡ�Meɜ�{sA�7��pA��[�e�0ߡH��B��;o�p��lxɧ:��̍w̵�K9(@�ʮ��;93�4b��=�k�����WY�&�7��>^�OF]��f��wK35
����@�Kޢ�����c�C�a@�w3Ɵ�W,��@-N�(�91�S�O��Zڡ	LжI��<�����@���\v����o[?��m�'�1��\%��WB�3 �>��^J��5��R&�l;�GET�;%&�A]�6э���RI{�x�X�u���.C�#@	���-a��������Gc�~���A'x��k9+��>Z�`�7:!���+�" ���#���}"�����1R��ϒiY��h��N�b�l(��'(C�S#z��)�Ц-��o.¹2E~v��BY%d���?H���?\jZ���b+��@3��i�+���ɀ�.?��F��H�=]������AY����0����Z��哊�3��x��w`IȸVZN}�r�h|�IU��u�^?8����:�LY-`�)�Yu��hO&On �^�PF�=�e�2��b6�l�P��B3#�	�E8����|�;[���CPdvxn���N2��ُ��_����h�<⏍QS�=[��q)f�FX�C����t`D�ڿN\�T����Qw9��W�-�(�v?Zn�o�i���p_��R�����n�B��R�yA�<?�yc��Blc��H�5Tx���j_8�[�P�PZY�B*�͠�:��)����A��P�P}J}�IQT#�CH�;�5(?�S_��3L  s���cqC�)�M;�E�t@�崏�n��K]�l[���T�FI��`p��I�
�9�`};�z�-�>�"�6��0t�r�j�Rd%���7v.TČE=q�4)���xe���^h���#c��{I }�u�/������/�pC��Й��$��*0����D~s��h���U�C���/G ����O����%0�h�?ZY0�������'v��d%x�~'=�э�\^��t2�/�kُe�Pg酩|:ǔ��ZJ���Yۑ�μ)-�,i�����M�|�͟�ȝ���>��t��=le�����2�a�SQ�J����*��ܴt-_ZZ,ŹZ8J�((��Ť���&�е>Ċv���(�� ��eO�f�t� `�x/��w�����w3�c��$��o�:�|wDe��d�Ga)RI��}<�y�
B-P����=��m���@A5��-�����n�ttd�=����Q��S9��!�0A�X���"~a_x:Т���u�_��nn�-q��v���7V?�k���sᆉw,\�؟5�Hs���s��JG��δ功}k�kZnUl~)��Y�s���l��KX-R(ՃT&ц�sT�:�6�v�	)�-����t��1��i'�	���2�3V�=$>��B�)�)>{�hـ�F��)�4������i���!�(�(����2�3�kv�e4����È��v�~k[��	��`�5�XZ�32�$Ue�Q��Z#s��|&[�i��E��� m����]]n�42��J󲹮4 v��DHoR�I�7�%v�@�����D~�������E�	�rʷ����O (u43y���:���U6[*@kDc��u����m�Ig���v��W�,��1&� ��A���������Β�E>��>,����K��xG��C�`��ol��^����(��������˭�ˉ����d�?G���(^ �ۣq�G|�3�B�b[�_\�Գ}Qg�^&+G�Q��oo����A���6�O����:�:$�)�'�Xb1��[o !ͥ$D�4�P96�t_�0^���|��H|��o��.��Jx���d*{�Z�VfA��C��fP����پV��1�ar�=�-��?�P>mh�L�:�*���K��r���i�6\Bt��]'}��ls�z�5iN�}t��6@~�V��Y�U'o��b��X��Jj����7��[=e���1�"�ә K3=̈́ͬ�۴��,6)�Z��#�Ս��w _�=���WҔ����2���o@�@�^�&��k��y#�f߈6ɸ	H�����V�U�HL�ƭ��;���uO�B	^%�fR��Bʥ{�7��zRu��t��0�w+��[�����=]�z�W+�QP�v�=�ڏ�~s+x�GM����B�:Č�,Mt�>�a��� ��.]B-"g�=�:�XUyҤ�c��X�M��m���xf4�W��Zn/!(��}X�
�zK^���"�5L�@n�ɀ������	��C�萝d��W�^<��h��z]&�i@�� j�~$#K� �����~�်��Ўπ�)qB�`ӎl�h	���LO��}�Dk�j�eq�+�d��4��d
�h{R�ei�|��.�R�fq�\�|o��XkE�����ה�Dq�t�Tk�P5��a��W
��p_"��gg�М���˾]����hj̠E{���=y ��`UFC���%�b�eZ��}pA�����K	���|='�]r����i��? �.��ި;-la�ܿ�
|�<M���l,% 8"����G<�|T则5a�3�_߿�R�r1W.Y�ɇ���N�Ya=�L�e�K��Yլv��T�:I����n�0=�6�\yW$�Mz�@��
���;�m&���隲]��N��h_"J��Ы����i?��HpyV��)Ŭ�"�	���,}�|'] ����N�QZG5��	���]�}��� �F��D�L�s�I��"fGO��3aL��r�F�,( �v�����P�^ӯ�]�pmJ\��9'��ˍ��f�Et��������X�֩tH���
t����@�=T�|�����:����/�rZcLH��q}��<����������[E~*�-فX�^�5��N�Х@Fq��������6���C�\d���6�B�'Dc,7��++�a���O�.8��Jo,�EZ�/r<@#H,�t��B}'*�S�EZ����K���6�n:88hХ���6��O&�O6iHȪk+�@p�1����D�*�8�imfJQ�����/��6-�\��V�V�S޺��l��&��C�Xx�}��1?bg;�=�"	B^�Qq�2�i�Ҝ�݊���Fe����^-���pS����|"�S�i.�8�l-��Kv�e)�`��+U�S�]��N����T��G���?�֥lM��\9�?��H�k����X�E3/��}Q�����h�P8�V�{$�����Y�ߕ���C�Mo�	<����Bf�5��"�)�K�Z��9GC��ÏM.�6��QqHDc_�7����w��{r�0<�Ќڲ-jﲄeO's�})��Y�etq�6���A�x�b4"z/h�"�oۡ����-�2�s�����Eg�;��i>�:��͌� QqU��[f"��*t=�rf���xO�S��b~�F�@��p�3_�?@� G����X�R��fV�b��7�~+�Y5߽R��#�M�@�}6r�-*�N抯Ք)6z1ј,�72_��bUu���e)#oI�\���M��a��o��o��K�I貦;��ۓ�����7�C�4��Rm|a���UV�޼̛�౧���.��d��8=�}m?`�-��t,Gg������W����l�����8�_C��r����qg@���#�1�m?��h(���h�;�����q�)ҷ�zkR���YA�֪
�_̤a�y�v	��Q8� ����u�8>,�6��X��꼶�s]9MoV��=��pm�Gԑ{�b��Y�ͼ�]�+Q�t�c@\�x�,��9�6�)��]c@�o�F]��A�  $ފ��ri�V	E��v���S�w8a��b*6D������/�+z���-p&�]��8�p�*a�B��K+��L�E�䐓��v�j`�UQ�y�0�ϩ�����YlL�@gT"�Zp�!��p��3MXe{�j5�!ܝ�ա�Սі#�񉚉X�>@���>y�"����UH!��ew5�8d�ZqA�3���_��Vc}��YI6��vj$)ߜ#��K^�[u�)p|�&�Mh�� ���#?&6�wdP� X	BP���O���8ݡ4	a�����ɏ�v�R,������,W!�� UFH^m�UvV2�\�M�7��5��6BR�/q9i0���_�C+����������8��O��T;��vخD�]�q���m<5{�Fm�烅J��bࡾ��~8=^�R^�q��X>�6�YUW���Qy���??=��|���3�=��P�@ ���~�L����o/^?�ᚒ��ŕ��;����q-
&+׬�G8���5+��p�C1�K���?�N��>��E!��aQ��G�4s*-N��~*N�c'y�O
z)�b�g8|�����'T��#I�V7�=F�@�buWC�eK�, �EB��o�P�����A#C�h$��ί*d��0��)���z�wlDo�
KW�{�٘�uS� �����`B0��{a��̶BkN��,�KvL%���c���N��a�K�Yi>�E��S]�#�x>L:���Β�g�re�8����c���O��zAJz�O Jl���b�Ϣ��4NG��*h#�ޏ�h�$8�eg��B�¦o�F�
�"y����������b����ApD[������j���ٳ6��<�^qEڪOW[J�C�i�d�.9E��'+�R��;��_��-�=�D��q[x��s�0P�*�,YÕB9g!��o
��:�[Z (S=�@�fIp��vT�`v�놵��)=88-��O�I�#�ͭ�'�JF� ۪C_�&R�vN�As{�A�NB�ø��r���ſ�)���l@u*������ffS��|#{"`��9���N).�k
��$���i?\��!I�Кl
^&8�F<�Nd�yF�B���f�{�`����arxn�5N��G���zs#t�[^[k��D�;X$��z,(VZ�|�)*�0v��?WU/�6&D���AI�������}^INg�P�6+D��Gnbc���7^�TKK-����$n� B+�Ѻ\`9�����S�3�D�_>�E�[S���ɺWp@�����9rp;g���)DIg��<=rx,��ء͒� ���
BZ��d
���	�v��L��1�C*o�]�RJ^L��uG��#!䠗�Z�oh��͒�)C%i��Q
r�iHHȻB�[�,�q0��9A�5n�E�2���R1ڊ�����cRb�S��C8��WdN���XP�ٿr����o�-�2>�?l�#�&���>���P�����{ƨ\��6C��KV��`5<�bÅ?�{oX�]i+e;���/*T�uџ����~�25����+v%�s�D�j�/l��7!G$�K)n�j���1"�a(�N�W߳d�+H�v�o��G�"y����D)�N�!�['����k�r���}{E�~�j���5�K?T���h��{��o|	]-Ț&M���8����(����zbk���+�TcOa1gIPe>P.��e����P�J�y��2uaB#�g�y�>�	�?+��H�9�X���'�	�sRk$4�����q[s�녜�:��0�Y�7w��J"�YOミ�j;�R��|=��|��(rv/Z�M�B1��_�1�cۛ�~Ϗ��	}�p:�(,����Rw@��?Y��<m�+I���`��D�I��<���hc���P_�)L�6�Vq����B��<���^�j����������S~���H�!�-P�+؄{�9�Ŭ�Q7��-����8 �ЦcsL0�����5���\57��U`V&��O�Z���M�bZN�V� V��T"�Q*��S��-�����`�@,�_�B�b b��ܢ����ņ  �	�fp�ě��8���Sh/��Q�������(���~<"R=$I]!pa�
�ƾ7V����������#�K�?�$��� 'θ�Ne����	�����rȺ�I�\v�scO�F���xb�E �s�R�Õ�0M�VEkT�N�W\�_��܁{�C�ܦ��D��5]P��DҍJ�tn"�̞�ŕ��l%����n���i���7�}�]����&�?:�esX7-qk�Ț0M�f�6�oWJS���A�ބsq�K?�F|mM��Ϥ]�3u�x��SK����{>:�2�q� W{�>sܓ�Ȥm>WAw�R���ٝ�+��E���"?�:�Hzdj��+]���$P�_*�p���I�4�X=<UdKڻ٦�;���ҳll�P�Bo]�
���iP8�0�8�S˜�;ƒ ��쾩������4��k=�A�
�V��ԭ��cŀ��]r9�W��sW�E��V�;��C	�ae�apP�X��-*�xr��v'��_�c=�&'%߲Sbml}v7�;���f�}c
��\j�o�7�.)�����o�A<'���4��w�l��1��0�Uak�y�FkԤ��L�
��K�m�L���Eeyz�j��@|0��1dr�&;ֻ�`����gk΍&�$�9���)k��cc8���ƅ<����hj%�~��L���ex�F	m�':��2�<,e��'/�!��G�U,ޥ�,�kW ��`�iLR�v�\4C��P�c�Vg��W�,���Nx��i},yI�a$���Xj���aG��s��6On#���n�q�J �e�RL��7A�˕��Ze��s7��f5�aR��4Ữ�V/c�7���`m�]	6�ֽI*&��-N��5��ɇG@��qɟ;���H�y��q�>d:
pl�,.A��Vm�XAww������FE��E6Ү��N��ԛ��p�t�6'_DyV
Fa	=�K���u��z�.��(yNi��������_"T�PB����:�;"QMF`��S6��'Rw<(�$��<�5���4v1z����0��Q�ww��s����Q�����A�Q��v�gb1.�Ɯ��K�"��״8H\��A?�W�b�O�e �G�U/����_ư�gV�5c�ж��1L��dV6���tvy�!�{�n�с�Z��}P��'��!ȝQ�¨'�#�+��x@���<�fT�>�4����H�DԖԫ�����A�r���H�)��@�naD� ��H
Aߌ��%�Z-�`���  +���8-8�73��8_m��ޟ^��c�ʋ��?ڼOPn���H�c�6o7��?� v�Ø���Yf�.n>%��ߘm�3��������!Q<��H]vo�؅ a�{G8Wj��]T|٭�9�oi/|YB�.��?��y{��ۍ����F���8 �V�5DCz�b|���Ʌ��+�o���i,p�� c��� 7���T ����7�w�`�O�-xWn=<�2�u�6F=@	��k<|����ÿ��d���k�(� ''�K=�
�������筪<+��ݐ=4���'w3�����4Ch�J6�<`���;B�Iy�_��eI܃�"G�j�퟉F���/7��PF���5ng*�(�l��8�C��O�Tn���ގ�I���#�>�2O&����ڡiO����z���[��t���O��@UƜ�K��O�r3�<'�*�g'�M�)�jѶ��-�|�r���!.���Զ2�|\WF�m~���#�^�CBL�c3&�cL�,y��{�e�����q�X��=2*9"�$�X�ǭ�o-�P�X���w�6���ݪ�p��]�t�%������rM2����J�<u�3R�ׅq�ڃ%�5�rI�!��}	�܎c�\A$v��S���m�5�k8��z�1t�tgF/ӧ��G�(��8�*^&0�+��,�O8� ?��!Y2_6��*�G�������!Ey��s0�����o���Dt�b�8h��AE\�Z\B��@n��|�BH]�u�"B+HkY��g�R�}��z��Laj��ix������(��jC8�c,�^6R��r�C�������U��ư:�٦��̡'U.�i���iǕ��:XG�y����]�cC])l���=��+%v��
(2��ģ6���kY�5�&��9e��оs����|[����T�@�f�@�-��Y��b������l�� ޙk�)��Nf#��$�����8!]<E�%b2;�m�<l9࿫'�Kq,M�!W��	�(rZ��!(*����N�80�!�[�J�:��c��A�v
Q����^_���݇�Fc�n����� M;N�l��}#^
��"�dI����,Vto���F�����,�:�z��Nˢ���n��C��GD�EɃb�P$c��JLh����=,$��|ߜ_�Y�F�f1�]��J�8H6�5:��F,~Ё��#�H���3�->?�s�9g��s-
�^��cUo򱃩����z3��u�¼/��6�~���$�㣳E P�| 5�%�\/�Ԃ�,��29�ɴ�����0o$Y���a��b�Ԥ����0�:��` ̚��-�\����MW��Q(u*�����k�Ǟ��-����u�@�4q:U���M�.< �o�tr[%v򭯙��T$"�Sk̿�Ix�l�B�9���vq �1�͞��9S![��(�1e��	o͚��loK�,�{��y��Gs㞺L�W���e�S�?�����d�xoXO@
9��(������șT=��Yk�$GT����5ڢ�-�̙��8�O�hB��PW��z�[)���-��:��{�@S,`1�V�ȝ[�<N�_���^۳zH��cI�A�(��j�}�h�L����t;/#��M��N�����(s��M�^L�y	u sY��o�q#��ܞؑj��qK<0�Ὢ�"��j��}!�V@�_�"���S�(7�m�,�z�g 㸓B��Ȍw=bJ�n)�Ē�<�N�>-�������]΋����L��������W'��'%S�j��������O=�@�u��8���k�/sh h�+<�h#B�eZ^���렙�}����� �d�y,UL􍷣�����u�A��7�r���y��ʭ���T6�g��N�C�SUFRGC-��/ܛ��bN.��f�D�pG���x�|j�v�6��zx�B~��0��oSm��m�v�W�-6���C����{��O�p���A��Ț�g�
C����"���ۡϥ�.�p�ZX�iPYI�y��s���Q%؂�6�@PKX�0;��YP���u�"�\���f�&e�;Ѳ:ũ�3Btv4͟�z$�"/'*����Εa�~�����~-O̓����vKߪ� ��U�O122}$���^R�s=G�:E<3�An��3��H��Yk��1��~�-J�I)@���iE2wJ�����d�H���L\�۹"��e�?"C�B�%�Gc
0���y�/�Ye$��IJv���٠7�������	�D�����ln���N��ւ�C�.!�ѯYKH �~f�>0�v��x�@)����''e�9���7٧s��Y�{�Ne݂��g�.ޑ�偱��*��}>}A��5s�h��k�mo�ԏj$ۘ�*�,�ϒ5�>�l[4b��Y�M�:eLY�qw�z��f�9Ǐk�+j���<ZDk�M�)��ȶ�6Ti���#]��5BI����jz.3���W׺��3�=Ժ����!�?�nɵEO� ��2��0�-D�o'3��@F�$֑o����o0Be��z"�����]���Xp3�t����$�Aߒ�R8DȆ��"Ɂ"�\�Y���Y<��b�nn�M���ܪ?��P��=v"�ez��x/zq������@���
�'�5+��h�F��������I/��u��O�4��F��%�&��B<�љt��/>'�jȘ��Fd͸���W�U���s�����Y/�m>im~i�q�F��k������~�ia�>���<��[�s.�\V)��D5��t�߳���CI*�`���pt��YFT����4��C��8ǟ��XM����ah�;�8v���&�E�7�T)���������c�ȭ���D�Bp��5�1�!`�ӑ.s�d˛�P�do��s�$�&��%[��P��Һ�qw���v�`�C��2�	e�����!�{g߽a�#�UmW�W��RN ��l���=w�]	P&7��B�=�}Hdl
�Ǭ6�5�M@�ڼh��jhr�@�|`���"�ΏR��6o݌�J�t�u�;�(��~�"(��/(x>� ���{��ju�i���g?@ʉfѤl�Α�� �x;��!�D_���zו�򛕯-�v�4�m�Eݻ��Y=��R�U� ����w���t��6��P����4hޓ�EϾ!�V��gg�|M9GD%G*� F�.�^\����w9�F��S_�g`H��9k��+|���M^��ޏUye���h��şNt
����ab�ж�6.�8�{��U�z!*°w������`sW=�ȃ�ʣ#<DMz]���H�����/~��1;f�zU)�a�N�K!k��e����˓����~RF�Rϙ���=��s���#K��3��N4��jJN~'��q���p��h��Nq�������&��*�y�[�6r�ᩜFM��@bV��Q�o�x2���G��?虄�pz�z�1 mK�������,b�L���ͭ��7��ke/G
��/���I-��Ye��or<��VGm��\s�I�+����puk�ԇ|�� V{1P�2�s�G��aÂ���8:�,��w��3���n��̱D��ZX�Mx���v��)�F!�=�����
"�m_�V��[���\а�$�Q�w2����!�U�{��'b�R��!���(�2:nێ6���R7s;^�=���Y�-Y_+��T��^���+x��ߺ1�>"�:�&�sP�md��R��͵*f:�'<aY��.|� %=�Yj#��������RM�A��6aY&	�aH�V�[��vr�Ӯ-8�H���{�4�l��V�RWy�.$��nJ�v�<V%���X�3Uiխ��,��2��P��
 �YΪ_��<Y��E-�I��%�m�y��~��b%��k8�U��ַ[���.5T��'��aO��6�����G"�C�t���춈�� Cr��K����'K@��c�c�`$Xsɧgz�ψ�mP��m����i���$�q��~D���a�"b�ط�I�r���:p�g�IHK�P��X�-���(�?7���m[��G2��H�u��\v��_|��k������ʞM� ���¬�9��\��E$�@$-�<��aNr��8U�X_i�I�l��t޹$/#��6��[a-��{��'�$F�L�]�L4����� ���{��;�H�,��ƖE�'� v7�m�fpe�>��$N/ϊ�]�Sp���L���J�4|kɞ��3�uD�R��s�>$��ω��O�g,������zN�PΥb1�;
���ڗ��l�T���ڽH��F��	�N���U�LK^Ⲷv�����&��Ri��a7���
����|Y���2g��mk��A��z,��|N�z�_#B9�q���6�6u��q��'�����!�����T�!�Q�r�,ވFc>��,��_�`eL����2�w����c+)W��Gh�g��LAmk��3�e]���ͱ\ĺR=W�H��X�6��4�[i<����J�� ((r[`�G7�Q�)6����q����x��F���ɳ��S����V1�8$���ã� ?���bp/{����ۨlWSo�j�J�'��������T���>�
S�i-�hTk*k�v}k��m�ɗ҆z�U>�c� �E�h��s.��.Ċ�5�.ʚ�N<��`E�N�'�A9���� :��<�&ޓ�Rn?">	�/�������M蘑��E�MVc���默���r	r���J�!�N�Ӓ���v�t��.���Y)ǜA����h!�z�n^ܔ�3K�g��߹c֜3'F�qW�;�y�i3�uD�^���o%�%����O�'A8Fޤ�b>O��B�o� �������<�๋%����D�����j�ЪS�m�|�TXk�e�á{�׷�kv�5pTT-&�<F/��[����_�Hê��]R�)��������S���ޠ3a�����_���m]�(V�����s/�(qIm}�_�>a�K�#��7C��Hgg�R���nJ���	���_���l&�($�]��>G)E3����[{�w!��6F5���qe��ӷ���ps��l>�u3"5����6��slG��:���L�w�
�S�Ox��=��!�i�ɵ1�*Tt���ڋ�<��Ma�0�b����\�m8�d��6S�w�ey�ykp�N]�b1
�nϔ\i/�r���;q.��|� 	q���?D��:z,S�
�ƒr?�G����:��M[��r��?��后 4�*2e}rtY��Q5�
w�jWQs�Y����A�^Z���K���+��@�R� �J�K;w���
I�<��\�B�J;�F>�C;u� �=)���C��d���)�,٣�����9���"J3��"���OQG�
Q���z�Ċ�j<V,�v�
�4���{00��1��9�\��μu<�I�ӃPjϖ��jӕ+y�bW��L9;Њ�ä'4�4>>��]��o9�iGzx�=E%����d�}ſ�
>�0�� �o�����G�ц�+XP�ǽ�~��1j��~�,4�f�)�0-K��:�?Z�A��T�w<��/_����`jyR��B׹�!������8�F�C!���L�ډ��@%����݈ P�����J�ϙ�ެ��a�_Iz悖0r�9,>�Y�8,�(���ͧL���c��ND�̈�g�"���z�,עo�U=�,n�hb�Up����M�Z�w�**t��a
�Z(����|��W��59�Paa��xA�-W�Cٗ���!��!��5�r�Ś#��1�VMZà�V�� �Zޖ��JC�­�����AZ�Eu�
��� �S�/*��� Tڀ�Z09r�����%@�Z
�݈���+՛>�Ƅ9W��qW��꧃t��"mճTh�Vج�_��.�ѕ�I����4����"h��K�u�Gb�so*��-o�F����跨�^
o�j�w���4.�.�`b�JQ�[���2 ��Hrۙ�m�h��$� ʔ�H�����}����T�]�B�a2��7qpkRd6�`e�j�޲��ф _�`�+�	b���`kY7��^DBlX��<7 �Hw3%�usm�7��)F_+i��\�G�ï5,31��Q�3���aޏ����:�
pa.5?s���E�b�V�|�@�`����w���K�"Z�c���������v\nAƧA���M��U��~c���"�*���y�es�K9��'�LL�e{wSpU��xr�I �P�W������b=:��JL�F����
b�=��Jt&���Jn���R���A@�>=D.G���C��UA딂���u�̱z��f)��:��Q����I�Ѻ���!CX�V���$P����í:�)N�f��&M��V�vQ�/b~!�v���	*�vY���f9��B�Ǣ�ƵOvA�/��2I/�[�W�>Vh�H�b��&Lש8+�~���=��3��IJ(pٰ����~��a���AԎbO�E&�Y�~�ؑ�~����;ÿ�,]d��3��II�H=ZNX�f��]U���J��:�?Z��Ћ���V�Um�?�'��FV~RXNKй�<�ش%	.��<@"���鿔��!�@gI[�n?�A1����M!��f�]��F�6I+�dry`!�G �9�F��^"���H�� x��1� ���F8�^����!� #-��|V����$4�����~��b�mO��]��_K��f���K�}1��v���M�PT�a�J�4�����Roў������T�Ԧ}÷@y=�cd�a�>�x�6���eYe�7��wu~���&��P�gw���!1)�Y#:��da)��9��b�f���;���H�[�͑�L(:������ 
艖�>����MmU��-���3 }��Q���E�@22
��T�ժ s8!�����뢃��Y���~���6��^����k�<Be��(۟��l[g).*c������F�_�)��"m{7HB�e�.t$���6�J�V����Lz7�Ax������\:EjA�P���H�%W�I�mo������F�)��Ď��ӪNe��������@�~
�E��7 F�!5\L��N��r�c�O��� #:�'�n K}7{�Bh[כ�!�[b�Sw��Hi. ��%;�2�t��`M3`��}L��=�~��]�B/-z���e�k��[�nϽv�NeI��ZF�o�B��c�Vd�#mm�/TK�}��Z���Q|�k�����F4aZ'iФ*_R�@��H3�t�N�l���D�?������n�l+���=1������cE)�7��?K��k/\z����,��uaFM'7�M}��/��j�Q�b��2�'�1�eo��rn�J���'�B��S��\�B����5_�`�Z���ݲ��<i�<��K�C~8�GI�D�A���]ǭl̩"]+ǃ�u(�?�{m�2z)�Pm��C��i?_0<�gz�v}J���`9������3@%%�"?������?�,�P� J�m����K��0�8��'���MV�+�-�.�P'�I�f�ƟҲ՚��?�k�V)����-q!�]��!���X����F�`���:oj���u�\����6)4/ja�dI����y,k�hCjw��"s�N�����dQǌ��mr`"�1'��\��T�p�����o!o�C�;J�����m�.�^����x{���u����^��s��p!�^ LNlGC�_�0$����ǆ��.�]���R`���`���*��Z�_Pf��*̝9O���V
�i.����{c೤�!SE4�'L��|��di��V���B����M�	��T�ĵ�_�;�紃�A���m��-��$_F!�|ˊO@�?��,o���j�y6��Š����$X�a��|)������/z�?���Zr���w�A���=X��4�fuD��:�/=N����Mr�Sk�V��xQ�4x[�-am�AoQ�	�����aݑE}X�����\R�5�����ܱ�G2�g'1���q�f�g��5����=��<u+���Yh��WB���*'H�1�Y���(���8?��7ex��,�cz$\�� ����DuE¯
F���z�o�i�wZ�x�/>@���,e�au73������ny��><�[��,��K��]�3k��T�8��^��'��4T�t��U*�	(|��Ӆ0g�$;�]2�����P8z)Ց�'��~�<�9ϧi���&]��(������ �H�_$G휏H�$/ʥVl�gm�%�����t9.�e�5��1�V/�"P�ՙ=�᮲ <������bm\T���\6����v[���q�8�QEk�B��% hU�\q�J�o���497%Y\�N���@�*6|f�:h�4-R��>)��������yS�" ��
�
z/�$��p(����/�2���5�����J^���sZ�S.����w�3�٧"�Pv[���f�P����
��;�=�1��������6O�x�i�-Gr�����Uτ;os6�Hch�/Q�m>Y��ϩw�a6����8�\n_E8�����C< n� 8i�e��!ECΥ���f{�KD6��=18�u�C��l"�tr��Z`|��B��s*S����3����Q��ZVʕC��m��&�I����ҹ�J�y�� �F�.��c����n����-X��-�.Od�����(��Vy�6�!�}��\o���6�o$&t���ߍª` �T�d���F4Kd0Y��"�?< �W��'C�ϝ���m�b�}^S_���:0�t�}L���G@�S ��h�Ӎ�pv�oc�ά�ڟ]�����@���Ɔ,lqi��g�O���zv���;����[�O��zZ���O:2.�eo1S�3x1S�'��@"�C��K1��? �`/{�Ŏ����Ug�7Vw4 !K�{��a�aQC���]GS�*�zq%4�U0Ӱ��UX���4��×�V�$QJK q�4�� ���0h�[�i� _�\�Rt��8V�5m�rv�U1x�b������b
���p̖�B��B\S��P���:�*�UIB�pv&�Qb��\�s�jѱ�R�m�JP��:I��h��{K�� �"]�����b����"
0�P��-�$�� �Q�§S�!ن!�Z�4�yj�6�����ݝ��}r0\(�~>R����Js�?��v�ɮ9�e�)�{�+Oz�7�%���N�mW^q�i���:�����e����^���T�% ׃�OY�	"��O�
���D�c�]K��VL��G�Ѽ6��+b��-�wk���l�u;&�W�1:�:��Y�}cz4XQ�B��Y7���M Q�|7�7��\�b�'S(k�f��`�����M��ɑ&�q��1\J=��5�_�'=��<��r����S�&~�OƆ��Ȏ��&��0�t|	ti�$��h(�t��^��\�ٸ r�|Cr�� ���P�__^����H��B��Q���j4���g��2��Y��	|S�����F�w�Yv��QTJE���g��V���b�X��R��0�G�$��V���,V) C�Fn�=�r�l�N�3�f��y@z�M��%mB������m���~+t�YN|�FY\Yg1?PM���Q�mц
�G��]�x&�n���I��t�/[#!������'>q�Hm,�E�ik �T�
�R��ҽ�k��>>��xR3q�A.b�#���!q`(e��qܥ�Q���D��D����Xe2`��~Oj���pg�Q��C���S�`�Q���e���_�=�]^yN�'I�*I�С^������&]]�45p��ޢ6�dSI ��R���Y�u�eF'�GБ���<�ﰢ�2ɛGdC�З�X4!`h�� t#���w�@�/4_����&�����٠|^��2�T��_���w���qD#!�������I��s��w�V�C��Ӛ��|�����G���\H^�����gZ-�$J;���UI� bW�E�C�;��(�x����K�
Ͽ8�߰�{N�\�	E#����Dv�b�~�	��ܫ�wW�o���g��`ܣ����S�}�Z�9��4�uv��,�\���>%��m�g�yh�Z͛�����YFJ�$`o����:�akT��^��i��щ�����O�r����n��e��=#�{���|��ʬ�$��'���&�#�� Z�w����"�4,i�*Q���{�h�F�e	�,�H?����5f�F*��P�ɐ6���AN_���sur�h``�֓p���G��J(@�6j���?J��(M���Գ\s��5IQ����)�|�N�O[27��{��h�|=�3���ÿ���-0�Z����=��J@+����u���@Q2����A����T�N:�Q�������i�h�#Ѓ��F�g*ݦ��!@i�螫��K�������R�ۯ����✧u�5����Z����A�-:W�߬��e��Ňl��⓰����$�o���[�_��9�ys��ri�%`�׭�܎�R�ӑ��s�g�|X�_���k�f�FeE�s�R���N��0����,W�L�!���4�l��r	 {E����$b�1;s��_�U� ���&"S#�מq��k԰�����k���(���m�`6(t������F��凉I4)�z[�x�+��&.���w/0������3����(լr���=�[�ɐ��C��cEs8�s#�雰���N�1\���!Fwے��t�M"�`%q�V��՚�������ݵSo�����mʸCs`�m��/�������n���������?�%��-��$7�������T��zB@��A�|�&�^�\�Y#w2YOH����s�!�R���9|�Ua~(�r�{�הOJ�>eɠ��D��*7���)�j��M��Gg"��l�i{��m{{��|m�!�tu���1g��@W�������T�L��z�q������lv��L#��������������)|��>�<������)�6=Ƞ���6b��Z������-_�ۓ��THZ 6������wꢣ������S�f��_�Un[�y���?<V�v���=_����Pj;��r��RuR�f�L��(�?�}2��o{����ޚ"�	E���������%�.�S�SK��0����*��+~(�T@���H߰+"��*�ѷc����1V�b������I����8�I"؆�[O���,����P��k����sW+B�wb�Z;i4�����3n5���'�]�m]�b��A�?#��>�ܮuPrT���c���t+F)��6��)�m���)��@��}m�]m}�y��&9n:�U({v��ΖU�R�2[�s�|RN��w����~����t��?lB��e�0VUݸ]�ӢkBa;v��u�ɗ����cE�r��"\+2��c����XCO��҆�y��)Ui�)���k�&���|ر3�ܹ�q��/	:�����A��|jl|e���Gn,���@�x����h*O5ק�>w�Sї�P:��rQ���"���Ӕ��0��7T S��֚iJ����,v��O��)r��y��Y���:��n��� �����Q���\�zO��(�;���/;	f��?�\�W�[�QKƺm�7��?5A�XI�+�v3�!c�	]fH�5U^�O�ȃ�r��Z-%>�خ o sNJb dzge�iH�}B�6͌��c`Z��o�M�+�ǫ_��q�a�7t�ޣH�Q�>%s�R�ڻ�w&����A1ք�x�^��^��dփ��U�k�6�+O��$�>ǋhF042;CC"q�F��~�g"o������0z4T�� �rהE�^�^�9<NK!ƺ��*�� IĪ+��:o-�N���sy+'-�͓KN���/�a�r���=���&>���4�g�*�I�ǔ�8�?0+,�{6��{��xmr-~>�v��-��2�HbG�"wN5ƀF���L���� �{�X������RP���KP]��O�icp��%����+jO�e�Nl�o�*����`Pg��o��f�b�hrK�,�{յI㇋m�2�X,_���:����k{"-��-��P$��F�]����+Hv5x$�?ցDb�l��%O��lIoD�;RiSG��Ty	��ک�39�ꩴ�ט71���V��k�q��g��'��Bn�4-5��@�X�K)��{bLk8�) ZS��qR��"������-����/QF�1�P�6Hv`�����x�����~�ۉ�!�~�֋�VH}�(Y ��2+xT�`��UaT�^iu��(��c��P�7%�����_ju��E�q~�w����p���c��Kk���[h}��t�"�T�9�vz���f]�Kp�ʬ��U°N�����7b[��n�"�u�T��� ����R��z���Ƨ�z�*�x�>�/?�0&&��b�*9�w�9��#�ʐe=��k��$�2!�@m��a�t+�uf����Q�p�*�w�K]��-)|����h6�w���[�3�t9NR-�qG�%Q�>4��,�ee�V���z��A��A�?n�fΨ�seQ�e�[�b���ߕ�#������z����0���������O0o�w��y	(h
\5
T��9Q\�"�^�Ķ��Z��ӽ��a� � ���Hښ�d��t�:+���.(2rJ���,�R�� �_;�����.(�mZ%��11����Yf�����~��zf"L�|�r%��y�z.��>�a����$/�3H5�����'O�^ʏ��h��ż&s�m�����*TD!��@*C|�P,v���:��ɨ�J�aQxs��2�ϮĎ{�mr�o�b%ef}{ea�~_c�cJ�����m_�@�ژ��M���D��b5�����FOj��ZRf+D6��_�J�y��m��^}�x���қHd�d�Ha���̚=$�	����W
7��A���:ϫRT|�c���$�X�k�4���w�>��l�ߩAb]����z��zq>P�V��J���e�����B��ƸF��j�)fh�g�%�+�F�e�����1�&�D����R@�0AW��F���ʇ�}!����G�p�S�����z٣q�Ӎ�e��Wpa�6-hnv2�ե�㗙Sv��:� L���לy��5=xŢ}n:�ߤ�I�㴶�Fv���e�5�����x�i,�Lq��`�\�E;a,�������8�0Z+)��G��\�U!�^�YnH˞�`�� �����1�h/Q�h�?7�����\V�h���''uLD@4}PG�R�ު����=#m�N��kZ�zI�e�9��/È�Rn�ͦ1ݑ�J�PcX���f�s�p{Q�(J���9M�r3��κ!��c!�e�"��.���>�Qn�}�F�W{��]A�O��?�4���X�U&�_5���������w�]ѣO�'�A��+�Pi�\���^�,�Ƞ�T-e��<�E�(�a�+�\Z���.��$��ܰ�cE��t�W�ōe���w�ߥG]�__�h��}�Q�Ix���P��an��/Jx���̗��r�<^��Qx�0jhM��)mTS_��φlk%�x�DB��l�����7�
	��息�E|�UZ� �� /��m��'��;���_"C�"o�%N/�Ftfe ��a��P|^��hr����A#@�&��|�l�n(��Q'���Q�z�I��=���I��r�?of'~�^��n�b;`Ask���:�[%�2� %�FY�7R���T�(E�QUs�Ѽ��r���9�h�b��j!ݣH��F.���_�ɪE��f���O��bx	ݧ5�6��b�M��_[Yf�b�鯝�(��.��4�,����&Mi'h�'X����Q2�����D6�u[7h&��r��؛�_�A_W-��0mq�0�{�ƽg�D�,����U!��l��I���W��k�v��k�Y�	P,�d�4���oǻ�V�s�Hk�1<�;�ӷ�e+�*��qa�!�ٚ4�:�ԣ��`U����`�\��6��� Wˀ��De�p�P��&��7m�Z�> O|S��4�H	!%%Q|��}�=&'7:��	�>�^���$@�-T���6g�b� @R���d�x:^��U��RW s�*�Ҭx�7qs�����,��^4����� I�{�CD��]9{c� ˮ6}��O�D�)�L8�%r���\ƿ��f)j`Y�]7pN~����N0|"��c�t��E��Oۿ�}�D��P�c��D%�ҕ����z9H4�q��� /���}&�W���
(BK_plғJ$�̛������7�/��"��saw�C����2g}G���.����\Э�tF)uo�$����Rs�������Ÿ���T��Xe��y��j+�/s}`�ZE@��yሶ<��h=�@���'KU���a,�`h��wQ�X(`�mc֕ǉH����qf���� 06����!�ŭ�r��@:9#������ɕAݲ|�1�x�Ed�Ȇώ(9!@�VR��A1s����m?d����9E>ɷ�Kg�������%��x�Gɓ���2R{�4��Ugy�2� �yf3�( N1�#��lh2�Vuý�G�� y���l�TȭI�>/m�&��#�;M�A�߇�Áb�L�7q��s�B�-#P��yA&�� N*>�h����E�_���P��w��g�{E;�:��ժ�h��X{BdS�J<Z�-��ݹ.IEjl��z�-P�m����0��/������~T�u�Jhd�(=�b���br�?�����+�e���ZC׶-R�Qg�=����b�g�YbS{�}�4�Wp�]:�M�@�8D�C��Ԍ�s��}���0qx�_B��#:J6ѝ��:��|l���W��˳ډ��t�K�n,
�o�Wd���ET�?�
ϟvf &�N����z� f��X�t�)x���`����C9�&J�Ls�<������#EPn�GE5�Y�*b��-�[�Jp�R�h�YV~Vz��~���O�����O����S�O6�S���jĻ�ϗt����0Jqgiw��VK����S�k]���z�5 ���e��J�(j��ђ��+e�X� �j��t4�fvw;}�ؽ����!u��Y�!�a��O*w�[[ŀ�G[�/��S�!B�v��V,K8-`M}Pjk+jPS7��4�u�c�*V:{Nԩ������~1�XcE%!�}�=�f ٰ�`��ɫ���fd7���X��i%�B\lv��ւ�	L��Г�4��P[�I�7�	��Wg�U��Fij{�l�QѦa���od�K�:0\x|�ю+�,l�G����(`�:��g��$rی2LK��P,�a��Ĭ��k�[ٳ$hh	���3�l m2������z�JD(��v��)#~\�˲.��g?���P�
�eF�6����$ ���yii�l��Q?���*ra��9��` �A�}!d�FY��|��`݃\���r<��x�wQ�����c�h6+}v�����I��ᛐ�%��f ����7���᜕)E�\R�wm���{n��[̾�Ԑ�.a}�Ef�xy�#�d*�"�ʹKyV��qyr����B/�d��)��/�-o�y�q���)�K�?'����P/��^�Xƨg�W��4?y�{\����z�����D��z+()�l��+^�\�Ϧs�i=���1�e�nA��!p;�[]�:�XMSk�nUK2�^�f袙�ʢ�E�eޡ�Jz��ỗ�^��ۓ���]a44e9zGݮr�y��@�=�
�:<G��w�X1OyrdE���š_�8�G�>���n��Y���i���w�V&m&�����X��V��`���� �Y}ޝ�sG�F8A�-�-��a�C�x��J�\4��u��!3Q�6>�8ú�ǣ�Y��gE�OpB�3���^kJN���`�OȠy �Pm���5��属x'N����#�S����D�l=?�Ѣ�:��UY!zɋN����n�Q�L��А�\���&�#;�b;�Sw���:�j8�i��ԙ/���y��T25������ �N��F a�N����r̗	ٚX������<8�K��|�̫Z��N��s�yv�)���o�� ��s�y��aj���l�]�Q���u�����C[����с	�5꺩���Q�ht�H���k������cP�	�	>s�&�a�Cy\��1�'��E�s��*��?�4��X������0�7�F�!��耹����5c���^j��C�x�Q����u3qW�]4�[��K�����O���gNr��߸������;0�ua�7�ݧ���k7�t@�Yz�i�,|�Jxb���?T�k���%n�ϩ4S�BR��kn��6��5�cY��!wt���d2(}Pi��
�Io�vb�JU��W�#	��2�u����&��B�xpP8���8�����bns�\��p�W1�Gݩ�d�n8�=2'h��{�x+�=3|��V؂������z��y�K�]m�����v�P��a�,}�֓p��ѽb��{Sr�k#a��-�Coi���(�>a��r��
����p�xrm��\�9NԷ>ԓ"����4�U��!eZ�zW�h���@
�i7f�nz��L�`�8`�=�ӵ���r_�%��5�Y�� g��u��=�y ���4�T�Ŝa�p��Y�_U.��4��ϘN��p��P�=�93�y3c��)�j')��w�vz�3��WLdiZ'���y�$l�I�	��Mք
���?�o,�2	���`��m�HB���Hw���]��������^�6�)g�u�5E�[��x7��9��0]�4"�5\IY���l�8�_��l�񒘄�UkK��;~��$��!C�ߊ$�x��ErM`r��=���ed�h���c���|�����#xa��D$s�.�st�������h�Bb+���Bl'}��2������U�#���dN_a����|��~U��
�^�>4�@��ҭøU�ظBZ�ر���Q��jF��F�&*D-{5T7˂{�����]u� t}M�J��3���p���gR���o�|PDw��[C��E��"����;�o�w	�(�^A�XV��dYs�Sa����}�^K��#B)�wO;�|�v����1\�I�6����7�K��|��5�Ƅ,��8�B,��/�3��󩲪I��:��${p?z���8�,Yp�Õ�* Ϗ��@"�i��3��eN��76X5f�7k�� ��9�����oHa�N�X���^X�Ek�F���2�qAH�\�-4!���>`���@B#���O,��	u��C��v#��"�s����jJ�X{�n�H����w���!�!��\����dӢWߔ�
�K���� a�,]����:�:n�ty%��c��G�O�s�q���W��ͻ?M����������9�I�sb(I7}?
1rb$�����SΤ�wB-h	�׏ڇa������|��99^����;7R �$�d���
�f����bܘA/Ä�?�F戇���;��#|ȸ&�`J`I���� v[�=e��f49`��*�R
��ME����f�����h7�ї'[�;_�ő!B�-6�s@�Mj�~�������:�U�.w�]����@�l̷�S�:Iį�4#Eه������&y=��߃N�1#K��q�&2�k}������+��j_�G�D��@n]�����z� O=P�/|�A�ސ�G{=+�EY�j�r>i��'��H��U�x�q5S�8q��gP��7�E��> ��H�9B�����|1�=���dM��G�ic�?`݈��[���Іs/�3���
�g#��ڝ��z8+"lJTgyE�D�ΐX��m��_�#��&���>���C �`P��n����%ߨOjw���9�0���|n�r����@c�lV���9�!S!����O�daE�F�4q��xN���P�����MW���.Ւ��k��&�o\b4�7 ��1�|�:K�-�iO3S�iG������M�i���(6��~����B��Z�מ��22�PL���F��p��P�|�e׫R4��C�in��L�ɺ1�f�Qh!�D�S��·��,�U�n|WV~@�h.�i�R�)Q�@E�P��;�i1š�T�9���&���+O����rj���H+��$�+3�%f��H]��l?r2��.��?�W'A���
s���s�,�P�]C؍z��qҘ����Yχ�q�n��@>���8G��k;2x�����uL��S�9�b�7U�;�#�\��V-?K��Nf��֣�>����vbK���\���O(G�`���A�ZY��g2xa@�%Ʌ��f������ѩ�2��g�Y"Y"#�?��Uvx�i��L��eR�xB�I8��nun�S��Cl��E�o�EO����X��a;k �Ëz�*���]ms�Ҫ(c�pF�
��h�cPy� �zO��$�iC��O�R�W���|"����ܪ2Ţ��1*}��Ƨ���͂�St��zH��^Fޠx��a"����:�A&\�L��gF��mq��%x��.(��+ng���rJ��F�]X�
-���>$��q���l<Z�ڷ�nFh���gX#�?��!�տ�9Ǉ��~��I�4 ��g?j�a/�N.Ζ}�{r���-,;��)����Y��'ϔ&���0�$�����	���ò�X��Z*Ƿ�K��m����_i��r%	ח���Q���n�>ڡΟ��PE"�YK��-���5�Y��
��ǒ���<Sl!V�2��!�h숱�����e�>RO�h���c�@�t�7iV�"��v��%�A���Η%�}t7��5Z���_����֜���x\,��\k�}+�FI��zu�Ow "=0֏��-��9���iQ{��GU��4��c�fo�ܤ�s�L#uK�.d�ș�2����?�$����/�B���f�N��>x���ަ�0<X��9*�6-��w	JN7l�֜��cDU��Փ��u�6� �l����p�����]��-W�*�E���j�F���`�<�#��ġϷ�XN�����]0���l�\�^�)>J��O��������0���2"^��sS�:y�&<{�4ķ�Ro��q"!��q�- $���lW�yu��w=#&/�`'a�E�Rں�z++�'�J��1�_'����`mZ��x���-���G�6����Sތ�,@�v�Gw-��фDn�/�M�� u�iy�h�����:��:׌�I�+=�F��3��2̡��Hy5�9��(�$�'�����t�KD�2*�b��o蹈�0�n�[�����W�
#���V����В���{8ۈd�LX)�@2�)��Hn;��3!�#��_�5Dv�Q��5��w�}�	�V�6�u�eFZ��* E{X��	D��h�v���R־t��VW=��@����h�� �����Q��u��̡�B@���G���L0�/��Y(��i5Fxz�'昗�-"~c��v���!"����.�ߺ�kS�/$>�27rU��#��*N��D�$4��DQ"�;ad�Hd�����3$	����W�F��bow��y�P�7���R��>C3�.�dz�R�3>�gy��u�f�Q�����gW�ō�Ѿ��y*V���keua��rd���z��+D�7��*Q���Ҷ��;G�l{�دU�4e����ea
IX4T�F�%�]����7�_�%�Cǜ&HB��b|��W�/�V������Z�FC�d�g��Xw��J�k���LuF ��Y�_7��T"�._VF#��_h�+�� ��T�[�\��J�x�;�#� ����f48N���ɴ�q�u,�N��J{எ����LY�>ydA U�D4d�'�P��	�t�C ~֗�!�l�-����ņ�{z/��d�%�W�<%�ځ����٩\F��N�
������ ��������Z$+7��Kbx�7�Je(�D?wۃ,m!��L\�J�j�jvi�ћ#�@�>1r��)|[
L�N|^�aM��t��؆��临�U��8�[F�I0�ô�-T;X#�D�h
�������t��Sp��+_/�������܅sN'�~���)C2.�*Ӭ���P.��6��Q�r(��P��u�J��0���I��F8�z���!�р�}��4�j��D�f��I��Y���肘�:c����V/)�X�d]�k�PM'��T�J�0�H����Q8`O�ǋ�]f���Yv����R�>>�U8�:p`�F�l��&Ҷ��tN��.��C��L�� L�@��v�O%
�?0�>q����wNO�f,�F8S0�!���뇐��/�Qg�y~��4��|'^fj��ӨF����9��ײO袍a��e��K�,���+C5�$Ϣ��T�Ѹ��#���(f@O�D��b�WB�+۔�ǅ��r��9Ot������'wl���~ڟ&�Ed���5lK �EQ����mXG�DH�`��i��D>ce�S��!��r�����I���w��o]�4��Y������2DE�dC>S6[���K�-(hS޹��m�h��Bc��Nh���A���[m���r���!$g�BCh�����"��i
7��W.B@�I�������,��nO<��.㑪Ucw��
0jđ�L�R�[�����c/�R�$qLr���}N�Sّ��u��!�Xy#p���ի�����)�(�K�˶��S8�s�U�pރG��(=�&xaP$A/�+u�y�����Ě��(��r+����B�x?1l ����ee�ӹ{@$�0�JQN�I)Uo���|�/,Ϩ
I�w��\?�P�0n<^����U�҄{3R����Z�9�0VS�W�M�Z�٭Aa�P���"D�ɪ�i<�����$�7�p̔ ���%4=���e(�|-R��1z���B��R�HF,���������(K>e�f�O��Z���l�t"B.*m�{�R�T��y��rÚl�-B�=CګS����2��w\gEAa~���*DȌUS�k���ܦ����m�3<2�ǈ+S��VC;�  ϒ6;�_���a O���h�����t��x�v;��M{�f�%h�ے$����%�l��)nc�~��ҷ����h�;w�'��Z3�¨�ز�^T�}�T�P���΀�/�tJ8<��u�h;���KX�p��.kQ����}�݆�s�i�����]�"�Jm,9�.�����r�hH�b���D���!\l�a����"ĥ�
U�?�}]r|�*��2�eYNi�!s�H��O��(5=�ȼ1�/&����`Q$9̶ ��,H|d���EА��_a�iY�;p��iA��LTO��M.��1��j皖 7RC��t���*�k���x��p����eC�S��(h��g���k�3�gh��� 5G���Wm��N^o!�3^A�,iW����.�ʶ&)2鴆B@���ˇ �Ԝj�M���M?���	��2�k.�s�g�>��q�c)41��_0��g�[����hrM�o`�'*"u�8!��(~v���J�PQ�Þr�iw=���<��9�d;�����P��QN�����4�eԕ�K	��|Sw�"��hEÉO�x�$񵙼�����GL,p�$�	> ;�m��r�U��̀��O���b�W�QM �vV,ˏ�N�)ġ�MW2X��,���asN}L�!��V�|��Ms�d��E Ww��ٖDp鱚z�q#@Lt��D��X�me�GyC�b���e��4aG��՛�Vx�7��>ƾ��ru�.�#�]]�[�;��,�����ܦ80?V:��i]���.��c����������P�S����3���Aa����9��2���ʍF�DZ�ve/�@8l�~� ����'��N��'�ݲQ���.Ϲ�EZ��i��=x�-�+,G�*�*Z�L�BNAS���W-���g}_�5ؓ��컩�y]Н%�K?E>�e�P���|��ƶf	N,����E!�@�:���ceW)l��R�ſ�cw�,�^��8��:܂Z���&ȓ�YIì6������[�w[�ލ���>��)�6~�/LR� Al,��H����Z�6�� ����*��!ݨ���&��S��^���	��p����cb����m!��z��Y���:� q!7���%����J�).OT@���a�b�m�f��P+�P�u�?BQ�IɁRz �l|AVH{�K^#Dk�(�wt©"V���G�wk s�3yG���ܴ!�!\ϭ ���6�'�!�^�X>;_/��o�Vu��h���L��˰F@nk�2�|��=�P���@Ƣ���>��'+roYz�	4��`>��R$�����w� h.|ars��/��"ҡ}3��GC�Y�r 
�P��5��4v�=�e�M d���R�6��#_�Cc,�3�\F�Ы.��Da|���*�-�5=l�]%ͤL�uN���*ʑ����8�~i�N0��Px"�>��;o��l:2�y�t�"�}�h�S�|��������́-����c#�":��6�'V`�,#��P��vP�ӏ����#ZVa�<���\����z�������$�E)榴��J���Y�W���6������=���n:��k�D1��DO�R>���;˅*:�[��J��1�����7+�_G��Y*��NGrJ��i�Z[6]$)�m{[�^�{���]y<oYj�/��6��_��4�P��`x��sT��T�;�w�u1:nc��<����Z���g�٬�����O�}��ӆ]����$@�[ �L�)�x`^���rꚈn����o�
Pٻ�6(�f_��>^v�/��eP�[!�=NE9ou0�=�G�����7��3����ȣV�ie) x-�^������OMm��4W������VUt��qki7�+�.4(Uu�Ì[B[��A
`-7��Ev57��8���U^Ԥ�<�m��_.������k�~cܗ�a����\��.8u�V#�UJ|���3�c��7��IC+8o߬���Av��15��2'��'�����_.���5�$#7�S2��$��.k�}�aK�Y��v���EWN�k�;��������/��q��MR6��:�͍Ҵt"a�J<[Ϗo���mu����A�o���D�z��T���(����&�:Wg��h�i���\x��|?�ES%���+�w��k+��7�������;;�4
9�Q�W�MCxl�b��?s�1m��n�1�6��,gE4���fb"E4�ѭ�nO��1k`�Ѝ��H�D��$�0���_L�����%�p�s��r�gBӍ|C��Ϲ:��Ň�vr.�vϋ��]y�p&�#%���]&q�$/��a� oW~��`�fU�<vO��ػU��tƇKmZk��Y�ML�ž9V�0vJ�6���c�I�I��x���[I:<Y��eb͙aP���B���}���<�����m^ش߀��s	�L�\|��_<�n��>7�h�A8Z��U��Q��}崎d�F���E�zFl\ܐ����~ I�QB_��'�`����4@�!�k��Da�S���lh<��]��<T�}�C���I��@ݥ��^�y��h3p������_ڬ����z۷�eO!�������!�1�I��4���C/b���-��3/��l:�Ο����H�2�G���BӰ�#v�!n��+� �L�,��Y-t�-�;�����W�q�]���0۽�-�l��w�ne��g%��T!a`FkC�{���JrD��[����OK�c�^�U�"p�ĩ���y�����#����S�	��:�gґ�wv��@���k�~W�I��'p�ف·-G���E��\��b�D��#r��R�(׷%��?�*��-i�[ޛG`1��[�^�F)[��<��Ha�h�7�W��FX�����N)߯Bbxm���}d��� �M����d`z�T��Yжͱ�)���������N?��Nf];շ&.�ipʀ2!qcE�����x�\\�T�E���w� ������O�A���B�wi&�ҡm��P_����k|�\[Ŷ�/,�#�[�64��_V��)���0���s˫�]���Kj��#���	����K�jr��k}���՛�U�8�k�w�����Q�����ȗ]�PQ�pk{�B�NIx�is�4�0b�yV� ^��@�#}kB��PM�pÅ��� I��Ϯ~3[�����s�NX2C�\�	��?B�jv��hj|�XQ�P�ݮ�3�?Ԅ.���v��"�)���n�+�_�	^��֑���`�a0���dv�|��{�[<�f,�<R��{�G\��1:L%�Rx3y�28V}
��t7�B��0�H�ޛ���pT=1j{h���c������̀n��gd�D5���<7.%�B������_7g��f$1���Xt���0�;k H�
�i
�����G+�o~ &���tT>A����\��C�P�.�ƀ��,'px�ī�quW�y��>G�?�]��J��&�E%���]�;0Y�K?��*�_���?H�Iey���7+&49`Ź�����t�	�M!�Sy�>2	�2��䲆љ�Qi��Xv9�̇Л��.y�Vt�b��OYB�2�W�èbs7F�
��f�CF���N�iP#]Bº����e�a��$ӌ�����ǂ���&/?�G��JVy�W5ˋ�~�m��͡���o���iS�ϝ&\��H���j��}	��6�t� ��/��D�U�Q)<~l���Ӄ���Жmtdu�mo�贅z�]�!&̬2pS�pe��%�Yt����%��SO7V2�V�� �cK����-|��D�sg��F�9�����e���)V��4�f���8� ��Ɯ)�6V|1%�e��9.c��U�{�~�R~�N=���r�,fQ��V�>އd��_���
�O�35�N�+�g�Ved��:3�(���_U�|�c^��C� �qF#�S����* �/����Gx�f��}�����,�����'��[ۊf�N�45ȏd���E"�?`�[���S"�o0�pT<���W�D���	��ך�P�)�X��w3�.�����7~�Gg��= XRA3�\�n�t%��,F��L�˥ӽ���~��}���L�vk�P��"��J�u8���2���{��^
��t�I%��J�g/��j�pBc�'��������^3���f�x�mz��!d���XZ p	l����?��W�R�o��s���K"y�G�끨^�<;hD�v�Z��H��@W�9� �1��$e�g%��^�~V��s��h[��Njl��T�*9��������u<2���(�ВWN���'�d8���Q��a'2GD��tbX�c�}�O�θ��]���%�|^Q'�藈D��I�j�1O>~-q�
�ج�n�[�	Α\]¼�R��t��y<�k����\�ls�sH��Z�xԣm�ڞ�I�p����^Nߠ�As�������f�j������k�}�h%�]�m���\:	& �={��^]�t�v��~�X�T��%`�ת� �B�Bz�^!�-�"�
��/�-��Lv��p'wL��z�,!O��4���Y���jAW��B�ٕ����ݻ���p������""��b�(ٱ�׹�;O7v@b��ʷ#�\�9,^�~��r7��>N�"*�<�}��s+�w$�^��5�П����Zm.��i��]�������|a��BwJK���ϠL��ߓ���|�H��ݓ�'u�mǒi(��p����#\�H6*.�ݛo=zL	 ���s~���d2��:�.�)4?�s����{5�8I�<����2~�S^s�Rw$�� :}��ö��e��u�*:�҅�J����}��ŧ��1U��^��a�[��e<N��V�*�Gt��@˺�pT�A*���n٣�dʒ��ۙt*�&��0�S³�Ϋ���Lò�wհv7�z.~-�@�-Rf������+m8��-���Yؘ>�*n���*J�l�|=������e�M��r{�3�=���/���#�-���A
��K2����:Hh�14��&^��f�[����?���{��7�`�xL�����ad7uA�R����N?r�Z��]������N�1Z1 <�Ad�$/�l0���%������yZ#C��Ae;�F|E]m��X4���1��E?+��xt���CB�3C��3���j�s��D�yG��yT�jNT�au����g���[���i��~��!p�wc�p��8Cf,'��
�i��D��8�r��O����'f+�+��V���r]U������z%�l�\د_��� e���k
k�|ά�]�X��>�������5�e����-qS%��i�$�5J�8�b����*�sYo�cc�K�Ȧ��,X�ȵ-�L�f���"�"�e��U����nu����l�P��ni�+
�v��(=�{.��>��{��s�����i/����`�+2�.7Z���L�lF-!�� �x��At� &�`���	���Q�Lkp�W�	��Ц�
�8�Iج��E�&�"C�h�ʈ�U�0w�}a�FL��3*��S:&S_�˕K3DIu8�d�1f��TJ��������GVSƁ��IgI�+[�@&*��q �q���g��j��.�k*N��P�8��Q�Z����N"V���I�x`橋#(׈��='���
����Zk�s�yf����5������wp�Z�n�.��+Ǫi<�#��w�"�SY��w�D��L�=���(˴<9���,I.F�>��A�G���t���U�����q�,�;�ֱ�IZ�F�Te�A������`�L��#�f��y:���Kbf�U�Z/sF�_J����6��L�T4��Y��h������#r2�����:���\ck�w���g�`�k�I�3y�G$b0����z�Z��C�s��L䄪�-�At�UoFc�N��m�X�{��O�[:�_$�rm3Y���9�+�ݻ�,� ��
)5ܬ6�(:������8�9���q˧G$�U�ȴ��{dnjB����=ԋ�ʢ4�Gq*��P=j�c��U��ƥjͩ5����b�2�o�R^!���{3�"�-{/>��K����*b:e��tD��/=,5lµ������5�GŹ�DP�cM�uy�t�߱%�$~#���LV����t���k�Q
�"P;��j�uZ������O�Ē��������A9�϶?��z���kq��ZF(zR��P ��U�:��I�v�x��sJq٢��e�KI� �iz;9�pt�9��^�)��3�%�Q"����Ư�Rlvp���;?FY��	U���-4�����C����Y	u )�M�?m������{��+��ѷD6E��۲p%
�S�#�Pl�F캽R�3�p����ΎrO�&��BQT(���ߧ�:�����-�c���V�G�����N���̽1!-"ݳn:�H������=��Č����I���O����5;.���,� ϗ�k�:͸\5���yP� oj;_�b͜��Fk�r9Շ<B�o<��*aK����C�w'+�";�ka :#S[J�ś�"{A5�0����cqX	�D����ɝ5*cVէN :@}����M���@U]V�mv$���3���_�������Վ�%��K\����X��)�W�XCe��sܬ��|w'�Nt�z���A����B�䍮�H0듺�kq���X��&��?r}Fz5��m��؍��cGoyϘZ�����h;4���L����Ӏ=M����z��w2��W@����/�NF��IF��	����J���.U��8�E��j��ȝl�8K�A1��[���??��~T:0��"t]28������3 z�nbFp�'#�.!��%�n c�����b������2��5YX���1�� �����oD2R�cV��0��x��Gʎ���H�Bx'�gec�c��|��q	P�iŻ^��<r����Ne,����P�Ie��#y���vH���q�����t	�6A-�r��I�Tx��C?0���u��Ҝu�a肶�'���~9����Ug��l�2�EIo.9x;ȍA�5<�&�e2b�T�xTfm��^g��pR���ݓJ�'�b�қ{�r�I0G��zku|�[�������`�
+V�����MM՝�.;�A�#��G 	86�����g�i5@���t���˶������ya��>��w�!�9�:�`���g+U�Y($�Xi�NਁYE)�`����*�B�у1�{:MzI�B���H�)�i:R�&�����wSN��,�ظ�j������d��0y'Pz%�l8-韣u�}�]�V���<�5����D���uM�;d�H�B�3������`��z O9z'�|qE�Ə4q'wQ�;���SV�2���y��5�貍�����;v�g�����L�����@|�̄���r����(�J��ǉ���g�.�@W�8&��7NR~7m
�n��9�������p�$��^f�T���_җ,?�Eȡ���*{'G��$��(����h20�>�ƺ+��4�DsQ�t�e�!�9P	��ޠ|A�D��K�f�'̞v���.2��ź�}�iI���|�V�t��.�C�=���W l��T�U�zj��i�L(0ZEf'��B�S,b�H����ǹG��g�:�+6�8ͽ`ӂ�WX���`��]ew�t�)��j�*��|���,�җ�5�01����t��@"Cڐ\Y�<5	|?ߦÆIxvoN�z�����<q�L��NE�3Ʒ�V�L@�?Cf�{�V��r�!�k���[4HW�>ky��]:��|��~��>qF�?�=�A�Я "�קD�ྮ�gȼlǙ � ���y�`i�IXJL�Ԙ},o*�P�,��.Ng�g%;�.p��M�ݰ���<�E�h]�y�+O�Q�g�K�F�eL$�9�������L�
�m�xU�'�2]����ivV���c�����m��Πfke�q�MG*�z���G\W�n�m�7c�9���"-b;�mL1(��������4��돹D�umA+��'��*���}i�=Ñ6H����PcO4�U��8�~]�b+�*���S�ۯ ��O���� v)���e=��Z�(��%��B�&�<������ղ��g�N�@rT��g�<�: U�0��^��E��V
�6���;<Z?l0+F�w� ����O��3�_cFIS�wq�;W�D��P�|<�ވy$P��)����^�pk[��]����Hټ7�bI��s~�/h����gxi����^�Lm��\]��PD0�z8r�e�꾳�	�͛��;��� �X-LJW�28e.=��N�配'0��դ����q��߈��X2��_��0� 9�� �#A��g��;�c�����IXnQ�O4�{wx�_�����Y>�Gp�ڌ�զ�HJ���اm�3S���S�U��D�kU?�������E�d�G��ٹ�zCݝ
Z\��qzG
;�X��܉`~���X1ar籫�y8K�_�kbN*�J⋛���ACuᜄ�h5 w�:�^#sW72���P6 ��=�A�h�VMX�^�sn�I3�����qa�"�Ō��K�x\V:�����̈%xsv�{?���Wn]�Ety �=�'5�(��;т=�#�M&꾗$C��Ԕ�k�*-_���'K<_ֿ(1��S��(�3�`�~����L��͡e��-��9�	BO%٢�V�|�t$�9�N#��*��G)$�MRM9Kmj,!9媮����c�?���/�֮�E`-�7�c��iTsP��:�6Zy��<�9Ŏk�*�C{���6��S�U�����a��ϳ^�P}Mf4k�>�&Ő�t"���xd���/�::е�|,�"ȩ�-�@��(h?�d�S�2aU����?Ɇ ��:Qe7�����j�'�R���_,���#�';ѫ䳷\��Z��C�{�_��|�@ޝ��l8L�A?��I��z,'�eb����M��{l�UΥ �ʩ��z/�C��Y<�?�w�5�\�z�OH�^G���$媫
���[I�>�t�
��X�9��M~�SI��7��ږiQ_�c���9r��C +�!�� �`5�1���6�̮�#��+J�'�Iז�H%֣��G��I]�����^hv��p<�%�d�PH:��mJ�QM�PkVl�?G�gE��[�J'ytA��6��v|jF�߽��i����35m:��>���g�!�B�W��hY�����ڒ[�����Oa�u,�z��օ���Z�$�6P�X����,� ���x6|G���^1��l�e��|r� E	=�Yf�nf.*y�t�%
Ű'l/J���#�����U����"p��j�%@c��q�0	^r.�1�hJ��fl����]![�m������#QC
�-8�'D����>m��)҉��~GRp&}�ܙ�ra��bd߻��i�uZoMF�9L:a/�. ��G�E�����hMF�$(�ET�n;�q�xb�ǥik)g3��7U�,�]T�D ���S�̞E-p��E��d�����e�#�c�C0�s�q�?I�6X�Sx���,���2Ɉ������g��st�v���=G�Qט�ɇ _���ccd�Y�݂��"k�t2%��&��o���x�S�������z����K'H�u�-7��cǫE���d�l.�g��6�k��=��p3z���S�W���,�l�	��#�r�=�M�v�I�rt)�n�N���D�d�ɏXM<�Y�!��G������E�gΓ$�#>��t�N��8�� ���	#ޡ��c��w��?�-�4�.ݿL�O�wo�R�@�.g ��Y'���u�>������+���PO��[6g7t���O��aSG���� ��A�x-��r3�&����oD��Bޑ9	���Ϣʦ�t�A7l���
$ֆ���V�����4�ђ.+�2��?�{/ڍ�f�U����>��se��ͱ��y4z���4�OK�p�t4%::d������VXM�0�;܎U=�L/2f���.0V�ƺ&��{��f6�`��$�(Z�hpt&�y>O�5���i��R����M5^۔�u9�_ ��!�q�� ����=�[�"EXf�1'��ڞ�e2�*���J�}-�E����k}2�`�� 5T�%Y�<��x/l/=�ʼ��OȦ���'��K'o͖��}yW(,)t�y��_8I^��xG�(�9�T�eؠb.��.��O���Xk����V")c]��!�qt�{C=����Ɩi�Dʰ���r�[N�җ���p��\�I�ʝ <�Σ����}���J=������g3K�c8`H"�A?3����Td��Ý�r�J��\В� 
��rFC���\
�e�v�Ce!~C���(I��V�`�zl��3����E�����j�
6 ��b���Դ��m���m
z���on�:+����U��eP�Eb� �"t��\��WK���k�������tɈ�����*�Qɤ�;������ۮ*|>1��7H� �%`-|�.��;>��Z벊���^r�FR��θu�{�LwGT��Ĭ�1:��ל�����} ��n����X�l6�C���X�m��pC5X�N���8[�o���A��BB�0U���5$lIN#vw7uAay;���Ƒ+�{�:�>\�	���60��{z�v\VU7���W˲W�,1�"��H��������v�ѵ�	���2��rb��/�)(�D3��|) ��hkE�\���F�|]?mA��oh��;H���6�6����^4�G��]b�h��a�����R���/iۋ:�"߭5��M�^� ,�T����qu��1�\ ��8�X�O���u�=yB�B~�~�}e�lIOX�	B,��&���<��[l����襯u�h]ݴ�r1m]R������U�]i�HA��G ���v�ImG��0��?_��ϝl.����o�Y���x�?�{l���ϑe��P���m7x�7��b+�į.��ݧ̽Ax�K�u���J{��%�c����$�{�$��\�����.�]��h�Z|�ݫSJ�b�rΑ���Iv�X}��A3����ϲF�^�9-���!s���0B����]����Le8*���O�O�G��eF�o�����)���#����S!Tmdp���O�E�%�D��U��9����2D���!e� �3��_Ơ�M!y�����8�=t{���x�v�314Xlh���'������ӷ>�I�|����+r�OnB��������w��d$��7�׎O�J5*{w����Թ�a_2��qz�\g$l������jE�%Sm�w����c���8ݲ��Iw`�V��e+�W6Y81ƀ�
A�f���I<�\N*E4�L(T��,���rP��j.3�Fյ����>� :�����t������Be��_"�'!��s���Q2���7h����(�=y�6j��vlU�ա����Bd���=�P�S�bOtCְ�"\#ۃXd�x�5���J�F[�3��W��2�V� ���mE�,*9�_s���ӖvE�\D{K/S~2ES�ҥ�7�!�O�o�҇���(�7�[PcJ*���ܖ�{<h'g[_eʣp�3O�QUt,7X�О��?��飋��팢�ku�xNGgq�/���."M���a̐=�*�.sN.d��=3l%��|&��ޑ��eh�fT�&i�#J��0�C$̃ɜS��)Օ��p3Ym˓w�����X�r�ݾ�v��4�^r<��[*
}j�3'�=�瑅c���$*��)��Q	}ùJ�3mϪj��견�@�2py���h6�a��^O;�4&H�[}hlT�n��n�=��'sk^G:�*�R����ƯP��ȫ���W�z��%�hP��>fɁ��C�>�''z!~w�4q�+�bR�Z{�t:�0P=���"�"2@�v�?�|F�^&��X4��<u.��U���L�u��w���ҝ���6��6��k������XK�C{?���8�ZaWE�����7�O%������?��҄;�:��W�R�-7A�ďH�F�B�C�%8��
��QXAO�24�}����� PÆ=�Bo��m�EٶUvrL�"&�1�t�vZ���$��֑�ytS��ͫUi�ŝ�#G��Xx�<�a^�M�T׈yR����`�u����ӧ�4sֵ�aS!1V^����N��K9�6�
�l%g�I�Fg���VjL�`���õDdt���USj_�O�<�HDK�N�D��${Mx��Z�j?1�Sd���#kn��}z��<��P,�q�@��0)16Թ��4x�0J`�p�ܭ�i��]m���Hg�e���z�ʿꢐF�z����"śv�B����H紇[�q�����+8\���Px���*Zl ?��$�4=�?CV��>ِ�E
�Mb����{9|�Zd6'��>W����4�G�:x'�R�\�9]l ��ܓ�vi� �gi��_�g�҄�C��w��;S�[eP���i���D�٤]p<�R�`���&��;�E@W.��PS>�5O�5�ɗ���DEu�du>�}w|V�më6��;�S��9MI��w�3o����{��qc@�>�T���F�y޳]u�\����&8?�j7��l��&�ҴnmW����9dh��q?�h^!8>���n���þ����^D�J>��,/�����:���&� �����C���w��lp���cNEsi&���sXbK��Z���9�A(3�挘�o>|ִ��!j���r`�
�H'o$�����2����GP�UV�Up���
�XB�Ұ���i����|(UX�9g�j�����Y�w�,״gL��� xQ/�y�����j�4d������<OD����syJHE����d���=����M���*2�íL�<gr��E�5x�@&�븂���A{�բ(&�"��#��$�Ś+�D+˯4pkpo����J<�_dx�0�|�M3��$8Q��)��nA)Gfp�9~y�`A~�`�F*1�T1�9}�~�r����|0f��x�+v'�0�m��v�ՙ��XX~��?z����w�&^�ɇ���n�+yt� �W�<��Ǵ��nSHV�H�o=�C�\>R���j�=�$�>J�[o��w|U ?�R�6�͑�7��%�~dTfE��������rYK�-N��"� ,e@9�ٖ+6�;9{<����x\�d�yD,�c$6��,�{{�����7����A��~��k��؎*m�G��q���T��/ϳ�p��N���Hr���"=���u����(`�����$ H�%g �T#��l9��F�6�)�	!���B�/e"flC�(���%2���/��Lj���WiJeUe�i��Ҡ%��N�~h�C2��5m�M��-�ա��5�42�w4�ķ<��WmpV����N��1&C��-�%��6�ņ%e���S����c�A#�=�"�gh@���Ĉp8BJ�ŋh�����"�o�?�#_�3Y<�n�   �f���:��!@;ޛ焬��g6�x����+�Hnh��?��J[�
���T��a;��,y9����u�4�?Vg��*��qVˬ�(���!��}~��������7)��>s���f�������l���y�Jn�^[-�{�4�(�+s"v�;C�$YI(֌;?�GKB���0����}�ϳ�c��C�vqx����ow*������jh�+8O^�A�����e�E�U6ʞB�����n�Xc�E"��~n��@!S�k�X����h��fz9jE\�Ζs����0�@��K�,e�L4>U��p��,�x4@� 4��(����g&.���*rh�Ȏ��_r_���+ZS�������s�K,	!N>wz����|��R���<���`�.�G�E�O|)ZM����P�N��DVk�WJq�MQ�����Vf��I��(s�<�~�<_�u��n��R=���zF^jHEJd4h�l�q�Rx��3���j��Ew�h�MeՈ-�b�Cex�T�qbK��[`*_x��@v)%���P=�Ӷ�$Y�ߘB�w�?��O��:��n&��)�0{q[l�h�tlJ-F��^���x��lV,2y�����z�@a>Lo��*� G�<n@i���S�~4�m��Ћ�}��~���	8���|B��`V��5_�/�@�}@'�k&���=Eu^�%~���5O&��p��{I8�޻L�Z=�× �U9�� �
H[�lET΄%��JdQ5u����][���b�����ʋ&b�Y�WR]%�^?�C �N]W���T�u�M$pd��m<w�˒ �F$x�d'G޼rm�ϟf��:�q��Z���_�d��ճ6�)�4� ���H]>��hEJ��hVV���bG��&o�!�1e10�8���\J(� �j�4a��K���\7��R�i����;4౗������佾�#s��W w�<ޭn��`��8�G�� ]d���C�϶e{K���}"�d�x�#}�_��E�����Wy����C[XvV2Ak5��hI��$�J��TD���,�����7�'�0����0.����d9����l�
�+-���Y�����Z�iP4�mH�Kͥ%�� W.)���]=D0u�V����!>�R�4N�4����Rq1C�A�ٳI��E�E8J��L5�'��1֐��I��	�2�1�خ��p6�5�1�$V9����y^25�3w�+߀V7����K�|�i�0|�wlj�З~@�����O#=���D�����\���}�D�9��1W�������cM#�?Iu��Z��B���(��hn�q ;�^qL��B�si�̚�O.�����UZ����=�������Ǟm� ��R!ˈ�ʙ�9v��A����\���*8�ߩS�OP�x��gKO��Qd_?N�����4w}JM%�	��X|/�|���5�hP�S���'��O0�z	�ɯ�k�,Ih��P�da>5�(#}[��a��DU��Xx����5�W��?G�$ǵd,ΖC�\��4�,����P����I[��k������b��%�C��Ӷ�G ��I�U�,��@K�6+��4�����c��=�N7�2Ë�f��n�Ŋ�a�v�q�N?�"\��x^����w�^�W5�Li���bƣp��?tf��B�y%|Tĵ�@1�ϝ ��ahm(�_�7M�t�==Q�}$�:�Յ\�)kAaHk���y�5�b�x��]�l	��vd)�e�ؠ��~apU��s����T����R� -��Zh0�h�ݻZ��S����\vBIee�q;
FN�a��5%��~������w���<Y�ӨF��&1M�"P��sK,n㱎�\�S����DiP!���2!=�[=�#�1?H��w�)+~c�b�4�r���W���pA1�,�cls�TY+r�`��l'��)}�0�ҰD%�ysI�n�_�s�Y�*y�q
�mz'-���;Z>Ԓ� <����h,ؓD0p��{�fZ ����/�m/sK�t�m0&�i����-�b�7��bS��[�d׏�)ޫ����L<�*W��4v�Y�r�:��	0+̖������{���\ @I�H~A�ğ�;��L�k�z-h����,(@9�i��s��+]�3�DR�Q5�_�}�E�-��f��D+�8����s
]}#����b�ӕ��$��}0�J=#j~��p�<�1�(} �S	��&�u<F����
���N|��ix�������"?�`d܄����]M�~��&G�A\DW�ߚvT�{�L�F�ʌ@� ;��g��*�`���I�y��u��<8��(�=�þ�#�Gx�qwis�+Y^,b�R����#�}��Y.�F/ۘ��W]S�M�.��r�� �8�-��'�c�Qk�d�#E���ۯ��@85���G]��pfY�?�{��t��+��|/ļ���j�1�� �!��`��H7M�$�=B�
eq_A��>�pc�c�"��$���:
Ҵ|�/x���G��2���eH5�_�FU�#�����\@��"�U�4�	0==1�^Y�����K����Ѿfֻ|O%�J��9u�כ���xjȁ���e��hD�b0��@wV�M��Hn�h��U�k޽O5��]�p"� �����0�k3AkX>^s�v1�m�ֻL�Ը�h{m��O��%v5W|н������Q�|�j��8�W�֧t�>��*o�� ���@���6���N���j\?���bi�&O�Vx�ƈԻr*P+N̚]N=t~5��j��ځ �R��(tl�Pk�?=	��OH�~]��C�3� n/=(�Y{�)ly�T+A��	9xX/}aX�j����Q�A��2��Yt��|Q���\�I�h�y'%�{OM�rl����u�?3h��C�ѭb��3���C%��[�t=����$��I�F��䱂�B�B�+A�ϺT@�7]ܫ_M�����s����M���_]^Kj�3������k���"�!�6�,ni�+��g1S´���mUڐU	�df���ُ��j��� (sK�U=�Gb�:{�@��QH އrx+��(���lm����/:�������i���z�������QU�w#��,G�7���i>l��V�DM��zg�)v`��{r�HL~�v��Z��GR��P��o�R,(T��\𭎑�t���'>zEGgo�� �x�sRqC��_�  ���1����QŊ�����_λ+�3C�>rf��~J��vv�GLQ�n	`{��W�ˤtu<&�Ζ�ף/�� i���(��p^T���j�JZ�<T��p�-/+\r i�$Ι�>����e�zF�gbf~m�gC�2
џg�t�MJ���QIp��Ǌ�v����Af��N8�b�kJ�eY��a8�� ��5�a��X�R<�� ���_5����v��l�L�I���ˑV�5��.	3�+")��w��/�7U�F;�H5�@����HK]��Nb.IVRm�	>��I�,�]HV$���ݧ�P*�%P�P%�(��!*��B��z�l=˟G����N�GS"����=�fP�KSC�eN��!)�"������gf9sΚ�/�%8��o{�s����)2
L;��T������)*e/Pq 2��Z�*�!#���=�ux�g�ᯏ��n��%8aWg�q��(�M�ak�G��{�+�Wh���l��~C�.�F�7��P�w�a?G�#�m��;1m��K`��+����~�s�n��.փ�F��B��J#��;)e$�D��k�g�	�L��~��!@]�C%���&-D�/5�T�k�~�~�V���q�|߅XpX7Py:�9Q�d��J��&[I�5���;E�빸,o���3��W����g�'OU��T��f��5�cŨ2�:naV��"�:���JDݮ���\����ơ�M��s�^ۏ,�[<yF~G	��=��4S�>8xwU�&(��/���C��H-2�ۛF�ڰ��vs�G��l� dRV/�Ϩ`��4�w��_b�d�96r�Y�Ϲ��a�
��]�D��˷��!7��}nI{�m��N1�4��!�<��pX�$^�H@H(�M��)�5��k��unv)�&CGF�5ZA(��µ�v3�둲�yG-�9��m�@M�K��uK�Su���Jw��$]���r���܈��*O���iF�&�L_�L�9{��|�������h��/!+X�ֈOaR�Vk��d���|=�վ�Z�ɿӟ���[���A�w<��r�G��b�#�!yf�d�
ܳ3G��@�E� ?��y۾!����.0�^�F���y�m �Z�ǃp:	�]�J����E��≴ :\o(�����,���-,.����I���+�S���QpE�k)�a��G�g~GY|t[5����W�ڷ��M{�1�"x}�5������r1"��<�N�Յ�5K^V�V!���4@Ƌܼ�|�J}M����^K�������:�@�iLץ���	��X�!GZ��w�{z���\A�����Dy�LM���fNj!N���g3���� {�(*��3��;hYs�pg~mT��0�p� �c�1�C�J��my*��`;V)ƕ���[P��+嗼͝�V96�z=P��N�<����G��NR���Δ��ڣ��U���9޽G8(����n�~��))�Au��5�P�B�8u�M"�C,�]c����'3��%��<��#��o+��m"�p�K�h��'���yj,�+����n��4kN�US�����p���*[K:�t@�7��qc@vv�$�ķ,��92[���i��%�̎�2�WH���(=�Z��7��C[/`������ƽ� /�1 �5w2�C����<�;�"�$��0o�_�'�q�ofh7�m�!����!�l�| `�Q��PR]�݈�$[t��w�+ M�s6)�^�e*t�{/�z���/�pc[ֈ��K������Y�k�@ʺ��{}�?���8c?���5������*_��D$��rj��ѧ����"=^I����UE��rKZ�^����,K\%��~u�H}a�rKI���4��ؓ8$�^ h�U��{U1{mP�4\�tP�s>%��d���G���������&� ��"s�r�W�=�:���������v��(2N���&��
��1Y羊��*�<{��2U�b�b.q?^��F�5`���W�:�?A;�/$��g|�c��)�{��;�;r�ا�$�d8��Y�:��20ב�A|�J�:^z�Mc���L�,�ђLe5*�V-E�{����JB{�t �;] H�t��}���j\�z�|�#�W��Y�+��W�ؑg~��Lz����;%h�(:u^%���#-�H�/�&����sW'%E��!���)uU���}z��r�x-Br�/���3>�G~�5��fTkZ��\@�h+��h`Œ���zo�e�1زI�+J��ѺCP��'=Gn�劒|O���͓�D�u�I��c� �����P_c��/�9	,vM%T���r*��9�)��EϨ��*=#&��p����YA�����zWT����M,*�!��'t̿�;����i�Ui3�{�9dtZk��&3}��ث,�M���=�=�Y�T���ђff���F4�'�����^k3�}�KM���*���NďC��|ͽ�{%0L%gɠ�!��n��w�8��ۣW�@���m��F@��e=��	����$)���V	&�؂	����Nv6E���[�'�Jj��p�>��l���:m��d=����S�Rh�b�0�	}L��)�a� W�&��C�)��@j��!�Y��er�[��1����8\���X�����.�@gmO�W؊������7�Qmx|hL6��2#�lk',��]A5�{Ar"5�pTK��"�UxH0�`��$�ua��f��,����h?�o�P��g�����d} O�8CS8�Ol{�.w�tHo�G�3eQ�6Ɨ�8
ڻD�*B��I�bv0Ʒ�0��b`�(;�78�*�h�5G*E��'z�7�cP�TL%+��Y���6��=��Je21��Q�ZG?q��{
�ф�����>cwٓ�!����0U�"�cP�Օ��c40�������n�������,='|�qif!��\��.(�>�Q�@��0�O�˧j.�N�`��fa�4'��4�� 0^��6ʝ��ڛ��ǰ�O�x\���m�1��U�E.#.�1��C`}�ۇ ��wG��Hݚ�:�-R8�oF�M���ttḾtR�B�-�����{�b�uq�R&�f��5�j>��x�G�+�x�ⅲ]��/s`Gv$��A?�,�"T��s�8fs8�)���3�r�lu�$�d	�R.�jc���O�C� c�l��$%�~#�Z�NR��`&d"�z��~�^=���7��^����fkP8�����!܋�BaQJ��/N��������M�F���im/�~Yl�݊�l��x��ux�W��dF#zk�k@����J�ն}=�@;M��(������m��bZ�A�?����3z�x��/����Վ�L�?5��84o]�{b[ͦ}8p:��6�,Q�'�j�� FS�mM1�R�Qfo��&�k�Ė����a��%���d�4�Mۊ��1��}=����S.����k��V��ɝ���N�x��9q�l�C��-$b�Ce�enc�w:n��Q�+�i�y�������7ha��WlL�T�Y��[�
�_���
p53+#�i����TN�?�཯BH��Ù2V��1�0��ABB�5���:�[�`-ut�3�~�ɠ����>��%Z��'to�Ԫ�ȡ�8���=_�%}K��9���Αj|CypN����e@��'�����I)D�rm��U��'��M\�Ҋׅյ�2R�()������	SU9�������{�)�0'
1a���ϤG��=Ǝ���_c�G�����kd�D���)��;ِ���W%��`�y���G7G 3�y�ڏ�J���%�\>7���47

�<�9�̴=�鄥���]�#7[� :|�EӔOV:�ϤUҞ3��]Рh+.*��)S�@5�`\�f<^6�HŮ�0o�����mkh�oaÜ7	��Rl�(b�E3@<Ƀ��p*��y�����Y'=Y��z�-^�󳼴�Y�V��TЗ*�:��CF�e�S�( �r��M`�Y5n���7PW.�	�>�l�_���Z-`6l��K�9`ȴVЛ4��x*�xB��%'�x��dSKNV8�/���~I�d��X��b2׵nt�Ԩ��qn�/@��,	WO��(�r���&a�ݫ�ks�SDza�7|�>�`[�m�-���\�>L4X�o�2~𳽾��EGNw�ԝr�<�I���O����4d��yw�qJ�9u��[�����q(�6��~e�m2��R�P0mF�9k&��!&�����]�kh�#��r�SX�X����2��
kT��W��cY,iXm(�����&��5dM��]9ںQ�@7�Q3�So:������&^>�2���ш٠qG2������T�.�_��Ǘ���;N�z��+�A9��(��[��[���" �#��B3����=�@�a#���ntP�j�u�&눶�D�8��Cm�n=������!�̸a���L���<�(,f�5A�Մ��{_��E7R,�ʓ���Bf���}ء�j��t%r��ႛ%Й�8�(۵:{Ӣ�(���7�QR��r�B�Ǎ��'�,Kl"XS�e���{��~& n�E�h&!ҹ��~T�i
��@>*� �t�o� �:)�q��"˱N�?�8#��]+�e|��BBR7�-�lٖ��A�T�����>�������V+�7��s�x�/�Z�O�wK�1�Jh_d�Vu�2�P������қo6�ú����[�� ��X��z�<�VU�%x��<de��}�x}!�Qg�AJ�B|�^@�2*��_=������9x��zRs����ս}	��Vy���{�TH(2VA����ai���`�W��$l�.�� ��'����?��������� wU��Z.�0�9sK��=&�|��G�
���u�8�F����A�X�g�T0�.}��&���G��S�+�ca�w'�mo�jL<l-�T ���l�i�s7+� h>���Ǯ>� 3�%T_�0H�R^#�	�G�AN
�M�@��k��k��ꦭ���%2����G�@���gΨbEQ4i:�-6�,»��n�7jR�*j�%��<�cÁ�J�E��)���)�4�Ç3%AX!���k^�k*�Ʊ����Ho[����}��*r���	�~������+%��}ca��"�;/�դ���"� ڦ�=���J�-���r�>��!�~�KBz��� ؉�Ύ�k�k�·�����Q7Q1j�V�nl�0?&Ō%���V阷������׈�?ˀWO-�)��etj}#)յ�{惚���9��>4�mЯ�8z�ZD4����肄�����zn���qz�1f�C
�R'�
W��i�Z���B%W5��'�Ɇٳ��6�{�H��-����$5��>ٔ�""�v��{�̃�]&���/c�@���oכ��
����n�������R�Gg�m�uX
Kt�m�դ����u�ڐzH�t��WVR�R�.�"_~���M��9����zw^}��`��7+�к�����
q�����%�Lq��Y��Tҳ�0�^�}�_"��b� F��Erx����E���Jj�T��
ƥY �����$��F�8~��G(��t7b�:ڇ�:Ӽ̨�z��w?�=�'�V��^��,�0Q�nL��]0�;7d4��M�'���X˽�\%�{9ߞ13Y!@�C~��Z��e�x�i�0w�w��9ܚ��9N����i�fP$z�U��W92<_B�Pa>A�kY��آ4�kuj8��;�r����Ʊ�lp��&��0y�=�aDɁ��h���$�V�GGҟo��0����|�"�%���n5��Q����$'���x}�*)�죏�~��W�K��3���JF����-�,���>/���&zbao�Fe�ʺ0ʅa jE�����[B��W���k�x~Dy���έi��ӣ·�hb"�k��ȶ��&�i�ɨ���L���W���\ ��:@7�	��5P�F�w����?v{�Z��`Ⱦ��h��A��=����-�՗��gx�L��G��t���6���C^����[	wx� ���a�m�o�'���7��@�7`..��S3Y�KÏU��p������\����(��u�����Qά?q�4 �z9e_�)z_;S�zi��	��:~����V����ug�[	�6(�c�N,������3?�\3|��"�/�3�i�_d���)jwY�D��F
��A�&|���}؜�r��~���O�����	��4��]�B��z3÷B<�}ւj��Z�<��bʢ�cӭ�C-���!'����Tߑ3_K�76x����Mg��ݡ�d�ݟ#�Q2dV>b�E��2���!=k=s���k@ ���ϼ|��C�X�������ǟ����33��(Y�x��'�t��|�BL������3��wy/�	8R	����0;�Q1���^���@�՜�$����d&�_�;D���a~�+W�(��a`N��v{�z��r#yZ�Vp`���R)��������W$`�� i�2:I��&{	�#)w�j�z��$܍�~o�M���E�g�(kR�Yg���e������g����g�z�������̶&���,$�gx��i#�'���	Q�C����1�n�=��_���s��g�W�]�mL�/��!.#2ҔS�ֆ��2(-( A�����Nw��Y�F�j-;ھ1��ݥ�0��u��4.���^��y���Fme�#��VI��YZ�H6���S'��&m.�Rd���k@#��Ş�.O�Nz�mh��;)[�N��kj;T�O��o>o�~Q^� ��U��UC��%Pš-d���pei�R���ua޸�����U�p���G-J�|�a�@L���L��)��S�@R>�U;�8hv��r����+���	�C��!7[G�aN�'���Z�A�\�ѡJ�]&�S�!�R���$����h��ר�d��Ǩ�.L�ޟp�@��*v�����g�=��vk��k��1�P��M�Q�p��
��b��X��ۜ�V>!���p"���-��ć�7�S%��k�
��oK�*�@_�`�T	k�� ��j��,�1��;��51��� ,]�N/fE�G�t�<r�Q`M����8���Y�aZ-4��G�k�a��q���/�+(`�PT"ۄ���D�ܔ��vw�М��.A����S^�1�ʫm��Q`J�y��">�nz�h.WK�X2Ӕ��ױj�*�,%0���;��A����l*�K1�V��D��*�E�s1Y���Ǡ���
���s�>e񏕯քHg ������;{�_F��n$�4y�,���|s ��b*:0.�/�6�\~���?��c��S8�;$|���0���s�$}m�%����a����,j����z����%��t́��'����ژJqd�z�@�_}�IW�y�I��a0��-���<��m]Z��s!c^3�����Pa}��s3-��;�:\*hIw
pz��L�nt���Mb��L�qh�e��B�����8b �%�5�&�0��ׅ��z6�� �
�%��H�S�Z��ͦi��\v��(�\�C׫*�k�+��6�C�*���^��+>:�
K�}M	'bN��Ļǚ��f�X/!P����dn��V�eJ�1��X�5��j�s��L\��{
�Ѓ��:��&�m ��l��Qt�p��$+O�D��nr�}V�1��n���ιkQ��r�P0��*��:5���)-�Se`�WmkVi�<�P0�poîQȜD"_�����;b���j%	��
�>X������>��ژ��EUt=�Ӽ&(�/�),��r���e�0 d�5�1D#�D�+���6a���]���8�!p��pb;��~|m!Ӌ�岙��[*:��Ǧ-X窞b^�������QO�1:����)�fR;|�7Qe���I�eJ"�~��m�)
,3:��o�Sp�7V{Ѷ7�7V�'D_���ѐ^�:��������DO�rr��u_{���A4���Mw� h��I��<�+��Y���Ľ�#b^'�pV6X�4�͝�����'���� -O+O�͘�Psڒ~���@�B׷:q���T����Cz�\�ց�q����L�4N<#����&��w��RF{څv'�C�1s�J/�����GN��u��5\̬�U[��u����A�&��g"X�'k��\V�6�M�.Cҗ��-��x����p�~�V��1Y!�g�O[p�eֶ�[������)�Z�Xm�g�/ǘ�E�d� ��q�X��P�ݫ�_KWe,���q�S2-�W���"�t
@$~���P�1�C�=�wxMܰ��@�V�?����ѧl��R���Θ�k�����!��H�y:z�\hh7m�R��`�m��]�7-�sCN2�,uI���ՔW��bǩ�t��Fr>��{�>�0�G.JW/��ۜ%
�6NK��ә��l����	&�t�p�b�M����u��*[�9Zf(��p$9�b!��s��rjˍ�I����LC=M��c�ϒ�Ag{I<��r�p⋑�4н]�oT�M=�6�H�ۜ��ɴ
�����RՓ�k�x�xS!MD4��f�kP�͝���Aw�'n����S��2o4od��"S�\�~'?:���y^*Nɻǟs��<�\� ,��:"x�9WoJ%������lZ ���E�s��1�p�ŕ��:�Z %�3n�U�?��*�ci� e��k{:��(o�[yT<�Rj�QW� �F����l(��gH���2U::C�x�`/\�Ջ����z�&��<��&I�">E�:nIԜ�I݇Jp�}s7�'=϶TY�YX�ѿq���qcH�&(��"���}
_A��w�t�"�ds
�7�67\�Qvt�n�;~�R��Jum����V���P�I�j[h�F@ٻ�Q�H���E�k�f��2PqE�'�ϖ�WI���C� m:��N�
|&�uj0��s�>�g(�r����d�Ƿ,�:~��e�x��h�/���#_i;Ŏ�=��Z|�C��[(Z�����@�s��w	K�n�m�?I����>�}�:J[D��h�F���B��0��#opt��ɶ��{0��0n�kŀ��kkd:m��|�"[ ~��c����'E��c�{���b�~����ҭ���'��74yz�"�̆��������>��Țb�#y��j���ǒ��@�~s9�/m˃�E���7���LXIg2̵�����E�����-=�rD"ʨdH9^�>���0����b�;�[Y��y�9?}4�L �l��Tewh���i�=8��q
w���=r�~�:��YU�S��X�Qc���ko�ܑW��]�Bl�v� c�g�s#P��B�?}ѐ;^�&~.��~�h��rF�` ��J�;�58�b���I��֐��D~P�dZ���`��1�;�'[�{��g�l�e�$���/<�WdMS/��!_j��K���Vz�Q�0bs�ZwbB��r� ����2Gw�������秓'!���4Zh;�6�+j�%��`U �s�W����ϟ�Nop��>N/�Px�^��;'U��KZ,B2�F������_��!$-������H��{�@�
�����]���2�wH��H9����H4�߃؁_ �d628������`$���N��J5��#܇(".X����#\b�xO�9��^i��µ�Ł�������^���xtρ�f-I�Q�@�ז�2���=_����-v����;:1�)�b�'��Y,�\#�ӟe�54T�D�����A�|��B'�pȢ� H���ܹL�3t[%��s�U���6�x��.��5�3"�a�1����<��g��jG_w���AH�df'gj�����|�������"G�K�s��6ɬ���H4. �0�Qw=IE�K<:���3��K�������gc����Aˤ�~��q�5�ĉC=��j��̦�3�0	�@��O�&�
ѫ���M�A����7ͤQ��`������K'��Y�R�l5�Qc��d��b��N��=�O?����Y�y
�sOJ���:A�/��2�%�*j<!�$=�(�N�]`8��� V\ˢ>-�H6D�f�%C�M�<�[����D���'@����Ԣa����V���a`#�~ƥ�n隕�>��C��}�  5���e��I�*��0�R?�V�x,4�V��	���lj��[�\���1��L/�'Ne��a�V&~<�X2�/�{M
B�Pfj�>�����ߏ�(��l:���E˹p�=l�V�-5)j2������#"H�-:*e���Vv��E���\����E�U	��
���]�_s+�і��4�>���lV+Kࠤ�Qӹ�*_xF'��&9��º�t��,�Sef�#	E��S�Q�-���X!Z���T��b�땣F_�eN�R#d����ġ��\�+�x7�ǋ��V	�׭�E�x:T��w��P��]ya�MV���ݖ�>4`?P9<�SԚ�qc!F���6qu\AWg�l��s� ��l���kۑS<N�I)ᖮ���%��� ��ɬ�9iD�#�(Ư��hu��Y ��2�i�̀�rQ�,ܒ�-��f�}ē��}�F�s�I�N��_X��e�n`%�B)�M=����k�ҕ�P�]��dG*ش�n���w��9��cM�,1�;di�e�[��p4?L?�v��E���Ϟ,o�	GoM�
�rq@�or��.{�x̝gJ����y/zrfw8h�Yk7פ�6�=��X1�w�]�����"�v>�0�׌j�4��/Dx�s�iv��;�|��/���G��𳉈��y�R`U*w�|���߮�}���C��U����<�̪���)�@~�ƿ�_���I�H�j�������g���[�¥�K����V�S��vw��KO8�j��õ������W�gC �'��*�1���g\�]y�8z/Q����I���#��9�_VO�\�0S�@XdU`��H6V�l:==>-X�3�"Z�
���`�55Bg�����f�R���S�}>ͳq����C�0���-zcۺ�nu�U]\���-���ȱ�V��J�c˰����߲	��ߒ��e@��oK܏$�)oj3����I�iF��6�Z^�g�L����8��C� �Ї� @��:i�>���+%eXh�Y�ǚ��F�����}�vJ��r�� m��T􈢑�n�SH�چ8�& g%T��ȗLQ<g���.��Z����A)�>|;B�pv$8�S���'�P痌������Sɴ����;~��V�� 3*�PC��Se��
C8��u��_�DTp��HH����\��u�.i��YQ�W�+�=��!�H�ߴ�����s�O�UW�yUT<�M��Ǆ���i���I��̍[$��,`����c^�Q|/^��*���/?:��&�ZG##���8{��ͮX���';��#[vyCc	����cɘ��<^V��E0��Pu�%O��E�S;��&�"/(�Vg�9l
R�3�J�N	*S��f"5�L�6�z.�\1=0r��7pU(c[
)1��� ����費�⌔?ev�K�/������s{�}���g��)���j�u�˧r��BI=�!�:��#�Qr�ce�i�\pV'Z6zm\1 �6�N�!������%z�0̇3�[Y�������<U��g(���9\˵�a��S�N>�_Ó�ޘD,4�?��r�!E��q��:n�Қ2��_�H,�:��꩸[v�w���$�}t������й��R�\�u�\���['��Ba)E�%��E���dJO�3� �t�|�(��#0 �<I	mڂ8��ip��V(Ŵ{�H���,�������$u��Lțx����$WH��6t�b��K���In�D��Ln��D��|�WZ����p-<^��ʣ62�$Ǿ��̈́5��T��8����t^�LC%�E�Ȫe86<o�n�]���c�pg|'	PW��էfa}����C��kK�����Ο���J�)�f�H�"��K*8�;afA�3b;�)��z��ժ��7��{��!رf�=���S�c����]�9��	�-N"�l�j��KZ��v&���jڿ�pgC�=g��u�bE����v�P��D�F��)��h�8���ء�\�D�P���zKL7�a �Yʭ�z ���{Z�0w�}��5 �-�&�����IIiT��g�X	!Ϯf|��'��C�[�a@�鑾����4�q���c�{Q��Z�c��[S���M;����)o$������z��/:Qƛt���8��/1��OW��C4��T)d���XhG��^L�&^h'TDbA-�)���!�N�G�6�h�q�qo� Q�Kei\�& W���7�!	}����/C�>'%Y+�G*N(l���G���(����v��Ǔ�d�WpeXS��E��[u�_V�u�)�T�]W|�R�.�rfUZ�������D8�킌�_���+5mX�I6���n�%8&�\� ���e�,i f�se$9���D2�f��l��)��N�(h�����	(9���Ip��ß���#�1�H��@�����J��'��ēO�eS
��u�]��<Ǥֶ��B��b������iKT���ZS�� �5�\�I7;�!�}�S! �w���Y���yb��2bw��Yއ��~q�R�P��g8�n)�~����%�����Dp�Y��٣�l�}��;�Vs����ܴ�A��x�H=����^�6�D������7N�;���@^J�Zԫ�ٔU��SA 5�
E���	LV�a�@��-!Uh.zb���L-Q���|�k�UP`i�즙�� X��!��yb�FOȘ �!�Q���Q�3k�O=]��3@�:��X�3\�:��#��)cI��q��ɔk�b<�[����ڴ]�`��mrA1�-|X�ĺ3���lߤ+4W�A�S,�a[}w���~���<�<@�lOgS"�K�5��$p�������]	�mY:���D��KP�s�ZQ?��� 1��^�	��r˪SEp��ȝmA ��)�$v�:w{�L/�n2��ű���۴C�j����&t�~,�Z��_G��0�.��P��KGel�^���RX�9R^�$�\�,iS�O+`g�#n"�[�Jx)]d�bJu��GF�L()�Uiֶѐ���]M�"S���`��E��&/k�K�K�{�ܴ��‫㯗x˲W���v@[H�Nت�*���<�X�n9"�������I� �C�3}����dT̲�]����3�]��P������ߞ��+�6tVR��,��V[U�US'��̔`�!�C�������C08Cm�(��4�Y�7��)���}S�;���">���JM)�8l1Pb��&�+Ϙa�:C	��v��D��FW�-�0�ͅ�4�E����`���	 �������0L��ґ&j�b�3��f@4�R|
׻�!v���)90���zE ��<
�z���G��|Ux�&��"s�p�M*��q>�Y�^=c�Z^����`a����9�F{��M-���dI����!��z����`�#�=qԇ{�p��~I��u�њ(v���Q?�ݜ�z)�'�m������[[���%H��};i��7�__�h���A�� �T�5$�����s:�]xX.�^�Ȟ,;���VC��I����_1/$%pk$k&h��=�wBj��%�tC��ت0���#٥Y�>��5+s��\m����)kTPp()&�k-a��ߞ��?��_Ι^��Q��s��J
ȁ��(��F�����g�ϫ�f��$l2���IJ��Ǐ3t��S�D3n���*�o���⮑%w�;e��Ѽ*oY�N�d�7\9���14�C��}��y㕱d1���H���.���1 fN���
��R	�"M.���ʸن��MR��a�-�C�~.�!��`r�x�W���D���Dz7��#w�/T�7��
�x�M�B���C��T�������ˑ����l]�C����j�9���nN["g�>������w�u;��:�V��S3��z�\��T���S\��/o*��	3���ō���3�7AKNZ�ؼ�����/�V���J� �Ȧ8��f<���56C,m���)A��ɲqF�t�":��ۄ���+OYA�K�Jt*�5
�/-��4)��9���!��(�A�������D��t>�c���]3����w�v�v�����J ���Um�40usfdEj0�g����f����|7�85�c�'�[���F�{n��_�PH�o������C#��;�Ea��V�p����١�}���W �@��hSW����j�:�{Z��a;�ړː�L{������F��(��ξ�Ov��Í@��u�u(����p���-�;w/~4�d��m�r�Z$�d�iQ�'OaHԒ��гݜ����]�ķ���)m�W��YL	�0����rxO����9�1i�R�j� tz���/�%A��M/βa�#���U�ci�g(`$.5-�D�b��}��n����MfF*|�ݯ���.%" 9q���p��u m���!�_�k�,�m�'7�ԇ=&}��+wa�W2��UU�㛧%f���p-�"�W�V@6��s�B��M���ۼW�[��*}�	ݥP2dq��(�E��cr�G<�၁��E"���=ƚhj[�u��>���s�9�
���F.��Ε9B"�9�`Yv��Q�a�[������~"��'<P���Y1�^0rtebM�«�Zgc�j��#ۼ�c��@�~�~���辦)zuT.���rݷq
\���&d��?����atx���y��{o�V���$���G���=�~��Z��'Z�m@�3X/U6J-���!8jt��}�%p��N�ԛ����3̪��-�c��H�6�W�� �&�}{�A�ߞ��R��e��݉�v������^	����o|��Յ����=�ʚ�%Ց�9u��]��x�j�D&��UT ��l�5n����	L�9���7���y����+a�<�I���ASy����YG�E9�G����+��9�z�;��?�L� !r�=���b�!z��>�[NC�,FlD2(�-Y�F�ń�?���?���G�+P3dx�̎	����~%��d4PY�ՍD�8�a&�Ad�Ó�6p���sT�oK�z�[�C�t�Y�4�vO_!�VVT�i��G�??�.$� D5��<�B�5�z�4\Ep@��\3��Ü),AN� �����Ŗ���}�����N���1'���N�dB�u����]�8��7Z{%'!"�3{���ѓ���0�"n?w�ϖ����@��
�^��g��q�MI�t��m�)@h����b<e'�Ţ�l��=����b�1�"��& �;> �Y�s^����
��!�TkU�����3B;�	�O��^��R<�ե�E�F��A�,j�]Їs]0Xg���H��^y &
%�Z�� �L�Lsz��Eg�a	�䉜o�E��AEꨑ2��S�g���);<�6[^�{A��`J&es�H�6��ԁds�:�nu�Hg^Xп��3��۞~T�������R�ݮ2YQ�O_�Ssu8�<E�������z�`u����jx�#���n1�
��"Y/�FS,N�J$
���bm!B8��\ �(֓�8�(��Fxܾ�>��O�R��4��Ѭ%����3����%�B,>_�0s{����G�r�D��|z�KL���� ~����vY��<�|kx�b~�?%R: O`9��N���mܔF�s��$���'{�N��� ����	0�^s�uL���i|Es�q��$����]n��7��dj��;\��Zb�� ?�Y�V_\�.�L�Br?I��\�o�Y��,*�b�ŏ*r|7��	�4����T����Zqu�.n�DF��u�\�n�oG�����{hqQ^�n���KA���M���e~��P���i�C���A����%uU�.�/�Vs��1�|E���iF����M��Y�6����D|��m���#�����]؈��;���u���/����=_c#��F�9�I�,s~�V�2���c���|��K�^ț�׫�)%H�?Rxk���q�~�LQH�R�I�7)�g��IW��pj�D����R��]�}��_,�p�h�j�\gy�Jd����m2b����ؽ3�_�(���g^���_�_8��S����ˮl�I��h�ѮAa"hJ��(-��X��c�x"]ɕx����������8jm�	H�{������<ܠ���pA�7�49�j�����<'Q�Vz�Qc �q#�hU�����G�i�b���G���8��Cd�����0�7�*ۜa0s��/<;��J�����qiPpښU;O9R�&ns���C�k����y+Pz�J�I�'�C�y�f�d�{��3�TR��AU�{�T�SJ��[�MacZ)W� ��3	�[��ݽ�8�2tR��R	�2��ynށL��8�c��rVQ�H�u�(����頋E��de�k	GAan�-/��c̨K�m�eˠ'��?�_G�D��DED/�A�K ��դ=9�&�im��r!���� �.nO4ů��	|j������f+Jf���Vl`�e��!�QϪ��FPg{ ����d.��o�p['��6f��|_�d>���Ve�V6�f���֨�3锤��j���EB�iN-���\�0��;#e �l*���^��x�c��&�r9�c0+���-,�$�W���W�ya<Ч�g�kfp#��ȅ�Kt�7�ֲ��f��T�Ð����|���)����{������r��ͷ���.;�$ZQ��y��f
Rx}�z4�x�
�a6��et�{5��i�9+���.>K[7�	��M�3I�4��e+�ٶ���B
2�l�¼�œ=21�n�6֌����lp ��p�.)���z��mEup�^�A1K�c��g�*y]V�\m�KTǉ��N�jȧ3����̷�s�q�^�����]CNhD&����J1IhU �y�"�E��X`��`�P���
6��D�D;!9���/�Z-��4"��;'5�M:+ig3b� 8D��t�Q�ݒ��r�x%�7(N��0{��Z����Bduȏ��_�������!��Z](��hd�P�Uq��k�s��'� �4
��O�20���ׄ��>;�/o�@�zۑR|�l����y���!��e���L�SN��@��όwf\`ߔ���
w��Q!�D�&�BaP2��F��*���Kױ;�0��Zb�q��
G%CP�c����
�M��4�ߛg%�qˌn{c�����˰��lCƢIѐd���r��$D�,Kq���s/���d�+(�ɾ;+U 0�D�ׁ	yE�Xrh�LwL.�����f!�	sWJt����߯��-�(��o_�˝��Q������	o4����#KǲC$�݆�-�o�N��s~�=�뾨�NE�g�TN��v��E I�D?���i3��F�c�����|�)��`���-�cծ7�����HIn��T����7��G$�F�9O?��v  �=w��ݑr3���<׳X%9Йx�KkFoC���!/y��?�kO��!#��f
��ę~��:2�p��nz�H 0FFg��Kj*qϿ���N�h�ªmoM>�f�2;�4qK�7k^��`��u��\�l�=k��1!�;3 4��}W�I�WP�����3��Y�W��u���If��40��д;x�~�np�1���%��v�Å���|vZ��--b��d��	����I_�E�<X�>I�;�v�٢���Q���[P=���M���>�"�)3��YdNȋ�ԝ.'�0�ޓ�������
(7U�_���X�ZF$&��Bɝ$49�"%�8��5�%PC��z׃6�r��a��o[y�4X�6P���t
|0��zdլ�8,>"��N�>R�z��C��d	������i27}8�j_�8��6/��ޔ�3�,]�1�	К���γ~}lq ��6����1���K�5�?@�O`�a�����>�N��h.X��l���Y�=�,cw����of\e�P�,Ť�?�p��G��'�����k������2�#�gt�+F�,�y}���"�"�3d�VY#�5����JH��q�v�R���.!��k�[���n�TRlrL#�-ox�5R�(!!d��I��o���Q61n��"Vh��)	�׬�ѷ�i�b�c/D3̒��SW[S�'9_�,N�������	5�,:֏�)�EU�6�"�$n��T�#!e�7��X�d$�]2C���68�h�z��FB�&�h:fWV��H녱n�X��>U,��6 _Z��A�N=D��/�|��r�;�X��^tqx�9[d�zL���8����8���~L6��f � �7[4��C�	:y[A:�<J��w��-}����(���"�(��y0��;�DG��O�h:�E��z�ᘐ�����]�U���H߼Ң���ϵŬ��fh�������lw���W���w&1�8X��(��ecc4�F*�����9|UQXM���S�E"~�"_�N<��\w�r�����E����Ve���k�e���YH��x~r�8&Ap�ҶU�}��>��q�WY%���~�F���l����n������%7���^;&�H���A]�N4�N���C*ɛ_g�i��X����Z�Y]��d�T$R�f�\�vW�F׽��e_#2���j�Ĭ��}�EcW)ׁ��دx�wN¶�p��zKs��C}���.:C��u� ��[�A}��G,�zP��WK�xvr���D����E�5��N�&C�ҵ0k\�;�m��q�D_�W'6D�K�<eBCQ��(�=WL:K7V�6�Rŭ.��C�'"(7�2E���h�.ᦙ���T/4��}U�nb�J�+핟��Ż�z���Q,4�z1Sϗ�$n4�"x|�� nY�l�R����Sob����g�?I�������x�12K&�c>o7XO�=��JhYCC���[�D�����}"�����!.�ތ�_rh����� >���)3l+h&VX5����-��s�ѿN�Ō�0�|×�{6��j^?h�>��Z��)ݯF5�,��^	��_�b��`Woa�\H��b�^jA�(�xi�C��}��y#l�5�f�:�j���V���W����~����G���|{�ʊ��!��t�ܝ�v�X@��#����49j	�&���zw��ߔ]�c�q~��H���濼�h�+���@�"��N���	� %�p6���M]I�Ǟ�}�Iwm��u��E\vQ����޳n�(�����FӱeiQ%����q�eGn�}����d}��깵�a5A�@�v%z�<�U=0X�`E��N��|�*�JԤ�>g��:��!$j3�9әԮ��u�@�BL���n�(F�C0Y��1ۋ���p�p	�de5�]�r����|����+��4�����4д�ڻFԃ@c�d�w�M�6G�lQI��j6��f�#@��!�ͼ�G��D�N�� :�j� ���܌.`I�G?�T=���J��>���H<����`�g�΄��"�0��R��ȩ$�ߝ��%�M��S�сͬm`��5��d-n��(�b��NU��rl�����e�J�� �L&���.]�D���G��@ƈ8�Ia�^g�x��7n�\0��9�hu:-Œk�y۽�D8��-�i�m��<�a����9��t���v���4<v� �{+��'��`��\�v�'�ؾ/A��cOi�юq-����������e�JM�5�ϫ|�|���m���hv��Q	���S��4��3[�����6c1��$Zc\dyu�����Ggy���C34[W3�H<�O:�6O+�CQa#5^<'�e�tG{)�ՔFM7�������rQ��;|(�n|����y m�m�d-Y�	���Ȧ�
�*'Y��6��:l�x<3}H��-�[�v��|Y��`����Ǆl���~�8�'��w�����D���A��"�7~��b?�G�V��Ấ�{a�,a;P'9��`����"�gJv�򠀄u�K��誒���N5l%�26l�u�{R�C��WkV�-��3�a��	��I�1!�,'Q���?�*C��cۧ,�[I�������_ӂ�s�R�����R?�� H@k?J��i�Lj������W�kF=��o�E�;��_�yc�V���*�#��p_�k��^�&�9,���d�:h�0�L��)1K2��#��e(�zI��޴q4sy&$�*�g�/��*\�
'n�Li՛�H�4ӑf�78<FRP̢t�A���Yb��ٖ}��+�(-\V�V�i����T���0��ز
�+E�{M��-�{`Z�k��5���gZ@�I���]�Fz�pdro�[����pD7u(T$1��ۋ]͒oho��RO�������q����H'%��x��d�✷�%i�x�4Q�n� ���L��wQc���[KO�E�ަ��D8�����rM��? �!%iq�|�Ö��qr0{���DԶ�a�+�� ��6����P��X�<��i�s�b��l����nI�Pj�V5���zq���D^jY)n^^:�k�8�5�8$��ImǢ:���w`0��L��ec[�KcLX����!l/ :!q��$��lI�P��}Y�0~�+�1IyR�7U��x`.�`le��:+:Ynd7U��S8;_���� �\h	o?�Ӟ��:!����?D-;0�AF@�RSo�G�4�s(�WDD� �<C�(���x��^6ePjo��o��<��ަH�;ێXN�+G� �x��2���y���ߢ�ß��J,�X#�m������t�+�_�S4��M&r�(�7u�7,Mv/HG��L�͋�A0t�]@	��]�&N�'�:����O�f���� �K���^%l���Y���1-�u�'��G���&NQ��Q��V �; ��z2dL��E*Bo��}���:���S2�^p0!r�Kj�kf��b���AHK��,����#�x����"Q�AU���S��#J��Ɲ������G�?RL]/Ʈ��J�$��x�� !cD�g���<n�$H��}��2�$��;����x�$=�tD�Iv`�1	C� �!k��yX6��2��[�@�ʵ�k��f�3�̕%��Š���[�#�i�x�0䩥o��pH���Y��^vT�삃j�}�'�1_5���U�;�PM�x#�}6B��]/~��X�=�#�M��N�g�� �l�*Y�KZP
�j�δ�9����LG�0B�Smy�Cz�u��(�����'��B,9� r}屳��.��#�K^3��������v��~z��|˞�e���0�B�_�Ƕ�p?H($�r����h5��%���r��X�A�~wl�O+��e)#�dl4��K&*
��,���s�,Ms��Y�ԠX�^�!���q���t��ѐM��4��vZm����F�ڦ�M�լv	�~� ������桒(�+�]�K�Lьwp=ǡ����ݮ�?*���� .�AjAo�~�e`�44-����?���߫��\��^��T����tz�2�y�9m�h�E�]ڄ�W�NC����魦�Yݛwᗦ'<߄{T����J���Q0ȅ,���M|5䙣������Z��ɨ�_�L=f�c�O���$+F� s)S��z����M����^�PƮ�-ӥ\Js�^�d���A�8_����@�a�0�dϠ���X��Y�;#c|_0���=����{�I�SF�z�d�YMe�ea��ʎG�X�2R�@�_`fmdEc�MZ ��ni`Y�\�k):�2ѡ>|I��i������g�&�b���>������s��#^+��Z�,�,��˴$�@��`�xPY�tv���E׊�ҥ˽p���5��]������̩	g���ݡ�u�u�X|{!<��>��ҷ���*r�Zэ�: �?sۋ�0��K�\yƀ���.d�]m`�ENH�� UZ-��~*�b�����o��UTR|�:���U��d��:�~�Tnn�⮓��o��Й�z�&���)�#q`n�� Oe�#��!Z�zhH����������O�p����~X�"۬>��HƯ���_�E�Q��^
�
�,�Mܲ�A���j�ԭրɸ(W�ߥ�dPo�[Wهo�9���m�n#�c�ljq��_#5ؘ��|:�W�,�7���bwZ���In�9�*{}��-�r�Ϋ�{[?ZE�~����I�*��G���2;eE�F��z:���#h�@�;�;nUԱ��O�ޣ|���o��;�� v,0�<ܞS���N���JA��	�$����U�����z�]s��*�qC����'�J����!�/�~���W*ݜ
[m��ӗ���2�����U�5�od��0s��ff�ef�*葤���&H�`�%C��E6��v@�=7dA��Z�~�D������B*�-�?��Y�3�����Wv��⣢��:H6q5�o�'5�c�ӭ�]K&����W'2s��I)9m�Df�9�3��d�HG�	�͒$��Wb�Yl���R�z�ʹ��pR��fþKg&k�$���hu�4�`�հ�������v;�m���e0W�ڴ�wFM:k�y̍�5G�h$ݦt]��>�8.FUk3�IX�Zb�p�d�I�+����`���;��q���:�����L�����$Ӭ�������}�͙Nk�S8�-�ō}���$F$��aK�1�K�.BS�G��gw$J\*hcA��Jm�0�c�+��6۶ {;�rnRoĥ�P]U`�� �J�n�{�p	�.]Z�<e#��}Lm�6�����$ѷ����"�k��(���,�k�M��!�$[�^-�C��U��D��<����m���U�APM;mj�ت��|�L��B$_,5(ڊ?�N�I�9_�E0��F�+���&h��놠ȴ��<XM������AT��7+��un�K��ιMm�P"Bݐ����+ �s��.֖ڻD��=�(���7Ӿ>ܳm���	�5��Z��:9b:�>1�� ��&��E��<HF/��3>�%�f��h�Q�cJ@݄��r�r���K/Bt*F)�	(�d�,W��47ធ�2���Yی��2�_7��M�'W���8?t��7o�L�hH���jܑ���� ��4��}�J�u�� A~�H]o=('�&�D��T�l@\���p��t�q:��|)�DIә9YF5��fy!\�LԱy��m�af��'��>p'�( ��UY�{����D��yn�b�DF�9�H��ןEuwl����^8�Q��Pj{8ӌ�m�p�o]����C���/�.B?T�"���0d�=!- x�K�����!�*�ObZM! �L0�߽�z�ƪ�V&�e6՝t{�-H�;����T��*bie&^����A'I���+�BJ��&��6�m���-��3�O�*�Yq=F�尛`��Y���B�_���w*9���]r�)�T�!�qS5�"k�̓�5��~�׺%��6���ʜvr|hu����#i��������+E�j|�ݓ���	����O�Sr���� е�~�b� d!!&��DY#cp��6�;[���2�Z�� a0���^_�$�K��Y6��*0Jxs�0 3�{O�R�,����t�����=���ī�3�y�.F��/!���h�{ݻy�SKc�Bov��S��Z#�� s��o&��}�_L��\��"�J�� ���)���v��0<�i�$	�=�I�:�2�Φ|�7~�֙�L
�	�,��M�rT}&��#MRFyB�V+r��ty�`>�_�e#t�mWA��^8X�Pfὰda-LE�NrQq�A����M�zVڹĄN�=��kVб��Íu"g�ΚlM��7��ez���ɺ쉗	rT{�@��.���.ϵ4ZE�i��Sp�<�a{S��_t����d�L���դ�8��+��i�,d���-�0�sT�k��6�v"D�!����lS�#�@�D�ٴ1/`���4�l�<ד�R��]+c$�.�q(��5!~ė��nFd��䙙K���	a�}<Xd���-m$�~�.�HB�$�VQ��O�e_�cH�%���<Bech�����z����g�ʍ~�,0Uٹ�O��@�HgP�
e�	��O���"�\��������9��H`��@��^��q�24�^�D^,��mͨ��e�x�>[-��C���ߎ�^��5<`;��L�� �2T�����I���C��6C=OpM^�qS�/��c&"2(��G�η�"����l�"�{��y�3]�M��~`,�e����ӽ 7`M�)�(��N@S�xZr|��$�f@qm}����&�ԫ� yJ�OLq (��P��̆���9�3��a�x�w�#U�#��Eg��T�f����Q��)t�pڨ�����]\�_���~yI\��P�΂Q�G�[B���K��q�*�#�!�<�������o����1��)vr'v��e��M�_���=_��f�$�F�
q�;���|J�}�WQ�_Ά5��F���=41)�*�z6ET5�%V�j=���(�3�@
Y.�Zf8���Z���Q@�yAב�V&���J���Y0Z�f4�߃��2����;F��_*_#z�������no,FA�g�N�0�����`R%S���y�su�Ι�XXVC����̈s��;�`l۴䗎��l� V�l�U$\v*Q8lN9�m��r�*PM���4i���֧��s�� ��R��u��/qsi�U�}VF��aH)���.P�S�D�F�'�p���mӗO��O��#\)�s��$�B��W���qq�O���t�Q�u��l�q�8e�'N��*�U��VH"%r.ԑ���ܴ0�m��t�fF�Ǹ�P D�6���6�Evv�F��L2�hE��Wl]���5B���&�[�`7,�V�M�Z�����O ��d'+>%�'ɵ5�1�b���EuX� ���?����0�Z��u��-�$� �-�
d��Z�C��ԓ�1Վ�u��T��DG}<�����^�L���������cx�p�@��%� ������=!�m���7�I�vl���1{�Lq���8��8��kiY'��y���8�t�����QKU�@��l��_���ݽԊ�\�}�'����H��m�{�E�70�u����_3�P�wε'�g1�VE���+����͟����Ձ�!Ƌ��-��
I���jJ�<�f^��ȀG���t�t�9{������dN�s��/�Po��}�XGC��ђ�ST�*Ց�d�L���5�%J��`/��uנ�\��L9#DE?�Y/
R��h>��E�C��|v!�S艐����D��	��r�l+��?ݎ�7I߶���o��{��pu��9�L˥g���� �
�3�g����V��<op��j�Nٜ��,��n�+������/�spg�8?Y�w����T�?
c����d� �H����Uz��\qoT�T���Ʉ@���wi}���_�pթ�i����3�!lu�_��Xk?�&��qr���Hݓ�$z	�܅]�^F�Ve*�4���b*�(�d�Mm�7>���{	6H��pH��Ӭ��r��WmXF�|
����u-#� ���*s	E*En�����\!�;�=�Sr8r빊-?�r�W�
0��g�&݋k������������Q����x �n���J�~gT�v4�9�seā.�{��G@��%P���c�Ȝ��~ do����ΨHhc�R,����gyP9�.2���:\��l��ݩH���C}��E7�k�e�k�=�G,�*����0S�b���#������
�%�����_m��_Z�V�3�v2((���ʾ�L��5opJ����Hs�E$��(4%�w�0��0�pt�g��S8��9o#`�(c��;��r�e�??aP��5镪=C[������D�‛���U�d��3d��+6��k�c/�R��d%�¬8�Z���%�"��`ƫ7�1��ӹ((�"�W�7s��AW*�w������8�U7{K�<8�B�E��=¢a>�.���F[��UL��MS�,Ӥ>����4��E���v�w41 �lݯ	��O{����Z
��v%�QۼgY�gN��'�Cq��C��/s˻+5h8e��Ӻ�fcBj^�ܠ��_	36��ĘC�[0ŉj�W�^�`�ı_B%�#X\3Q�-#�����4uU��G����mL͔�.[n��U���Œ1��9Cm������?����>�/Mo6N3Dl��Y��}؜�섖t!W=���Ҫ(�cF�hxSY�f�C��P���H����h��4�A����X�p_�#��Ԧ��x�g"�M�}3=�u���0�^����Bt����@\K��k�>��d'�,�Q�^ϻ����d-z̜��r V+�����x
ڲ|���^�d��9%�EF1����>n�����zJ��+��T2�#����� 7,^)G	��:@97�>����d&��Bf�0��:�\�'����|[���=\�*�ũGl��6���yM ���g�	�����- Ɔ�J^gd��K�.,��UE|���'�d-�[�5.�>�������&O�,��䀂`��ҵ:��r��'dv�#��rC� �&j}��C-���摃��I��3�F��?�R�{47����� <Q�!��Pk)"�綨������8_t��ؠ5�'熵��8��!	4:�w�4�7�~hG���ѭ[�F�k*$_֧.M��Nd�yz����%��@:M����pjBC�²o��H�V=�:r,���G���	�m�ӥ7���,=�,�"S��D�v�����U��Wn?�Z��y,P`n�$�Mu��ǟRc/?�沓֮��k� �!; �b��y_0��F��Q�ؽR⑏ܛL��3�92�{�"H>��:��� ���{L��ݘ;Ʌ�R!��ta+���}�56x�`��Г~�Z�Y�+[�������a����q�|���ªY.�}eBNU��}�g�+���f/"t46���]/߭H����%Ђ��ɂ�$�ހ�(6?��̆T�+���� �۔o�t��:�u����{��G���m�d��)�D�  뉇�'�*�D�ov<��z���!nxvppn[����a�/�{���kԸn�/�U��赾L)�qڎ�EP�6�\<���7��k�m.��q����~h:.z|�I�-��Won�R4u.ch<y�V
��4�����竄
�$���E�	U�gS��O{%�R:��VQ܀a@E
�T�Hh�)�t4�b��2̺���D����+Y�5����=�-�X6��p��ܠ(B�GE}v��[�m~��D��[�n}��D�r5��Zc�@�Y�� �NH��������1O�^eL̕N�L��ۦ>�)
P</����%C �^p	ǹ�De��޿��Z��O<�,%���n������뻨�,�����z����_@\���}g��!������Ϋ=/	�$� 1Qٌ�w��F� ?��^Os�Y�.D���`��g�Z􉘮;=:�J�c���]���p���@���0
t �ܵrx��y�eR�<k��6�BM[�V�Gߐr}^���2��tP��8$"$�^��e�f@�}4bpR]��Xge������=�F�1@�b��v�;\b�"-�B!�Ԟsy�Jn2�D��_k�gP͂ �X��<�v���3�٥��s�j$��R#�.Z�>�9	x���,��>��?�E]�l�5-~%�
Ȗ�w&3����O�-l`-��>e��`�P�	+����zV@�ۀT���f��	��^oޱ/��ߟ��n�y��>{6ͣq�'�|7N�k�^kIN��|��L��1�Uh%�.4?Sf%��H���sG��Yo�)�Ɯ**��[_�,���ږ�V^�����T�ivMf�����&8���(��q=� �!&�c����݆=��~-���WFv%��9�r�Am	a�б���t��=���rf�a��*6M�|�x!�H�Fˡ���g%E����ձKw�/��5\���w/�Y��?)u�6���!�Gƴ���0N^�0�w
$i�pr~d��%ϩ��H��Czd��?�Ҕ���˻���-�ȗ��ѩ���}����K>� ����������wBN�]}�+��?i'x���z�m�l�P�TRl/�����,��?��F�d�IH,��C
��rp (�n�i�ǂ2����ܻc<s��~�~�9�-f��-$�+)Qوv]"�BN9x&�k����4}��C.7C}#.*tL`�#�z�B9s�TG����y�6�|�m�C��ďGm\#�L�����p���_u�R���b�}�����jC4bR4|�W�W^5��%G�n�]��ݭ��ћ��+���B4��(0!��7vřb.Lֻ����u'�`�,�/u����n6���0�<F �rbǆ-���Az+`<#�,����gc�������L��'���R(=�sT)�~��|[X:x��gU�/�ߊs��l�4��� �Ȭ1��8.��%���G�l�7G�y��<�c�`7��R�3U�����\/3�Z{*�f�45�<Tt�6���΁Lm��o�ۺ�`��LZ��@S�c�s���h�W��kQ�j�7����ռg���/X�<���VDvd����
(�h�֛~<���ץŗ��o:���n������� �M6D�����]fAfV�1��gA�%_X���wƆ.�MX��Y9�����a)n�~9e��r�v�z�ky�A&rs$h��YUQy���i�����$���0ğX�	��z����
|��J��M��ai�Y8)N�V��F��{Y��)�X`�6�C�0��sAC�b�;��g�%��	�u�Wt`M<�{��GN�n�⶜�(��fg�����9�P�ozD�z.�?��ajs�\/�w�����c����D�9�'��~Ez���@.ϒ,��E�hwAV��Kyu��H���S5��H����({+�nR;���*?'f��	�H�7R�	w�1��v~5j�^��/�P�Q��dQ��ԄX�骞}��� ��V��@�g��uo�ЖT��Dgo��4����z�j�/W���p�>D���J���; �!�)�dTO_����I����oE�~aN���n�iЬ��X�㝽��l��b�'0�_ȃ�6�Fgot8�L2`�_*4#�`di���D8��4i�2��G���FR��0�þ)�mO�'
ބ���<�S[��m��ʟ�I�":}�~��I4��c �Ť�e��R}@�d���KI&q�D�r���X�W����o��.`�=��4�S���/ֲ52�Dߧ[H�*H��,pp�؂���m�o�ѷCL�;��{*RP��	]�<G�u\ٽ�%�t���03�P/yx��w�G��7a�� *9����튬�Oɴ���<��=���!6e�=�!	|=���~�ӌaQ�ˆiI	�-�=Й�@�A��*��6Y������8}U�k�@1q�˒C�ͦ74I] wdi���]n1LYA��j~��}��h��~��� o���DLT���2>)�$��N�g/�s/0��A�C�����a�.s�M��#`�&�.��j���c�%VeԽ��ol�7�m+�;�/�&ϼ��_��|��L��<�`���	�s~Te��01��j��L�s���Ɋ��~��>���l��Y<D��:�o�dneJ����(�D�i�'z��>��:���8����#]v�>Z�o� �k.J��QV�.=��������M� ��V�OjD0v�A�7��1���n_줒<?s*D�˃�z�m�J�R�q|Sa� =�:�@��[ह�$�2ˁ�Ѫ�6X9^�_T�'ժJv�����a�_K>M�-��Ww'���c (�P�{���Z]�p팻�FAW9����y���\�t�[��T��{�@�b�ώ�ܾB���ȵ�TVPu�-_f�-D����Nu�FM�I域VR���a���f3��bʄW�2����`+�9 �`�����s\	��z1n�>u�̣#�a�eY2���?��J�ȡ�S��> i�ɥ��S8��a]ʽ�IS�0'$�n$����R�������J\�uqxK�����h9Ж�'�x��tɲG�YLU��F⋡a�L.|��ˀ4��~�B��]�O�6�K2?V�3�Ŏ!���B�SՉ*H�)�r�-�
���/�؉���{��-���̓Y�1�밫J��C��õ����s�w��Y�O'8R������*A�qvQ��ʊ�zķ=�����0\$�9���̀�ڪv�=#̓�Ͼ�=3ىD2��U��^DX��l�#���4�)93�$JT�{�B��3��(�+��H}5���Qe���)b>~������<�lur��fp��M�'h\ZiR����R5y�JS���w�lDŠ%4��N��>2�?��[���2�q�~Ycy�ޙ	1�yM��,�v�Ë����z�
 :�#�����n�����6���.!�k�R)�%��}�h�N~��(���2t��i�Pų��w�@L����R�%?X*`io_�3�'TFCDS��� %�<� "$�ZC]���.���׿c�T�!M ��]�4k�V����=Ck_�8�8����q�\�d��/����>,����� GFD�?G�7X�Q��/::rԁ[b�盇��Yҥ;��������<���*���|1o���Wl��Wƪ���^l8�qT�:}"�Uk�>[��˫�#o�=��>\��DT�Y������1�P�w�V��6#bS�.�%*�eӻ}j>Wr����Ri�}f������	}��K��c1�����%|g������8��=���<eC))�U�&�uSo砏�TMWq�A�{f��]7}�&�'._�T��絹������^�SU1F��Ac�_*3���nv[�����a[jGF��^�q���o}f�F[�2tov��0��#�j�{��:s�޼Z�|LO��@Z4� ����l���PS�L������^��FB��]}_(b[�M���L:��C/H�.d�:*΋<��@s90q� |��_0R��BӨ*���qu�*�u�u������1�c�PA�*�	y<�ὲ�f�C��c:��J�]��4rz2,�ʛu�ʇR,"��ɫ������K���w>8�!���)_���]��/O���;���_��zX�v`""��;����@�F����`�>L��(�>�g������>�,`%K9g�W���'�Ib8%�{���g<����͐��ĒZ@6Ҙ--���3P8�[�1���A O����>���5��Aqs"k�&����@:r�	���:iKo�U7����"�&�߂2��
u>2Jǣt� `�E�o�i�UK$S�ė�9S�I���j1��+�2�S��� r����v������Y]\נH1��@�5����!}~B�]k=�Nf��'e��eGV�̄}#QQY�<u�@k������C�0�����P��x�tR�x�P�6k	Bǯ�N��AՋh51j��x�Gӎ����չ����5�9S��V)ȴ���A@�&��3p>'��W/�l	�3��8��?C��ŕ=��F`2i��,�VY�	�k.K��Υ�[7�/�U��q�g�)�/q��B�sg%O�e����I����f�o��95����ҍ7�}�5���-tD�GvO]�s����[�OdNB��ƶ�� !C�Xr4��v�ef�7����ɶS�,Ž1�j&t�x�p��h����~�B����|3{KN 3߮��$��l��b�j� �����7!l�;Ƨ��L�ٗ����h�G��0a�tc�5C(��\�{)e'�2��G����v6�&aa��	�y���ͷ��a��,]��$̺aR<m�8�.��32`d��c|��R��`��t1%�����7[���W���D�65�r��FןrF�i�ֳ�ah��h���LP�Q�;^,�?53��V����*�Q8j:��q*� (�!�kt�<&�����0e��ѷ߾�u�W�� 4qW���R\��+�Lbvm���K�o�����P�>Xn�l� "�a��y�_x�}��nD��9�ۑE��������2,S5�^��!���A9�� �5n��ǆYS&�q���=����5p�g����j���	+C�{E��댐4�z��*AW�(�RD�A�Kq,?��MJ��U)������XM�|V�����&l���f[I}.�wY[��t��78ɢ��v���Ns���Uk�%b���9?B]Ƹ��u2�/7��λȪ�NE��	�J*��|��FP�hյw7����~�'k��w�J8��j-�6�����+1a{!��ϼ��j~G+�����R5߻ru�h���%��(c�q,��{�[�R{L@fk�Ă�D<�����n-
�{�*Iyo�p�ܵ@�E����;4-�+KC����u��`�`.���ݤ��9�$�:-s[�07��t�(P�E��0�Ҕ��<R�$���
n6E@�}�&� ��=G�H�a��=���.�0j�/>u&�5D�+���'Y���"���(Ҵ���5�f�v�Bv1��_�	�U�CLtQ��5�<e���:�l�t����*����.u�/������0������D�<-p�%��KI=�-yx��,T�{��x�e���z�r��l�oư�;�|�Ԩn�`.�M7l��������W� J-"6=��֘[��_v����F�)[�Mu ��#L�:C��ryt��G�d����h/?,���J�CjX�ZO4i�'3�H��Lw��q���m]*X�k=�C~=��/����+�J��=�����pB�'z� -d�=*1���_��2�x
���,��PL��k��-�ը����sO�d����G�[�G DS�sj?s{lB�fW'F��n=�u�`�U�,[��o�{�M$�����_Љ����}�S�D���}�:����/j���"%�U���M�㢄�o]s��V}��Z]"H����O��N���Z`��@����V�wl!�N�猟��K�zJɣn㭀"p�8�+(�A���n��P\�!`L1��"9贰�-;�9�x'%T�������h%��}�'@��׾ͨ��eP���Y��X��j��pO� �&��7k��|�W�,"o��||����K%ys+X����2�"-�Zj]�c�Y^�Y�r��MZ1� �u�0��.I!�(1 ��%eqI��M��0��Z]wN�1��o=)�/� ��$uq9��K��o�QK���������#l]|6���>�z`b�&J8��-��ǖg�%�("i���#���{�Yo3�ˊ9�T�:[�����pV�ՋWᑐ�1t״��$E��_��7��p+�lK�R�w]���;�E���T]��۾�Ҁ����Ǐ>����NXo	-��|v�!*��� �-h����N;;�y��g��Ϧ�w"�6�K�ݻ3Y "0I��۪Pq�2=DmM㣲�������F�y��9Ϣ��1"�Zev�n�q!fN��{	�2sx)K�G�m�P���6���s\�m�@v����Xf�O�^תlyk8�}J}��B�?'����h��`�+|�n��ϼ���nya���)!�W�ܒ�[��������p"����	=�:c~o���� k1�4/x�^<�U�>y{J�)" /V���$fc�.��l�U��b1E��K/�gƍ2*d�Q?HLv��,��-�O�44���}�Q�H���	�S��;���Dzw:����rM��E�6F�xU�mCJ������ɍ �K]����#r�li5F�wZ��Y�����oB���۪��clu�^��t��݌�v�"���3ʾ��p�$k�����/0�L���� ��m�?qG<cGvj u���<�aE��~�S����Vq^`NT: ���%O�grvLJ��L86�����}A�f%�͛�K!�L�β��@zh�"֎��5�|q@,C,��züp&��<�e�M�֛�n�(Y�:m�?z�G/��Y���Pr��|&,L��I*���-�7D�,o#1���/�p��Ο[�#�H�c��������G��0�+�J�Fp	����"Ŧ��iZO�Z"8�sL��d�(��Q"p��0؍yćI��H�v���YW���D	�����'X��b�p��_r'�UMi="����b�"="b�+�G�TU9�vJ<��\����P\��1�~wg�!L-�;��Н-�@�׿=�)�G�DI����i�CM�uӋ�4���k+�����f`��?�؀���F��Z�q����l�K:zSOy����ܧ齽o6or�'�����E��K%vy3r�_h]Z�Ӣ���E�IkrA^<Vm.]f9�_-
������v`��O�;�Ak����L����G��"mE:�I��`��2���q����v�iT{� ��w�[Eֻ(F 9�o
W�K𺖹N��(�QX_��$~<��\�?0d��6L삼ػ��-�9z�rʹ��6eN4�_3�8tP�Љ�E�I�H�r�c�MO��kws��d��k��++6)i�a�	c!��y�qX��/[H��^�� ���Ĭ�z�]�����u�L��_���f���qฐQ腱�)�4l�^QP��4�p1v`������Z�W޼��}�ǿލ
Z�8�/�\�d0/m�l"'~uY^����8K�yӚ�_%I��]�W����l�5�Hac���[@����.��X���(�fR����(L�;@�����Fz{K�!�D�͒�7��}���VG����^��0�A���..Ƅjjo��� m�����H�>v��F#V�;�hh���6pY�����b�^��eL>���&[���M-2f�T;��3�d�9{+ V���Cat�y�� �%�D ;���@Iy'_C��Zq�Q���d[�=�7!�{��M��ݑ�-U�����d��u|��ܡVL#L�ETcn��ę��I�,��~�T��Li�����d��b4���$��gǭ;4�]ޤ5�WV>��J��L�ǁJ'a�Lз�\wiO�gx6U�ZM������K&t7���#fH��o̐�nyӠ�[v�L15��g[
Ӂx6w�5�]���FnC�ER{�0��9ߌ�];��+<�F�o�Y~,ܻ�SO`���k��G/6��b(��Q�/�n8~��%�"���\ߖ��w���vבH�8�{"a�<?8rao������1� ����,���W�{qߋ�ޗ�qΠ���T�a5e�zsn���0x���=�ӛ��\}Z�Q��}��;mV�?�^=��G<�/�Q�Ԕ�3��6�?�[.i�k�%	
K��F({�}YD���,ʕ�dRέ�L�z�u��ґ��-�%{��[Q�VJD�1Ak`w���i��͍͠�"���{���c�]C�I!��M�~�/��EvIM���Ƹ%$*�?E����_�&of�j�^�c&u�����K���U�U,��AS�xd�-L�IVE��3�a"F��X��a�v���Kn�:x�1�=iWm��7��#�3n� ]r��4�	*���6E����>���x����"_*e*iO<��>&�rAܬV(8�����¨2��qx��7�������B�8
M8|����m�f���[#��P�����F��d*A-�XsJ�ʋ$+�"\ 1��<{.�R�ʽ��[������,�D��7�c�%���$��0��4$�:(��	X�9d��be�bP��~�W�'���,Ɏ	~�"�m��3���l���:v��#�N�'N����t\�Ss�ی���x�J_0�&�y(�`�+C�kY�AA	���S/�n��cvX�]�Z#�i���OE�z��bg��C)��5�3s	���N:�85UYD{_�;;���75���i�iTtnNf<�s}��#"3ה�҅C�貒nM�q��Y��MVz�kU9#}v�Zc��ܼ�$�un2�ۥu��rSi����ş�U�{��1_r%h�E8@c��P6¯���5�R��c��;��7�u�9���aM[:���i+kމ8���W���܃!�8	RJ����L��Fz�ὧ�	��K@5�S�vu$y,�/9���9jF*쟰N��.�wfV�PGC��������e8�70��&|�����F|�`.}= M R��E�V��d�2y�BIK�Qoa+����l9RV���>G�\��ד�H7��p�U�].3�WQ�f|'y����@����L7�Jm��탾��a,Z1 �s�`1V���x��Qu�0�z�o��_%��'�,(d�	2>��ɡ(ˁ&�}2Nގy��IN�2������ �%C��l�;��?^��Wx�-�{#�@�E_e����X4$��=�⿔��Ou��J�A����Y�$�Z~d%1��EO)�g���N�L���)ȶ`�&{����|/U�?�3�	��p�́A�G|���1v �8���@o�m���~]%���΂�];<+긭p�X0�}Se�i!�J�~՞�ۛ@�B]
����VJ�ꅠ�0Ld�{�g���/Qi�j[(�ҋp?���r�S�K9GO�g}ĥb�!u���E*I;����^��&B�6lF.H����kY��9��[���|��^��tg�fMӭ���klL�;�.�B�7�����@���2{2S���S.G�Q`(N��{�V�3td����`j؏ ߞ�D�U �߿(�.s ����C���X���&���KNQ�_PC8���v�X7�;�fpƇ�U��Н��D���u%(��i1�TN���AY�!=-/���<@��J�3-:D��x�́#�~�iQ`�/"ޞ��̧��J��^�M�)�0~Q-�=�<򎤛�1�F���l��nS=�'�����V]����Uxv(҄�[�|Z<'�<X���OM�Ɋ�g��W����ZK0P�3������L��U��>�8d,h�S}-�R;4�s�U��m�r�=-�$��|��a�!�Ӕ�]�5�T�����N��\	���`q���SaлMs#��8�4���m+���v0�Y�@<��D+#D!�-�� nU�tdsF��W��{	/ɰ1���b��%�[��2_Jg�bt��brtx��䷥�.�)�˙"X�Iܐֆ�g_B�䙳�3R!�1�n<���V��dLw�ń��z��͗���ݼ�����l[�ЁBR�vCo�Vf��x2��VtC�?������;L���m:B��S;� �=��ۦ$����zot���H@oa�S�R1c��R����U�;XZ��!����[iD�A�����*��W��$� Z���~'�Kʠ�gO�9��p)���4x�]���!���_d��#�?�d��٬י9ֳd(�bǡI��"�q����u@�:�����6y���=��n�k�'�鲏"����������m��j=L �T��5^�:�-Hʀ䉣�~�|�ެ�V	#��5,9�[�E��m7f���ҊC�1�>��Z�{��ù�&Xٌ�()�ʹ�p~���9IA��r�K��Cؾ��`.d{�:���ţ}`��{�^���3Ű���V;D�mW��g���^��0�:D0�}�T}��s:��D��S �_OekK�4�H�%
ΐ����+:t:/n5y�x[���ge�PI�1F���'�FJ�'�de;V����; �����%*��4�>�,��4�_�
�ğ�|�P7kA.^57&o��cB��Z�|G��<	~W�q�;�Z��e�2D'Uy��Hu����v`z��l�x�&�	�dJ��#M���� �5RG�͈?�>,�m
"`�"4����*��YB`�DT��}������ѕ�)��&b�E� P��?�Ч�е>8Cm���qo�	[�ߗ���c`����S�����\�K}��/��������{���c�_�O�rB�ŀ#�#�R�(�i������l�m
��GU���:����u�A�>3!�0T�Q�,�E*5;m�ԡ�7:[,"RM��0˺��WKqCnx�Og�]+�=�䌋�����'C8�l���ɡ#s0��7x(�mk&E��5��&DL�d�:���f����5\���Vh�~;aT͇��i��w!-�*(~��"b$��yLj7}h5o�܄4��	�AA[���%�4��\_�v0�3��-�u�I�.ڗJ���=����ak��ʬ�%CUV��Kr� =�Dػ����խ0��)��Ԥ��h���ĕ��˴7J�Q��,GC�;�ıY�0� n���`6�k�=8po�?a%`�,�d��y��&���p�_:$��eE������?l��p��sX���l���v8&�	�o˹ghdG�PG�d���Z�o�
�����_F�~����A#3�U��<t����X���%[/�7��?��s���W�2>nQ&%�':Õ;[����w`!2|'���]!�<��֭-���ǝ>DȲ�<F`l�\W�Q�Q��L����{�t垰�ƍ��<9@�jƛ��	Y���-z�9��A�,�l��-��m3*�j��_�j�����r���%��.�Z�c�G1�N��p���d��=�w9}�pʽbѶPg�>O8�W�u�5n2�5��s��,�y�n@(�K�nM�8��d ����[���c���t�Q����rR�:��9e fcb�����}-����K���9�q�u���7���(׋v������%yn7�H���O���1���@9� =;m������%:N��4(.)�P��&�ۤL݈ڱ�Ŵ�I	^W'�(5��vvM�d�}���z�͟��(̣��Q��*���9X�q��]���o��~��ٵ^]�W/��8XΑ�w�Z�C�8,�踁T���ɝ���Ҩh���GUk,"��,�+��p�����EN���8F�z�n�zsk��A�!��#Ӌ"��������Ē�_�K>�a�P�
j����_�TfYx���vϼSNwze�7�������n��M9��YM�?���e��� o�q���;����&�3Rr�ah�)AO(�\<�y�,��0�8��ýn7�8������c���j��z�i��t�3X��_��|%��,pP*����E����P	G��̯�SF�#^��Y<v��=H���5N�B&���2��r��:l�S.��f�{���9��(��*�r�ƀ�L�e=�x/���*���cc[�����a���({�K	�g˩��$V�MFF���d*��n:�eV�V���s7@W�[����|.&v���$ʶ��OH���|��f��D�,	@BBA�lE�v2e]~��<�#������A$�8f�e��s�tƴ�P�cu�#'dZ\qC���<Oˑ�~���u��Y��H�U��CXf�F�bɏ�[����^u�PI����?��z��ne,�C:e1=��憠��[�h'��-�Ge�**bw��ԣρ�V�v�����"��=��>������������,cK*�̷XÈ�(�Ս��b�г�/vx�:�,+lbZI��a��_z%��G�p�3 |�"��cO�U��g8ﾘ�훟���w?���t ��A$��?>��	=ߥ�Y:���DjI��ov�$M����b?�y~ϝ��{C(���L5��ր<�t��'pI>�{&C��? 
n������z!gO�4@ ����\�!�j����i	����L�{�g�ۤP�,~��; " �9��7RJ ���fMl�鷀/t��~�!TW��a�N�ź#]&Z��3	ZM1��g�T��}^�`8T4/� շ�='�O��V�w�b��{u�X�V/����W�~��)ԧ���ۚ��V~�T�[�y�#�?�Q���o$}臅#�ֽ	W�_�P����]��j�]
�yز�y�h��=���wJmn{��G�6o�j��=�C�@�i͙2q��Y�>o[�o���<�{DǕ�Eg�\6c9����a�0�_��`�=�RnB��W�������Ȑ���;��7�R�*�7u�2)~��OQ���X��@�V`�>���,���}����ԟ�����>!�'����YL��c�C�����;�4�� S�u����Z8_�z��Ѩ��d��!~�C�B��xs�Cf	j4�w���8q��]⡇_��
6�������������~��������;b߭aI-N$0D�TN!�:He`ܟy�p��4��Pi�p>f����6�!O�R����hE� �����̇$ƕTd�6'�U�����)��0b����I�N�C��I����W��Hc$I!�^�����޾`;l��D%�Dհ�wk��qy}m��q)��/
1,�1���Ŏ��Ze�Z7������}ZQ���e�Q��.��׌J���e<�"�u��"t�ד�H���ű!{�D+�4y�41�Ϗr�C�ڔmg��o�_��dÎ�J���x6��h�߇��o �*��$P�P�{��ji%�pKA\�Ѳ=M�f��Y�PzB���o`���u�w���
�!���g��X�66���jU��/����boii�[<Z|-�'�o5bf�5�|���j�ؘ͕@UT�q#�^���s �:9ۢ1Z�ʫS�BU����Wo���G�� ���Ն��X�
��(u�Dg�L}�L�e��h(�/RYċ�8��H�����z20M��K���/�W�/ߛS�	�O���>���.( ��
�8EAD�v�+83�%ғi�<�az��7�~r��lwE9�2��Ÿ�i��m��e�h��e�Y��{-ɴ$�!���D[��з�½���]�͞Ȗ����A%��'6����,J�M�˝�c�V�z����x�/|Vn���ع���"��,F�Ѵ���/��ɣ{DݥJ-Q�fY�LO?e��K��Ic=5�"m(�Ydc"^>����q;��_�Jل���63=�B��;_�~V& &�G��B�هԾ�U ��Y�z�9���`����!4H���6o����Y������,F�~�v֓���U�I�J;��[d7��F�ip&����� �iT��$2o�����
q���Ü�n(�ZЀ�N�Y�f�"{���[���������E4�ü�D��|�NɳϖL<�yf|�������V�f����	A���\)���BfQP`� '_�u���tp�����	:5�a2 �����Ul����I[vF�C"%>~��8��Z���n�$�8�e�A���4/�>�_���z���r�j�X�J��,g���4w�@=���daXn%`pe��>A
�fΆ���E�ۧm�,�.������㏔.�S����Ӭ���wVx�:�	c���x�N��(���,�zK)$=�np8,�d�C!�1�y�Q��1��V�1�^�G�ޑ�u�a���pl5�Îˉɨؤ�F���H�Ya���
|�^8��ol�%v%d��$b�����B;���kA�#�#�:p:�B|��b�])�&ъ���KD��U����0��]���� -� �]�/��K��1�� �t�;��>���<�l��]����賞�jᙪ�4���ǖRR�d=����X00�F���|�t���݊mf��9ݮ����_y�x�VX����Nێ�S��V���(���M	(dui��;��ڗ-4�2���T��믯�w�z��6�(�;`.ZƸ0����՘5����Wz�%)�?s@��P��P��*9y}Jw�v���,�&5�	�?�sf�i+�u�[�:�&
Nl�g���<�����7Q���0�>}�uoU�2��ձ�Rg� ��Hq6���%m��$��cƀS�,Q@�s�3N�����N��BҶt��co֤���+��}��Y)����K�����:@����P���m-���aA��ΗF�?��57��;4��+��N�k�cJ�KVr����^L�/���f��b�95�(2�A�\���9�c��|6�+v�S\H�P]����2Y��:^���ݻ'T���_Li���Ȓ՞�E���m�f-�[,cle�>H$�XJ���1|� ���j�A�6˟�z���<q��:�R��x!�W�t�B#����3y�+r!WߡG1��D��UN�j15���%2����,�J��d�DL�qt>C&�N��E��?>���y��#���	�ϷM{�E?g6C��zE�a|�$1bp�<�Ľ�[�*�?�{�`9!��e���� ;�Z�}���p�D�(�.l�$�;�$��Lw�����O ��G�#��F7�P�`�%7q�Ʋ�4��B��'1e�j~3��
m�0�����S��>/%����Ĥgy�^y!�K@M���"�|��R2���a���Â�U3�#uj��vҋށP:l��)ZIOw�vR�C��w�&�������ڦ����w�LGS��B3)����Miws��Y�$�z��f}[u㙜T���_e����<� ��!�0`�n�ԭ5SKݶ��D��*�X���B�B���	R��|!���([/�-�B���g�*�c�Ƃ��4��DSglb�Ѣ ��ҿ�K|�+�ҵ�#������b`���(8ҥ��,�z8n����>E�$-�g)R�_K!Tc���K(�j����*io݄���C�B4uPP�G$�m�X��R�K+1JA��`C�q�m�y��|�rsƳ	�}0��P�<�[s����9�E1�L���"E�z g�<��{�eG�6e��"��Gc�me�P��'G	�'{S�W�$ɯ�w����Ƅz�i��E�?V�.���6�?0�8���w���{��M�������}VK�$� �cg�2cF��e����#~�0���Q�\��}9 ����%˃j���,?��|��s�9B5r���+Q5R�*b��F-�������>,��o��$��+�����R$�X���U�+��ڜ;Y�0�=�3X39b?�i�`�'I&(�)��r��,��Z.dfU����y_�o��~#� hYn��l��8BX+Jp%�o�ޗ�����"�cn�XU��bN�ƹ��X ��
d� �k�	�
�k�v<�C�F��D��#��W�!*����-��j�9[	�6�S5n���	�[e|�5�\���"�APl�9Z�C�z�Yaa*5Vܱ����m&�&�1E�Px{�^��v�vL�<1�&SJ�[N[{9�Pu�2�B {pu!t����N9}�F�*V�������b���ͷ~�o���-�d�����������"�e�ߏ���Y���e<����(��YP�Iċ	�Wb~�+��=�)�v����<y���o�C32��&WYjH�O �?�'�VDȸ��������
�Ŷ(a�-d�����jQ��c����ٱT�g�����+Ÿ`X�!%-At&��L5�O�m�O��r��8^UbZ>��;S��-�Rb!��p^�üKz����)��o�|��  a�F�'!�>�o�H[���k����ief������$i;�~�h�X�"Rj�"���Ak�=�D6:w�}`��d�A&�Gs��Z�
�4sF$Yw~���1W����u��a��0�
9�݅
�.���ci�f]�u~-�cfar��Nࠝ�E�at�`*�QV�gq[tv�7y�g�T�/|am�g���*��b�p������T�(���a��vk�@%4Ǔ���v2Ҁ���̭{.{%��[�a�����,V �K�<� Yy����M�h�c�l|�m��%��_qg}�����-��φQ�٨��0yOJ���;`���|��8K�'8�D��D�j��������ޔ!?8�ےtja�R��:�,~e�����s}�\�5Ho��� �υ::���`yC�d�Um�I�%�ѱ}����&_���	�T'(�Һ����D�����xj����{�q�ZS����$�>�z���`ݱ�o,��0����EX��e��Y&7�C��]���z�[/�5{G7��h��TŠ�Qĉ�a��+�ѫ�M��q9�����ع�hmG�ae��X<o�B���'M8y>�]}�BS
�,u"�����A����f�!���U��7����F�Px(7�����r��LL�6"(=�A[�J ��� ��2O���n��Y�eS�Q�F����$�����9����e]lh-,E�.2�: &�>��qX�����c�m�L�K0?;<jL��G�G;�;�[�08��W+n���bXo��?��=.)j?)g����;��F~�I���hW�+;�d�RbV���}V�����X��d�~fp�����O�l�Z&�����d<u�U��HrX;&Xe]Z�<��p��)q�xW��p�k��wTb.i�V1'gas��uRb�t 8�.� ��?���M�/��W�)�p1W�J@Ùm}������J�R#4��`�����,�y-����d���R�����f��M�T!
�)^:a)!�LF��h�b�Rj߉��Щ��j	Ĕǧ��M'��2l�l���p��!s��h���}���a)����!��X�Z���|#5�wE���B�}n69�lAG<�AR�8������h��La�!5*У��^���H��>���9������h$s��*#P�k�y�bE/��0����BxR��yze��vф�d�ݮ�9�]�@��$ŪH��s�_V	y��Q��ݼlZ'2u�,�d��z$�)�A_Q�|�+@���ZpxC�d�R�®G$&!�����D/M'n�a�;J ���
�Mǣ�ݻ��5�5k�]�
�ۇV}�Rb��qO��X��g����<'&�X���&B:�d#��fpE�'i�����IG��A=��G����1�E�b�7�7+5fw�Áw�إf��dS#�(�JW�6@⒒���8JH��E��q2gا	>b�����B�N�c�m9�������TU3֛���@��%�u���i)�o����kS�Xa���yEg��$Uj���:��/�~�^)����y�`V�(�MC�b��P�[���-&�!�֛(����4F�g�w/��r,j�4e�gN���B��/��ȏ2�ŦY�u��W�O�^'� me⼴�LRp�IXW�0!�RnC\��#kg�>�D'���K��F��^7d��L[$����t�`+f4�}lI���r[B,%�Ta��H�Ļ�f��A�ԏ%�2�9��@�=��L��'����\>M{��a3�=�ڪ�|
4��J&.åO�T�?'\}��CX������B�@�ý"��1���N��Ot�۱�Z�)���<=b�Qe!����B��^̿.F&�]���'$e;��=����\8��{�f����\��}K��o���A�JĒ�!;�}
����Ϯ�"���H�]%	{=Pst����$'a���-��(�Vy$�I"ˈ�sF5Abo���cS��[=��q�X�2&��5�����
��r�f�S"b�]�L\��쉺 .�k����X5���KB$�!+���}`�xm��A�ġ��uf����w�W6UZ�Q�JQ�����+��6��_��s����P��>��3��p�
3]�̟e�T���d�z��|�u5�J���9Y������K��g@Pߐ�"�6x����[�,��l�F{�K#�10��l�����W����y6��U��k�vWܖ��<o����o���
�~|�hwO��!��AԐ����nL�Ї�O$A�/�(_��wK�(��$a��b�"کm�/N�"���Af���:�L[���dyH)��hƏ�4�=�5��S_ul�sX���7��ٟܱ��x3�x9���w0�텚ȗ	���Z.F�ry$8��b�^�?B V��xޚ�w�$�*9�J'���J�q
�����.�:�r�S�"I��u�5X_��=��3�6ŧ�hl;����/i�����A<�%[��(! ���R)}7���k�g/����W�0}�B��L�ŭ8E���D\k��
��x� ��o�{�� �Q-ܓX��8�����ݍt ꎱ)G�A�'�
#Q������@��坍$�ˬ(q�����ԓ6Lkz��l8�oX��ހ�F�x�m�mh�8}��d�e瀺p�����(���T2u����l	 ��VT����֛XJ=p/��|C���
RU�$���!��<_R�#�[�?���f|5H}b��z�@�&�
Q����GJ�DS�&�V�d���J�a�����D�iٮ,��t&��2��;T���Y�'�S�?a۲'�� ���d����
�iP"1����߆C(��|#�" ���*��j�Gy��z�M��⫡Aj��Ύ�T�q�"J����H�W˴�nΈ������ь��ۅna�JM7e�6(�������xw�׏�_
�NѾ�E�
�ȧ��Ń������d�Z4A?��5���P�D_Dڂ�� G��esx���z�
El.���'�ᛞg���CE*��G�7���/>e����;R^��R��� ;$���
�:�Z�4�^�_-�9sB����E6;�����rܱ�9[���j��g�ّ�F���p��W�f��f�ݜ}'�̂:-$֏�1iL@eX�}&���!�~�����^��rq�ʹ{��#�+�lB���Bo�z�z�����Ń��3$�ONlqr���=����ƍǲ���_���x�Réu�\�	o����yM7����g;�pA1iR��9�:O\�e��!�D�o���T*Ҭ�t���=��uD<���&b0u�?��3��]p� ����cК����K��;e�?�-�9γ�JX��^cRw�����] U��޿T~s���tr�AS}�3�&IC��<{�n��F�e�I~2;�WϹ֔z��4�qm���,�ە��OM�����d��m1�n��cA�P$���8��@��K�+�����g�4VF[V��%G2�a*#��O����Ձ��ct��mH���vROls쇑[ݚS� ��-&�l��*�H_6�8����Q9���C��
`n�����l��Pd�u��lH���@�#-x
Fw�ץ�a���k�����p�JA@	7�VН�ijA$2��]*�����a`H�~R�
�~�Y�"a�y۩��7�NJ�Z�di�_L�E@��h����q�������������H4Q�D�co��ÛФ���(oN�La�1K�������KF}��~T�W�G� �u� AA�(��Z���Oi�� ���-���M���y�����{�?x"��8��jC��=�$�N�.O�F�Ƶbz�ޤ�����
�\u�9ZJ]� o<���L��W���)7`�Y��i*�cS�.N��.������r.�s������i3�c�t�y�o��x�'�?,��'%�������6o��!��&��&t����a�mm����~+�!�fS)쇒��l��	N�c�4=�j`�Ǌ�Up���t���OkWSp~�Ce�k��5N�Z��Ϙ�Gl�Pk�<\M{�.0=s�%f4�Iw�\�r-n���hpdW�c�&�G_s�s}�(!�hyiz�N0k�`7Vʕ�G��@Y�B
�otҼ�l�MKq�i$!!X;�tbj�k)I������4�_����A��o�|ݹ�1R���*�F�U^נ��?�(��!c�]�>|I�CB��4��>UV_�[T�z�"&�un��D1��+�3?uQ�4d�pDce���9C'sK4
�f��*m>��i�^t��j�C��2�JY�8�'�ʲ�ɠy�g�^��Lطf�(��� ��$R2A�H��K{����.��˽v��� :h�l؞ wX��/�%�#���k�M�}Na���w�π�P�X��&�杞YI c��T�ǀ��{�X�d̶�Ά =xmN^�z��Tl�� �qu�2����0��;�9\s��_i� ��{�WWK���� -�+OD��qJs�J,�n�jh�Q�L�}�΅������,6�����b"6�A����}(�2�:w1��E��`K��'#)�!���{BM�!�S0�>IjZ�hn�O֛��ٟs���^��ү]�q!���^d��w���+�Ag9�pB���Z�n#��x�0ҝ�N�n��!~<���	�{���s=�9l�~툜�7���.|z\��.NQ�O�n��âĖq݋��'�zȑ^�U��#A��MK��'���6�:(��;�u?�Z �����T%��E�k��� ��O��ןS�!s��rm���N� #_���N}�Pa��Z�I�]�˺9)��v�\���,�X��|ރ�#�˴�{:������i��{@�BF�PE�/��N]�}0�o�]�~����ZZȀ�r���Y�@.�H�������w��G'�_*CgBO�9d�cm���r�.@?��(|8|ܮ�����S�]��%3 ����2��j{���Y#z_m����[C��یw����6c�O�]8R��ŅM����GlP�&� d�1wI�ne�)�OL&c�nG*Ν=��L�<Ե�Px.?|��v������`���{��B��������(L� =�9�q..�,���������"����x'�Y-��T�?)�Oo%��m�('����q���R싱w��Ƥi�'Nl��&��ᖻd�F��>�rG��7��#�]㵍����E��$��dc�&�7J%J�{�F�|�-��S��_���|<,���ۯ�!:�7/�e�GI�~�W�g�J�j�\��L�򅍂���C��i�����%�kyP<��;�®dc�s(|L�5��H��׏D[������V����(J�E6
�Y*eo�x�Ѧah����>�5_�8����ݲ���D�a�K�*��2��E���ɒ�@�?���1ҟE��P����Ò�4�v��M۞���O�.6������x27��t����,��1���qΉ�1����|B����:5=J�6��[��S�/�j�_�:�	��5�E����
�>�����ftI1�1[��FZ�$m^��v؋�7����ڭ�a8��*Q�1݄ڕ;�y�����F�@���{�[;
AyY�=����4&ߟ`?��$$��u���o=e�j�Hr���Ͽ&w0����{�5K������:8�k.�FRc";0nAU���h�t��I$!���K�0�f��ԇ!�|J����!b�ٶ8�U�L�D7HbFKu��qr��3���#a\B�=�J����j�{.�9�Z�'��g�E��n7D���ӏ�FΜ��v���0�-/U����e�JӜ�����V��p�r\�A����e���%��N:���o�?`#q���&�p�
���V��a�0���4^���$&��	ti�K�
Bw�E��d�'��s\��h��}�-����r�V��ח��k~xhco�����+��B:���O����6k������d���DנPb���:�����+�{.�7R�D
R�7'lO���ޝ��Xc��.�f}�um���Q^�b���Z�~���@�SN�U�vGkS��������	f饲�ɺ4�%y�$�oQ��A2(�_~����=w�Ŋ&n�U�*�Ƌ���r�2,�R {��q��z�2���(�(rѱa3\���&&��pН��G��_���&�N>������{��$��6+#����'b����l����"%�>�Frv��%��Gx���Z�Ti�ݥ���_d�A�W0���Dv�l���EX��:ik�� �T����⹑Q3�����,}�zv��B+UUu��Ll�f'�����҂�lD�xxao�D�þ���1n}O���݇����U�_g�'=L�ͪ�|��E���%�8�1..T���J��e��Ua��l]��Y��e�f�	T�4!�z����'s/%�[�����Oyc�fLC�3���h�񣏷�Q����-i"� ��e�^� ��ÒQ�4!K$�
ѬK����eczGz���4�ð�dQ$Mbw+��4�s���O^�5j$��IQ�o��أ6�M��P� ¶,�����rh �'d���hK����q�O �%o���1��ܹ�i4'��r]�n��t|����Q8t1�ĉPT�R!�<�f���#���g��y��kmuf|�{Ix%�x�n쿙�����qqn����Bt"w{M`������cv{�T�Ebo6N��|�/��qDu6�r�۵��<g]�b�4YK2���b�{o��M*6�,��hW��u\ݖ�~��~6W㫈�i+���n�YI|${l1l�o�A�1zl��[%b��A�{3�a7d+���w�ҳ#�5����f�����,�ϛ�̕#	rϑ8{h�F�3��3� 5h��,$r�x����G�D�/׮%J9��QN�_۩˩�����[v�*�w����v�9�e�ۧ�Til��x���z.��ܟy�{�w�e�]Q8�'�a����N�(�<�A�����C�C� �L*"���B�V�[F��v	k��9�ɐ��{a�!#�w�:������l���C�.U���k��7�T�p�N��ky� q��I��w	�$�����L6u������7-������X��5���B�ɭf0���w��<�@	�k���j��9���ˠc|u4p���������á&s�+Y��w��	�8��?ut�o�]�E�aI;w�-��!I��]��΁���u},{�߫�P;w�(�4�LE�aZ�#��"�<��[?��U�ϠA�#ĺ�^��K�g��K�˳*�U�U�̾�ܞ))��VٟI�����H�+�[&H��[Ê%�lr�S�R|(J��HT�Ƹ�l9��Q<-�0��-��Z�L0J�}nX��������v\����j�햓u�ĸ1Ă�`d��&؆��h.�ج��>�?n������;}�)Ĳo,���pq����4J���]�>A���5�[`���	h���$�3�g(
�%�;Uc�>#@R��N:�/,:�+���ƌL �>��^��`�'���!�2^$�8��T�ɋ�s��	�J��?���o����-?��y'M��4A��y�|���A�!˛�A���,3��E�b�=ܻ(��+jo}�D���E��u���K���Jl�ېl�i}���oIh=g��������I� ��D�~͏�����n� ����5bD�����E�7A�k-Q��]�j���K�D���K���.�>�����x������+o�����hU��ħC�UԳ~s����,�:2}����m0CER��X����Y8P!���a�Y4T�Z��p�斋�W�N��&oi~�O$�N��e}'k��>zUxSzz�������i�,�ez�M��B�����6�C�������]4DW�C�0�4�����m s����g�h�뚠��	����|�	4ʹ��K�o�	gI%r�*��TT��)�݇���:�]}u����n�����;na]�4E���P�Ԫ���0qq*l�%�`�Ch����z�ȫ�(��U�x����]{�� l7�_[z�V�ۻ�O��gO��K)�x�E�g�0]R���Z���v��:�"�� (�n(^5����-j܆؆"x����d�&�� ?з*�g���PJ`ꊖ7;��M
i�@�ܥ\�v�s���Xa?���j��aH��fB���.>XJ������u0kq���:�m�jv�������/d$�ƍ�Q� *����
T�QX������:��̰_e�����y���~�j�Dt�U�(���|E���0����VP�f��0��P����p ����o\+g�p9��QOv*L<�y�o#������w軼c��Yc.��^c��4�C��#�m�9b9j����xQ G�U��"K�"��kX�@��
8j�L�s�h��X�8�Q��D-'���U_��w=�!&���O3¶
9C�Z ��s�$NN���p�$"k�@�r���/C"�v�j껍g��g�J߃>Ǯ����YꚖy� ������wI.r)���T�+mV�"Ss���)��3�o��\����������� '\ u� ��=�$8�4��@x���%��c{���	O�i'J̜��i)��X���4�1�K��3�2�~`���rE;q��i�ֶo�f�B���;0�����Eo1�1K�钣�ff��΍��2(oH��t���RA�?�G߁B6�iě؇Z�<�.[�]�Y�/A$:����ˁm�^��@�b����P�|s�@.wF���d�HX�(��SO���cN���E�� X��\o�=��HYd��+e�N`k �3~��J2&�4/pQ��܉�� ��1�5l�f� ���Y��(;��4eݻۛ ۉ���FSk%��֑_��8��Bl�Fy���k騂RC�D%m �r�����+�l�p���Ty�j̫ƵW�̳뽅��dEō�
m���i�
8���,Y%K	�8�Š:�l�"�҄��}h5��>l�3,������S��7^3X]@�)�H��/����썶��>,�/��p���~ʰ�당�����\)}I��N�Pv5�r�S�Y\����J��;5���XJ�4Y;[�U� �2�w�f�@�J�0�̤�#�⾓q~��ak�^���?˾QV�b[�0a�1��͗�-������Ei����H��!N>LKpY�NO,�/�6ז�m��3=A^հ$�"Z��Uŷ����
w;�V�U��L��e��L�7VP/��)��X+���<TDt'��B9`�%�����vs�2J��Q��f"���߇6�d��+P����d�`�F��^�yz���A�_�h�wT#�(�СQ��@��<��)��yQFM��:���Z�9i���ϛM��0�I%����fH��s�u� rN��R!�rY�Yt�aO�Qո��O��s-�i����-]b��,�Y=3F1�eAb�INB�j�	6Q�K�SlmT��nJR��8'�'E,�n�,��$Z2�^���a�p�LCI��R�]6��	TխW����=N�ĸ�
���W)PT�X�H @w&5�2����c�J-ff��f�MH�B�.�H�CiD��,����C�n�S$1��U8��IC�iIףQץ�e�c�,z��ȔT�x�T��q"��ߊ	V��J��g�|j����B@3J�<�tIk@����{���"�=`4;�Y��Ag74�\��T ��a){&t�b�ֱn�D��	��j38�$���P`�d�q�3��ҡ���*�B\�@/��뀯����E���U�6�6�������l���v� �tD�C�-�����%�������q����5_�쏲v_��k�s�]�IT�d%<�hLdU~RJ0�l��9��yU���Xy�0X`��C1̕t�w7Bt�����"'k^EW^��L�J��&#�W�d�[��xٛ׀v�%ş�$s�Y�q/}@K=à�Р��q�h���xf�yX^S�i-8���F��C(�X"í/er/9!8Π=��c1�N�ز�ZS���LC3Yǥx0ӠNX����-H��`2N���~m�p��� ���;�����e1����w�ІL�!��F�e��UE��r6�G}���m���7�|=��%��r:вdu]
̦����8���V�zD��L�5��"_������(���b�Л��|���猠`��T%�'~���Ԫ�,���O ޏ��#:.7�3��D���zMW�C�\܅W���7֡况ц��k��Mb�-����p|�i^U�Ǌ[��Hm;i������U/-�,��{C�b�B��2d�,2��v]}�W�����r���M��e@*�$C��W�~��
S �(=7�
#�ƈr3�X�8]LWɲ�����r��<�K�S�s�p�h"C
����i|��^4��?��S�6G���KF~ձ� Dm��4�qw�ϮٯnOX���b���v�(�)wǡ=ӕ5��!�ѧ�I����3«��W	Y��Z��?�/9]s�I�����9���M��17P_��'J]����+y�lſ=���@E�bQE��'�1Z��l�0�²b���X[����y�&g~�xI���^�>ڏ	Q��U���xR�>VԻ"?��ꯍH}���<n�.s�/`���O�8d���E�M��`ҩ��7��c_�{���񤏝��	$��F\3����t�y)N��n�@/�sAJtPEo� ���Ɖ� ��`(�Y���2U>ppjV3F����Ze���@����/�����f��A��s����"e�F;�<���'Xdsj�.f*���l��׵�|F�kg�����]k�Ա�����d �_����	����-FA��|�������4yU�����X�VBQ����	�#E^�T��nJC�9�XO��tȼ�6�y%�AgTMlp"��kPK�ދ3�J�Hu%|O�t�C�xb�OO�I���k��0��Jļ�M�ꆊl2{�������|�B����/�2U!�i�b}�{.ҍ����~ـ�ƈu1 p���c�4��6�+�D_s$�<Z7&���ʞha�gmHQ0�+�P�A�̃~��E)�/�J�輱�R���"�՗�i��]v/���&Oh���V���`��KM}o�]U��I����QXE<�)P	y����Յ�f樂�I�����0'*�]۔�.�~�L���3\��3�)�k0�/�Z#=sv�t����6df��?���[>D�W�U����.F_�Eo���0�~ܢ�}l:}�A��p���=M8�ƛ�T��0q���T��+�s[��a#���q��Vu&WA��x����T'8�Km���I�^FJ5��{\G}���N�0|�G�~�}M���V�BeݼJ,��Q-�|��<5 ��Z}1�0��b�A�d��m�8Y�f4��W_��d$5sN�C�ےOݘ�d��ԔG���]�|8�ؠʒݾ󷦰����[�t8t�7س�>�F�_V/RZn|��-���C�R���b~
b�%Y>̈����D���f|U��6כ�\�7�Z�˴T����[i<ɖ�Z�!b����K���Rd�}z�
���:gw��ߎ��7�簤�*ڕ��o��
Z��0|�`�e�nIOtJ!�`J��X%�����6LhQe\�)����)c�0�`f�85�f�fm�/q!W�����4u�@�$��6{�q¿�>S����}�Nm� ����Yf5�;n���R�l�&�D�s-�ȃæ2��|ѩn�ߊ���c�M��rS%�`�T]�?u��ZW���-�ۭ�7R8�B���(�e��W�ȉ�'a��-/A�/����d����0AkĨ6���N�r�_5�9%�f������^����̈́��L��A�}E��<"��%o�]��(�uz0s�� H�!� �wae�������a�I6�{��hL�D:��F+
�gbE�w-�aEK�%bOOi} �M]�Nf�̵=Ζ"ȷ�g�N�
�����eO�4	{;�W�y�谑~�}��y���=��X��]�JS~釗#8�p�Ok\q�����S������l��$��W���8�A�n`�jL��\�4;(��|��J����d��ܛ͓�5�4O7��
m�0I_M�C����<u-a	(��J���ޱ������R�Ma#�������ݧ��z�8�y�����H
h3�Q�={�PRD����Ŷ��*Ғ��Fҙ������k1��&����5�����4y�Z$@$"O�I���s9d�
w��u\�"H��S_�x�2��1�J��2#��{��C2�'D���rO��0n��C~�߲w�tra��Ęh���Z�#p?�mSP+����xxZ��[F��K���1��-;+��v�'���:�%Mt���ک٩�u�)Vi#��37��Ɂ���������F��i�T!e+�0`	h��&�[����n&-,w�v�IO[1P?��%�[�����ʷ1}�{����h`.3�!(�?Sg����n��N���6*j��#l�|���jBv��ɴ����3���_3�ĸjuDu����&�p��?��%گ
%^%�IX'����C��Wa�v+�?�Z�P�<�:f�{mE��'[��g�v�
ύ�ZQ���������������9]�U�9Si��%�d[���x���!F�(��<�¼�	M���o���Ve6�q
ȥJ�2�*EB]�����۔I��bD�� �4L ��Y�aP%7��]���t����q�_���Z��$�G�]2�xT�1�don�<�Ax��A�!�POh����Y_Cd��+�����/��	,�6^�f�����aH\O>�y���TF�MƠ8��vw[,�R�0~��c��x ���DP"�Ӈ��IJ���[�96��".�BƮ[�?u� �1���HO�7x�\a�LQ�e�Q9b��p/P���r��)+Xi!	�]�r�r�j$��q��ts���oH��IY����Dϻ���5���d�`��oo�)������B�0��] �8<�-�6l�W TM�E����㾼�2k
��ׇ�#��>(�$L�Kf�o���
@W8Ԣe-:� ?�b���w$�m�+�Un�d`|�Y@^T%~~��o�z`��Ґ���OXG�|W_��ap��Q�yc�«�޺"��r��=��S˰8���D��vi�5�.W�$��JF
\Y�Nۧ�A2�4Bpz}��:��$�V�d���h*�Tg�?�{��8
q�, dW��3f#����n�EI����t�*���C�eW�^��ui�g'IG%�x� ������RP"kdV�O�5n��q����2���{��[����� �mZ! ����~0���Wp�c{�DMN6J��F�R��?G�˻^:��Z��"�;�k5�j+#�YI����p8s%�wF�)�#|�|ݒ�׏����`�=�����d$cc f	ʤ�Pt흞F�(X]�0��5 �"5�"���U�˖b�'.2&�&��'`��������#��~�[��iOSV/n�j�L�������Z�6Զ��v����;����zwB�F�g<u>��b��0SCo�|��3�*��l�I��2�ۺU��G��3Y�Sit���e����*,F��O�渕y�!�P|��ık�[�*��D����Il�X�9u#u��/G�f�ņ%�����L�? `�(�O��]��?���y-�E#���OYʊa˳;�O��W	b+/~�`%�j��}5Tׄǧ��O��� p�h+�Ѝ�	/v�3�YÎk����cd;�<��"8gh����3J�B���3k�N蠴�H?�0�̣;ܴ����Dhͱ��}������f�v�a<}�ڶ�`7��J3�g�z1(
l�6a��^;[k(��H��VN�O�X��#Y/�q����䍩-2g��9p���`�^��Y���{\�Y9ӫ�߅���w��3MhpH_�ˤ����Ko�z Doh��M�tW���I�����oE!���%�ժ��G9T�	Wf�S�2ֺ;�ճQT�Ё�%��VL=��]��aYW �c��]sw,��R��M_�>���Q'���,�M�mw|CUy���.�ABy�f��'b�`�7��j�4)��ˆ��O��
�G���e���<�Q>���E2��j��K:E���<�ȸ�
��m���Ǆ}2�h�W�(�&����Qg!���E�3e]Ս�63&��w��\w
W�N�wQ�[��aa	P�7A�}�x�q��������o���wm"�O�%�F�=�~f�9/����Y�����Uw$_��x?R �#D���K��<�����@ޜ�;u�vm���o$4UQjJ���V(�|3��us�M"���&Uߋ�	��皹`��6�Iw*P ����r��k��a�;�JN%�(1�\�<�����J�;�'�=���EL'��@���º%����N��Jtj67�C�,�<���if���+T�+���t���r��WU����s���`z����9�������	��Yٖ_s#��h9=��1�N�^#��UȽx[�wg��@`Vl�O1|�9��o�R톟ib�w�/
_S���[4N��y5�	A׺�1�eP�S*^�
hf�;y��?���h7<�����n?G/��[7� T���P!,�(񩝒Oje^�(��:�|���d.��֚�;���Q۟�S*9����Y�T�]�k[|�$~���==#�P5�����Ɯ���1�W䙝�� �B<]V���z����hw�|����Ҵ���f=���~��MH.�sTl�@6����}�[l�9LO">�4T��SήV� |遞f�L�'�l�sKdZAX<���;c�)c���J��v˷��������Sx�o����Wx�����Q�b޴?aj���KYJ|g�cZ�?3���_jp{]�-�;K�|�����h��.sh�Y�����*�N,��ƣ����'B��ޫ�|�~
N����Q�L�a����YSX���j�{#T�ey\���'��"���3~n�����i��yf0�z�r��D~;�����.G�~>r� �A���r*O�
An��o���j��?�K�Y^�����H�:P_Iy�#����I����1�C���g1K�o��H#48�g�O{ƿ���c��u�е�O���������]Om�.�Ԙ�2"e�;��/�Hl�l��բ|��AF�=��w F��43S)O)�2o�1`oּ�Tl�Tw��J���5D�(�����of(�X+���o�z	��b�z�����68�XqE�<0�Cn����;����hK��JgA�n��z�|H���<�t�H�7�V�׿�5w�����.�m�G%���Z��`k4��)�'/;"��,8-���I��{Z���0&���E���Xش�����LEj�K1��g��S$G�?�]9�M&�=�V�ʩ!׸�l(I؍;�uK��Q�*W/D�R�ߖN]��d2b�_:Aju��1K�7W��c��#Y#$��M������0����1m����<�$���:6���	�Zk�mY8lݪ!�� ��<:�2������s�󤙀�
~�k^m�Ͼ�3�U�	�Y]r/c�V��͵�z�6�ͻP�S�(��#���k7���+�K�WN�1�9x�`.�E�9Q��Ӛlaղ]�!�yO`T{��3 ~V!2��h�g��(�*�n�/��p�ve�� ��޸�ۢ�8�Q�3�p�,����i���x��`���?��/�)Iެ�m}�3�ja/���ٲ��k)m��}X}�nM)����i@�PG�	�~�[xQA�=^�!*k��c�u�޶�@��:�p}�2��;��7�	��a��$��HM�E�^)xDzHe!����+[=����f���{}�Yo�:��rW�'kI� ��
h~L;�ufe(�SKbuX��z�}n�)��� 0��xn��g�*,����>���~P�Y��D �%��9Xw�$K�1�Vӆ��Ƽ��{� h����!��$�\�����/9l#����g�����!��^Z:�>f�*m��Ԙ��Sh��k�Zq�9�:o�����0��]=]Qd�E����	ȥN����o	�Sy	�Q ��'�y�Fߗ���hz��j���$�8�?�֛��#�b����ǵj�xP�k�
UpЮ�a�!�������C�@RK&4޽x��V��$/�r�$ps+�WB����&N�vt	&�Ja��P����g�LO�/��7e�������6*?�G�/?��ǧI,������3�*H��y� '�?W��� �� ʥ����#�4���:�-�GE��|�xN�ߴ�Y	#�l�Yh�џ�kx��`/�b9����m$d"�Df�s�V:�kS��Q�e�r�@�����2�p��}�:�����rV�����5�`k��6~	s,�H{H%�W}eL�*}��:��%'Ԁ���R�V�t,Tf�������>Z^:�~@��ö�S�8a��3gM]J%S�km\��J�ˌ�ȷC���-Vg�#��,�p���h,�g�� ��;�W���*�.�I���_���tr����0W�#ٻ�<(�N���ڿCIn�Ĝ����E��Ʃ��#�U�;>�42EBػ��S%�[��u�h�ӇTZ��9W�o�|�Kz�K>Ԇ�5 �Յ�\\�$�Fq�䛬��ZD�-[���c������޿2���Y�WUS�âP�&��˯�bs��K��i}pAh�٦vTKe�2`�\OFH�ur �a�fz��N��<��9�;�w�8�� �m� ���*ꔼ�ޞ^����C����0|#����8�_����� ���s�ToϹz�IX���}	`�`5��<��M]��5Q-��/�I����8����>�K<�6ě��+�.� Z;����G0�CiʳNu
���fi��t��x!Ad��qg��e;�UJ���J/bQ^mx�s��Ml~C��0����z�j��h8���_x�}w0��ճ<	�l}��S�|�l�_!G�-W5@��WKz�+�֪gA�g������0d� �@�t�]m��VD�bt��?Ӈvz�u"��֫H1��w�=���[��C�	9��6�{_��j�@1�L�]�""e,�*p&�$�t�n�Rr�ۜ����6@?��򉆱=*�	o�I��* �r����R�Zz��|���нM��]�
�����}��70#Ao�L>f�<F�s��U�Z��c��؆�+�p����� ��b��]m�Ҙ֝�r��W���h/�glG�_�y�qK4x�=76�i�=��,ߊ�-ø&�A���
�t�����`�\�5�:.�ʦ?�+�v�L�v�s>�V{KU��sb=�K=u;k����p�)1_��r�-�U�{7$�H	�������͜䡚�z�BA�+���SH������"�$�����ς5�?��q�P�M�Fe����X�fa���L���!Z�4�奂��D�N���B&�# Fm�� ��N�k�\4P��`c��.���A%Q��zV�2s�s�!����V��=�ȡ��rX�	�f�6�m0j@�lM�V��j��?U�aӪB����&xR�+��'p��?��5�������k@�1����6J�V)R���`�{�~ƯҦ ڿ?z�!6�00�]vܕĆ��:a���RUk��`%�Г�ǣmP�;�fl����U �� ..S��	��D��+T����y���R:���z�2/��\�ݍ ��;MFg�����C4H=��ׄ�s��B��#���~_��/�n:Ÿ`6N� �tH�-�;��_��0$t���G���Gɪ��m�ޅ�egC}$�,d�j���X�)I,�&������%V_,L���fJe�R1����\��?(�Ͻ.}&cɅ��9���]T��lΕ�p�����G�-�
'�����8�5+��)v�Y��~"I� �e��~�Ua��������@�=C�9�&2�|lS�7⛮���m%O��'p5�|&�C.Wb°  7��H��+���y,��hR�0ʫ���Ω���
�	��8$zB���+yB�Ī(��t�*z�{��=�1��yl"�
1c�ɫY��\��U�i{Z���������±*XFzf�[R��z�ne��ŋ�f+���jPQh��-JOTT�A���2`��k�q�
5���T���k�����R��/!�[| [u�g�$��a�5�R%�2���x��i9�� �T��Vt��a��}��}�r&�	���Ig�[�u�����6ۗ������שc��/G툠�
 �9�u���Go�myjkG3w�~	0j�����##;�I�b��;o��F���{�rc�˧/xa�m�6j���;���B�*S���2��.�����Vc���ױD��Ht_�{ܐ�?�W�S�г�0<�&C�
�S��I��#Ӹa��B��i��ҪϻZe
���
��y��v8n	T{��R���Ʉ�h�՟ò왜T9p�6l)VUv��	�롗���3�V�w(Շ�X��+�+�	�C�]R�r��J�b-ʷ�r�T$�����`J�{�dR�p�q��F���%�2[��*H:�����;-��O/�E7n�Z�c>�b�K���~�gNq��0h�t������m?��nO��8��o�7�2��֒$�0�ExWfW���)U?�c�oYb`��T�^7M���7�" �.���T(�-{s�B�n���BZ=/5i|,���z�B��Dz	���ɞ<��C�G�Vu�Ūҳi�u�|e��st� �'	�<X�՟*�����+�++� ���+j}���?霻p}��u��gO3�G-	�ֲ�)��B�y���ky�8 �����z�$�6R���"�.R���7��l+⁗Aam��A���fy<�E�g��|���c�`贵`���V=M�P|��o� ^���z �H�ӧ�	!�a�7����ʟ X���8��}q�}g��^j�ph)�ƻ!dx�k���N�4���A�1 3W���Q�!1{��Xj�����,�{���2���מ�2!�k��Ywj�}G[a�S��!�?�*�@��I�c,3n>=<�"���h<�-'����=�f1�!h`�e�=X�O;F>G򽸙�&�0O���_��+^)��ѧ�TgU�i����<kv�(���/��K�����=�O��������k/#�<�̷	?s|}��#����gl����Ŷ�{���W�$"-	�1]��|н�����#�}����;�wi�ңN�
j=�6�vH@d|ެ�Z�c=1XB2�o�"�{9�Eo.���@�˷*�Pk�%����ea#��l��a|Lo!���+�+��\�zWG�+�����')�Ǹ;���fC��kZ�{�*�v�ct�
I��%e9V��ń��/�`ꭝ�����w֢#���fzF�v0���s�F�I4�@��џ��LU��C<�� ���Q���<?`�GQ�^���7�
IQ
�;F��t:�����J+�{���V�%Q���j�����j9�zW��)����8��#tvG��LLFژ��ˏm��kfa�C�ȟ�~����'�X����O� �|��A�1}1I?�׵����-���-G�:���WtD>ɢ���``�h;M��nW����G-XD˵��(���!��X\Q��T��Ԓ����&�����y�>�]��A�'�zb��^�!�̚�'&5��o�v���F�i����B��A_�j��'��l�zZ|H�I��i~�KΜƗt�� ��_#��=��$mb���2�1���9�K�����2�7�F���f}+-[7����-��N:&�g�������w�|��d�;T�~��e��'2lZ�a�Ҋ]aN"͠Nf
#���ذ"��.t�k��_��r3'���l�=��`6�����X�_��a�B<;��h�E��"��Ǳݔ�� �i<�)L�>|ʑ�ךx�%�ЁlE+�����Μd����H����PR��qm(Rݎ�/�rۙPI��m-�h&�@�	��ǂjV잁�Y�	s�g�n��P��Oӂ�tپl�'�R�}(�z�z������Sb=�z{��d� �� �X�	w�͈8���#�j��,5@k��W��G[��9��[���(��,����/�[A �������s��t.}�fsp�`$jHK�^���Q�GEt9|�Ϋ�����E�s��� �C���пN=���i@K阛���1�̣�%��(Y��iFi��Dp�_������p���&�R���w��nk���a,f�Ƌ�����d�lN�a���A���o�C.J�u�K�3.���6>�'�� ��p��7 �'�5�9��s�]�j�"���%���ő-#[l�aDI��&��n-�I�sXD���\M���7�����u�I�n��#�"p^G_�:�e{x�+�in�=���y"�v���ar��b�P�Ӽ2]]��|��=w\�z���'_�����}]�3z�뚟S&���������43�8E�L�9k�Q9�_�U�S$`FtݎQѡ�}N�J��*)� �^�(����P��9;������He1�b�c�����ź�@�*&u�$�46�3�Z���ӎkI�����L)~3�]�=�W���d��B˜C�3h�"g?^~��2<�=*����.���@춍-�}E����_�����������a�37	�Xw'�8cU��&ݞ��+�H�)Ww�'[��!�l"���P9��e���i���X�&�3��z��c߫���v]F��S��ѭ�-��������+��=P���*5�HP%[�-�h��t*"\爹*���j�5f�Gj��(|�:�J�'G�/5�`�\�<��w0��2��i���F����GKH<׈�� ��Y�댼x�a1�1Y��ݪxf��"�~?$�)v�}��&�����HY[«��FG, �;ȴ�w��z�Oǆ�����}x���I�ROU���n֦�� ����'�v���T��A��V�qA"����ʃǽZL�=�i���:�����N�DU� �m� L$̈́�F�e�cA$�J'��|8�!�(�D��L�l(Ԏ�ef�����!�^:[��(�����nK�B�jc����U5/�:�c���_�g�1rE<j�!�So_���g�X���0����]��Jd�����tH-x�Z�Ɯ��D�p����b���1R��d�X7�/n�܏�@�����{J�ʙ�c�IB�>��^����H48��M�k�œ�[��@��	f�-�; ��Ls��RU�\�,J�_�G�֢~X��EV�;�$�G"6$6_�k����@ΐo��4o%qO���n 8�>�j�����Q_ 2&��vuɗ伝|�a��H�'�ކ�Hƒ$f��x���<u)�D���f�z���
�c�Cnضyf���X8)H����m����E��<��\t�Z�F9F�9D��%"؇ �o`K&�	G��DZZ�~�
�>�*��r�Q��:z�^Q,��c�R��,;���`��-`U"�	@VǫmAk��`>��j�e8VJ����Ŏ����V3ko�a�̒Ec3��rV��[�O���o�v̠�4�+
��T �7�q�E��4ky������[m��}WBa�=�
�G���H-.28��fZ�}z^��I�+Ŋ�3+�%,	H��}��R�7���#F��榠mT�4WO���m��{O�#��wf��mV|m�L:��N ��4��Y��7�+$�w}k[S�4�Jy��p�H�Q�f��c}����N9�8�>b��h� q�7o������iJ���m�x�	n[�믙��s,������Xr��/�+I�d���pN\��3�)R��kCR�t��s�ܵut|ǧ(��IlB#$s�3��x �L`.��Qa�#�k\j0Z&i�uK��HC��>̬�6'[���JjV�2G��Vݾ�u`ժ�z�a�0�IeJ�H�l=�q;���+��ɗd��ʓ���;S����R�32@��J��C�(y֥���n��sb{�6�0тG����qX��WL�3�<)�/x��^�J7�
�╁c�Z�A؉�_UuB�:i1���.o�7'�ɪU	�]�BSo��S�:7[T��0#���B�L��6R�n���9P�N��f��y�Ew����%�?�%�M�����{)a}n=�{�!G_�w_��&�Xv����i�4�5��iΈ�[��R	�j X���[S�)��w/ܨ}0op$�ˮ���5��O����^m���騧Qa~vu����F6��)�4�߯�i�T�J�њ�<9l:(5x�	dk�}��2�x���ɨG�Bnꪅ+P��Q��1g%�K� [g��9�)���%��gKE�/M��C�mS"��tԚ��ԕ�}�����Q�G@-�����ˉ����k�a͙1���y~�O�bO�	��`�l�x�`�*iY-9B�*���d}���QPSŒ�NX���S�0��2[|a��]snn+�c�ר��v։��z�M�+���Mq�����&��E���Y�D��0�ݥ'�����9[H`��Ч�~&"���_�|87'Q9�@��sܶ2�<깂��R���/,�OA�W��>�)��E�����O@�#��~e�_۲")Rx@�'��W6�$O��P�B��l&���A@�O�Ɣb����vv4X�m�����l�;�;r�V�����=M L2+;�6f����o�F��l;�s� �0Ĥ��ޛy�%p�9�� �`�?|�D�F�i�-�EDT--��A�}`|D�䁶�cR�:Z�Q�VK����cg@��">������]`'�vx;ZS�p�����s���(��p���|ED�:*�}{���n�"�)��8����o�!��I^�m7/�Z�}��*�ֿ'x�|I�Wʻ�.������ǎ���f���g}{��in�)�TD��)ж��wG��pe�t�J��Qh�x��k�U�Ѡ��� nMr9��̙f��*�^��!��P�''��=���5V�k�`m3�����A�y�R$d���<�쵚Jn,�S�!΢U��V*�&m78�R������F^E�jc���J��f��X��-�_�����oH7��>g��?�c_�܆��GK?�!D�@<Ͳ��XVM��z+�-��$�g6Ϳ���i�4��pPC�x�g�0�b��_.�~������w��@p���~��H�է������!u������y��[3@si��t���袀KP��p�8w�^�k�N�`��å,�W
�w'�_����W�u�,?���A�F7%}q;�#�����&�;I2�?�5�h�Ȋ3z�z���.u��{Kn�:o)��,�Z#!�@d�
��lAy�x���D�v�x?��V�+�XZ�������}�g�&EM���bgQ�x�aH3��՜��Ku4~�{�7ʘ���l�����]P�� >'���/�3�ߺ���'�����,��%���0B-��F����V�5�w�׏�2���ᒚ��򑕠j��c�;'@Xț�T�����I��%O@N��8���>P��J����M8�) �lH�C�zq�sN)�|%����t�f1N=��
ծ��	��=�K��S�|Ծ�!�?���#Ҁ|���6>>T��4/rK�h˺Qs�yjgN�� �Ƥ�k�\��YD^��W��(O�mZ��Ymݬ�P����hEg�т|)�櫛�a�#��ދ�[�trf,�-x<�7n.���l�S<ڔXo�����CꜲs�S����ivF�^@Ҧ��K��x$��rD��PxW��(�[�0���#p�x�e8&�;K��[�!DqФ�>bP_����'�(�g�B�P�Z}��N���.<ؽ�p?��ဢ,#HuQ~�����V�HΑ�&�=ίsZ��N�%�^&�^�C�v�*5(�ñ�����[7���%��r,xO�xsޗ�hC��(P�a&�}a�,� ��~������Z6�w�І����Fc���a�Ӣ�L���D¬���·�[��W�a�P�b��I7��ᢝ<_�NA�=�׌ ����&�=��{��%��p~�`u?�0��Wﲲ`j�3�FM*��^G87��H!N�R6nLxd�r�x�����ND#�F>�1U�/�*�=S	�oiw�K����+GaV �oH��Fm��8=Wc>~��L]��|)k��1Y(Sp�0a����sg�eMIk�ݺ�0v������[3>D����vS�>�~�5u��}��W��hhL��%ߏ�����Jތ�\j�澬a��ۉ�-��h��Ŏ�%�T؋Xhe��][N*ꓞ�=��&_>�Q����saZS��X��C���z/�Ű �s�Zc�S�|�(�~KN�C���Zy[K&��2y�jF6�������}!�0�Y�)3��� �{�T�r�ko
�J)�݈Ε�v?t[�M��صJ�_ƶ��olW��#������J�@.'��3
�Ig���h�ƲT�W�[����X`�Ƥ�8�����)� #Oko{�Q�5d�ˏf}�5<���h�B�w�[Q&����\�!f8\i���9
rZ�����W��`�А�/��A���ؖ���^@�m�4+��<ۣn���5�0��nk�gz����� �Ե���+\A1t4Z��O��R���4�B��a�#�ͭ�!�����&ٌ��P�;nlo)���[��
-�Y1�W���#.�~潨�� �_L. �vq����7pTA���A@����+��Y=J��#I6�.�3�C��1���C�}���&)��+����2$�|�s�$k�〱�݊��~����4yi��l�^�8��(`�v�q��/2Љ���Q�֏�HH�_��_��#��s����
c�99���']1����J=��V�YRRr���p�)�g]���$�3ta��E�+(	��H&��4�h�M�j I���V"��o�'OKe�W�x<�
I�ҝ��0'4�s�U �5������0u�l�� u����>H�9m����(�����ɹO-[朧X�Z_����Oԋo���9o�އl3"��8W�oD58&�$OB��I��	Y��L?U64N17��>F��L�w�+ �%lc�\��R�S����R?�\vĵ�0�Y�17D��k����z.1Y�)���Q�}��%��L�l�XQ1���s�3w�#Cܜ��r6��D1h|�����M�����ڕ�<����0�:h�|��41JѴA�����l/�1Z3+ˣ+E�\����|JV5�wV����te͸���_�R7߃���J/��	�L%6�������z�ܭa(���>Em܄��xƈ��D���Mǔ��<ϛf
��^�ր& �4/0���T�2RU�+�6�R�K�gs3��u ��~
͠�ؗsZdx�ƔחL����g`3.���\kW����8_Ҫw�R�T���z"���Q��X��״ �8�G���I��wg,�|�
�P�$��o����2ڈ�'��{K��"��q���:}��}OB�]P�J�q�$vl����:d�]��<���H_�T�#��U��7t{��r�0����!zC��QFs(���*>4@�s�l�[�xz��e�k�(v1�yW&�0�g�^��}~}]�{b����L����s�H��)�<�'t��+	�ex�#�S�ǂ�PTy���=R�~�Yowox!jT�!z�E'{��o�g�_�`߿P����H^��_�@@S�o��WK��,�Z�c�OJm�k�t�] *�\�����#פ?t\��X���𲅂�S6�$��?T_�S���%w $j����W�W\�fW٣Sh@��qu�gme��"ᛗǽK�z��}��r�ǭ��\���v��/�r�gw�=���D�lu��o�A�:41�����eXa|������8�>�8�Ud�����TǷ.ٮ�x�n���B���f�Y3%�ɕ��x��yV�Ú�w����2����}����S���=CNAzٹ���Ƀ��ߖ�|�Dx�n]�o��ZD�*z��87�&P�),Q��+�ݒ��.�B�,>~.6�]	:8X" O
���
3���G�A�1�;�}�I�T�� �ǂ��C���! ��|-�EE%�6al�Tn6o:bgG-
�,�9�	���Ϝ�N�Q�������ʭRI}�=$��#�slJ(%��C��e袄D�-VOr�/��9@�c��c>���%^�%h�������^h����T򷸾`�����]�8YQ�p͑�v�!�ҿ�����O)R�P�Є�Sr�{M��l<� 4�⧭��:,pzɃ�����!��bP���H��ێ��@oжiQ�V��T|���Lw	�
�$��g��A��x�;p�C���]8�>�����O��<��Mt�/>*F�A���rat׻2��i��L�X�u����l��+jB��ŀ�+�E���ބ`jr��	���I3��k��si��)DlK�zX�{��&�kG��m�o����N�vU�����h����N"!Y`6�j�]8���)��x�/jN��)Nj�gc[�or����WkQ���_�����'7�:�E��~:p�6r�� �_F����R��b~�|ى��%��DOy�dǜ��;�N��
�N���Ac*�$=}��5%��9�]|�=飘uY_2�v�d ^۔L�6����ſGm󓢍?
>��R5A��'�D�(1\[;_�&���>۽T7v\/�p��]���Z�Gj�m@�쩔�)�[0��x��}�? ��������qSW�Zm]@��a�n%�c��X�N�1��-�|�Z�����%����}�a�~T{�:艹]R�j|4R!�^#7�/ᎁ�G� �^M�����7�m�nw.z����v�F�6�_h�����O)Chǿ��j�-�
9r�\�{x_a�g���|���-���AK4�?�m������b)>�\�D��k�Z�
ԏ
LX$#0�ȫ�4'�����쟐�P�6K�AR�L逅9,W�Յfc#����H>�o�q.]Zb_��O�^q�n�2w��z���8��}����uDl���M���8�|ccװ.f�X������>w��4d��|�DX`����t��f�[>��>�"�jl$eJ�Ǜ��QR��];�+Ӗ�B�
���W�/�ʶ�>E�+4A�N��!P�:�wJx�tLK��13�K�mt�ן[��$4�Imv�}}��R�9�%�.���^5�v�#��s��H�`��C>�������75H�@ٚ"����%�*�ߢ"�����4f=��4w�����HA�f�q=a�/�%�v/D��i���G�d� ��F�~��'g&�[a���h�d;Tq1�xv�%�4�T�X�m�B�6�$���p�Y'�	!¶��!*�<��8�.�&��sNj���{�' �h��q]E�tM����^]y�<"��8�شCe�3�~����%)Yx�l,]���	�]��	g��9��y���`H2�������K��_jfB��6�� �Rs�.g�,�}�f�؅�oB��)6I�,���4�s
L���)�?W�Z�o��i�Y�?�L�.�j���ͷX�6E4����r}wCl��~��?(e�������������IQ�$-�I��U��E"x��;���@�t����62>����Ffde�Ƹ�����<�&n+V^<8�f�j]�nV�o�̕�rl�궢R�ч��C�˧�KM�~��ש
nH� kQR͂#��h�Z[@Qa1��'?cPҾ~6�C������.�݄i9�\���Y���%2D�JOlD���v����	`M4=�Y%/v��M�Eo��ύ��u�u-3xF���Y���=�+�^;�ft�n�c�[�� )��N ��~Э�'�PƴB����ɩ�BL�m� ɕ����uT��~M�\��,ϻ�Z=���İ����I���Fީ����m�����h Y,�XOɓl\GE4�ߐ�^�����:k���4��S4�N�xO���`d�'p�cq r�j�U���|HdkN�o�3OQM��`�LP�x�O���R�h-�N�[��7��%֥Ǉ��$+P<��J�'q�<�Q*�����N���]�v�x�-Fr�>��:���s,"m��D�����U�Qh�G��:'
���67~���'�m�=�z�;�0>U!����*c?��r�>���@*i=pIՏ]�v��uj ��ۀ�w��AG��n�.��{�m�bb������e�/����/[�x�M�����\X���:0���O���N�����`��V����t$���
�cJ|\L�����8p N�WK�iQ�&976�̬�k�8M� ��P���j����J�$�'z�F�m�_�e5�x�<�/Y�p938��_dy&~�_����^{�e�)l����4�#+���>1�k� ��]"��#4=F ;�) 
з�����>f!�$Z�(�q�z-��
�M��ǽ�8�ܳ��x?�c�>A��&,
����J��Zq1EP�!���HV0����^�\t�8��������DRJ�'�T����"Ys0�"[̊��@a�Iھ90Z�I^S���v��q���M,��k�5��џ�\��3ZD����B9�K�,�F�SC#����u>�V��z�O���[�{�,�7NT�>:Y��a���y��]�t3��	�J[ʩ
�M����;lޜɻ9���~`�^�)�bpIp�-_�*���6@&ѴUm�vi��FZ
�i��WBL酈�hvU2Ak��/n���ﶽ�B+��-��c�^s�d� ���r7���2u��z�ߑ!��ZiȠqվ(��)���#/JM
�[j���tn���y �b�[�PH/7l�L�8� \�� ��U@]!"�e�"��d���K_�LU�/�8Ҙ�1�����n�h���ǧ��`�!GeB�s���)��q���T�;������6~R�s&�ѱG�S~3E�V˨�k�^CJ��[�l c��`;h�Z�{���n�1��;�0�_������K(��v��Y��Z�m7Ca���^�x��I:"�-�-σԑ�y�^�o�(U��Ml�� �nb�z��X*@�	��ɓ&��Q��Q�����I�ȸ���4I���JS�K-d|�l�j:����l���/��Q�5,�9�<3������39H���&}0t,��w"״�w���0����J:�����c�A>�D@�]_5G 8!�њ��W�<��F�DT��;eO��I��2�(�a�@H��	��!��6��R]	����Y�:���.�%����U L��B�B`}$�d�i~K�o���W[WjZü~�P�c,_ᡔ\�A|�%�C�$7��Aa�����"p��= ��B��z/Z���2�J�ޖ���x�v݈��P�����}C���/��rg-w:�k����򭌫R؞ L	c��W?���>��|�Z���MDF�m��t��m��0�l�{�T.�3�M2A�$��4Ag�i\R���ML�*��ܾۻ�9z��3�~3HQJ�X,fߣoϿ�vSG�_����+*#�y����B�	S�sǲk�3q��m��.�rBy��w1;_ή�
���(����=��	�Ka8�Ty�B5�m%���l�V=�Rm$�C5vID*ex�g�L}��IYG��Sh/������ ��UX	�#T�<����5�������	r;4)�t�Z��F��g\vy@z�D��]
�N���;�S�^�ߡ�������p����f�[\s�r�AK�mrv'$���z��i]D�6�ŖX5M�J��B��i�������k^)ı�%R��E��8�� ��9@B�w�xX��4mK�I��{�S/�˔FJzT��Ҍ��SpH<��:%��Q��v�N��wj�6�s�`>@>��={y�I��o��c�{�3�a21Y�l�|�p'C�p ̅��%�c�f�qu)?4�䜻f�S�A�d_/���2�����_�i�w�}���z{�Aɀ��{�W�m�p�+3���җD�&�3�y�������ۦ٤>*S�-�D�W�fY/�/�͙#�5�N�5��\bf?!8�%0\S�Ta��C����%���2 �	P[����<j� ���&*�w-��<�.����B	��q���5�;x�*���*�!��ޮ��b�P���c�kࢱl�J�6"�=��A�8���g�ʅ�.�#�˳)D߸���}��Y�q!Z�R�8���dL]!ݡKeEHp�T�OC��7�:zE��̨<�>.��˿�o=�y�.�ޕ��K�A/N�����[�h9 ����A�F���[ �tE�sCE�ҳ�w�A�&�m\�Ģ/Qp�7=�~���}����F*�)��{�]ϙ��_2}Q�`p��,F�x��d���jX�;ٽ������A{�ͨTQ*��e9�Q��+-��Cŉ�ƉB��왕�������A���b����5�l��,�'�6��J̶vٔ���V0���s.{t͍�c��8��s+M%�}�x��D�
�]�\��ur��YP!˻3��p����)U/'pߘ)O�݋�o>�����z�X|��Y��&��+9���8�m �}��]���`�Ǯ�����1����Fw�,�#�|Y����8m{|]&*��ŧx:��>v��K �e �,����m�$y߻�Y�Bu4�[�A�{7��?���l���@"��`��u�t���rVǒ­d�fv:��Z|�t��V)]�`�����(ԣ��P+����	����faF�9!�C��޳Z�S�G�<h�0G���A�m����0��d��p��;~�j%0��v�p�n0��� |����&ɀ�)]'�X�Z
�7_FCh�Pul���ЍG��Eu�B�|ˎ���`���� �s��uHt��/���k��z�RH�`��vx��_\�S��~ɧ�.fS��8*'�Pwi�|��;y �-^�E-�E���|�g1�\��������Ԉ�]�I�����Z��}�/0�q��
�lZѓzTA�!��**�'�MR\Ԉ�G9�Б�̩��G��'�n=)�79(^,�=9I����KCm9�kF�1f_�q�|������(;L'g2��8 M���	�\TbGV3��g`e�硿�RZ��)�4�^�5&+��6�o�j?5K�Y��lNT5��5V-��m��X�qS@ Р��Vw����e�ݳ�AT�_CgT���N}��Ζh=�$E�8�Ż�s�[h� `����d���g�Dяx!�qB���I�j�{;?� �K�x�?j�ѭ���q�"�ē���E$	�y�.a��7;��T��"	S����I)����N���驙Y# N�z߰�� ���.Rn�V�B-�QԒ:%@�O�C?]	ƤL������$OK���*�ψ��p1�`?�J�k�x;O�~he:��#��X����t� �ݖ`'+I;L�9����6|K;LNҺ� ���j�N��W��r�z�`�q-vk<��29�Z�e�D�|3�'
��*'�'	/hz����r�*��Pb�������R�#��*�݃Nw�:k���&�������G]��Ђ���Rd�7F恊\���v�=�W;YFy��Q�1��#U��r���}����a�pj����6�u1D�Q!ۢk�ZP�5�L#�<޸�׮�T�cF��}�֔R����-򓲇J���$J��;�S�	��+~n�:#ɣqh�AJLh�<)\T͎���7�����C��f5��m��
��Ǵ�cwj&�Wg����]�����ҼOr!����~NC�i*��1�F��[��Bi���:�O	��ة[_pSI���}�$x�M��'�h��и���#��?��L�q��e֭#0L`>}��M�v����2O���;�	5�(1�k"��W��ne�!@�IOI�0�Q�-��zP`��`�#�j�ͤK1l-�M�	+��bI)wn�^�k&} ԩ�,h���iݷ�;:hT_K�����#�N��K�gE^A~R$�5��i2h�GF��&���ه��S��M�NH3g�Q'VC��L���d��x��G��"���28�$�p-���5:%�J�2׎�ґA����6#���k�K>�|])�)���|4c���E?�)�N� �!��TH.9�Ti��ci�p1)(��C��F�"Ϲ��-kI����8N���#*�����J����h͂)A�Nlȴ�^11P}BM���P���z��'#gݑ��9c�N���㌠"�����z�x� ?z����Ai���G|b$���|�ʃ��ی����*q����鴇'Hw}q��Ў?C�T_i�Y�;oY ���\��Ed��_�6���pU_��T�)���|�E���*�Zp`cb��&2)g�u�лD����0��P6s�e��r!���<~�NH;���[zml��,Vwϋ��ҳ~z=|�#���%�H�n��rݕDw�n1����>�/�	�쾉�9�"����3���K8�G�T�l��qA�Ϫ߼����6���Y�9�h]U2Y��?Y�B�|n����t ���gІ�$�SeO�3CޥK lY\�B��������]�E�
����A��"�9�i��V[j�H8(�,�����-��d4>�)��1r)�.ry��^���޸؁����0�Ce�22������I5;���O5���y��[𓠕���ߦq$6�|���� �B�ҼԆTeq�⍏����z@�����;�!��7�ߠ�*�j���� ���]��t5�`ѱ�w������,a,���K	˛��K���l����!�R��]%6��F& ��Ȅ��3��G2Ȅ�g?���3��#��X�ʏ�5�\�0�s�d�LX�Lfc�j8d��Ub:p��Ny��5x��PK0T��<eK~Z��6�GK�3��,Tw�Q�wwhU(��o�����W�Q Uxv�J}���Ŝ&�C��������i@�#A��h� ?�{
{e��m�@c�p���c ���mN:�v��0�sX��=��]p��t�2�2� ���6��n⟴ѣ���b�pU#��nʼ�*چ���8x�KԺ �C��Z�_��V�i�P���[IWF��}�GÜ6q�)�C��]]����Sƀ�;ͻ��E�����	����@|�����
R.���,���b����� �J!�k]7z�i +�)���W�%a$�wW��lEō�(�����Rg�q�eF~hr^�PP��˔�ș����k%-�R�_U"v�������L��N����S�l�N�\s�����K��.�@I�=��w7>� �蔩��W"�@���-߫Q����S�[G4�_��F�y��=�g��ZX�@/7�������p@�j�$��-�<)�g��&���"�(HfՑ=��?`��{���-�>��|����u��H� �;����;2�:i��
�R!h�B]�靡)�j"�[Xo��mі�	5�?��.�S		)�p�oW���3LI�I*y0'��Ф��F��j��������mKT��K'��j�_�.2�j��S�`>�v��-dZY�]�x\!K�r��ZA��ј�|�1�����-�I��B�9�9�.�{/+����?��Qç��1�/aU���<�'ߓ|bc��#��� ��W�}PQ�Y�'���ٗ}��F���%M�dr ��6�j���A�2�O��0]�3-���ZG��ƟUD�p_���\�!E��J:%¼�z��jy��{�P�D�a_�H�7?�pB���k�h����i�OA_���a�i瓵f�ȳzH�q��$i�7,�J����,gU%�_�x�,&��h�cY�pO�#1Dڔ�� �����6"YU݅����]K���RQ�8�4����x��w�h�@���,v;Y����[72I��x'n�3ԯ=��b���
��_+m2z4ǸL��5�S�KRE!z�����a���؇����Z�B��n��������%2:#�l��'_'ӏ�Ȧ��v?ǌ6�~.�U����u�O�F�M~�c�Tc�k"��I�YrZ���H哮_�:�������Ȃ���_��� ��R��п�#�${�.
����e�xD����W<u[$S�vF^�hgb�h��.I���u�ޚ|Z�k`p2�/�Bw��Yrܰ�v����x��e]����yF4B���έ�L�Ք�zu�C]�Uɣ��� A& @(�ӕ��
��bZو��lF�f��exP�:ԇ�����*ʥ7�-����fY�,��������<���<"����\ciYR�/DE!vU dm$	�e���٫�e�,:z�����H�{��{~*/;�aU�AHN^�eVǾ�Q�O�;]�m�
ͅ�Y�F)���Cc��74'���d癬$�""�j=e�M��vk������Jêael���~OFդ���B�z��?�ټ�6���������Qq� �r���v.��)s�"����w����Dj�o�����zb�mΒ�3�⧍�:���h��m֥d[R��bcr�x9Ȥ�%��CتՖ���XK��?:=�u���M�h�H��'�(ƬJQ�,j�!QftgR�ͺ�K��mXd���5x�V�Js�rf�'~B��0�*2�s>��@a�ă��jW��{����i�1��^1?q��B+���aѽ��];J�8�����()���A�h"���D�s:��Ph<E}4���]�x��H��:��
^� ,L�"Ex�P���^>ۼ�q�W6`��s��h
�e8��m��^`�г�GNyo.b�,�(U.���2�O�m��J,)�9A���B���x�J0an/]=����,JP~٧*�|��B�Y|2���ow�_�Ԙ!�r�3)��d}[8_�������с��A��O-&ڸ��� ��}jbr'~�˕%pg�T�K%虠��iig��LW��k���h������	ቸ��Þ��I��.m,�c�x���TKf��9��3m=ύ�t� �N
�WuU�>��P+c6A�� %�i��$��Փ*.*���S>Q�	[R�^�+��W�����C�As /�� �h�o9�]���P����g^+�w�:C��m�W+�v
��4?m�)�g���/���:��17e�J���RcP�S��@�J�*����ϗĵ;���enS�S[�!�D2#����!�~�]�⬨�����F�sQW��9U������) %,��>�fj*IؔW�k��鮇MD�Pc;~JY�%��-�*��/���0�{��*��o��R���}����oo�H�u"�ρ�2>0�J?2�Xc�k�+�^_7�w�YY�`��7�>r�?p
��kȋ=��+?��ݜ��t��	M�jh�	��"TmG��e��7����4�*O���<��a7����4���O��V�j��9b���ǻI^;�8����e�H#�����S��0"Bd`���_k�����gd*>]h#h��Ztr�U��o؎60�A���K7��ˇz�m��|ݾ�G@�e-9c8UCyW&�h��RR\[4�����5e��=b�j����{�,�	�����*A��_��o��fD�D֥l�\t���?`,���i���+S�-�,��׺��N�B�a�e\G��goP�_����}��i�3\7��{#Vg�w�����jZ~�k�h!iwv����4+���G���ϴU���8&�:�ԚG�F�-	,�3��K�w㟩�NX{�`��`�D�L��\�<$@ tpW�6��
��Z�S^�7�d�:�rUԁ�E���衱إ�o@FC�Z�hY�R?TT�<�����!aߐJ*s���π�cHz{��t�I��hH�_/"c�5h���NDk'D�R�#Ω�K��ӜB	��{���i���e0Oٲ ����T��fLг�㟤t��=�!`��~#���B5.H4b'�p�������k
�i'mt�ӆXG�ap�_��X�oH�x�|����p4q�Sr����~��@���t��Fؤ*W�MMm����H��e�+f&,\�³1:M�����N��P)���n�
��ٺ���'[6�G��2dY3�ޥ�7vڷ7s]��fMb��.9O����)�v��@����))i�WJ�����̾n��x8�:�N��;�(<G\�l���9�������O�$P@�j��QK�2q_�)=�����&��h78{<����iP�+��K��������\�l������`��n�U��M��!�"�\(�5���߷BR����A
�_.0OV��D���;U�Ap�`�����M~��퓳`["'����%r� �$?<-nL��39l8�o�;\�5�иr�!սc�����0�B����3�$����A��'�z�3����S���6��e�x�������o:
�ւ�)�"S�b�*���fw�v�]5���#37ĨF+��i�R;/�]���,��l��E��c�v����2���;y!\S+��.���c5áC����J�n�c4��v��j�w��[�<�y���7(dU��-�����A+p��p�������}�u��p��h�n��[��p�ń�S��[�l�j�i����ò��MY� �̮�W���t+Z�-�� 	-�%��p����g�����D����H�'����
:��+�1`�O�����O�k���t32կ+hV?���6	3��.:\�/�$�:6B�t���wF���P�b�s�!��� ��#����ǲ{�H��WE�um��<T+B�ߜ�1B���~ ɫJ�W��o�6�\��P��]0S 'D�-ٟ�Mk��a��J�o�u:̡B�����F/ilrUۙ�vο��Kܘf_Q�2���ѧv�_NNF��n9 �~k�w���� ������b�g���Q�Nہ�LU50�g���l�p^\`3"9�@R����]K�.U��ūvMJ"�V�3K�=wȩ;��X9�Mę���+,ҴQ��\��B��z�ՙ2U��[�X1+���%:�+W?���wˬo����ߖ�ҳK�|wj����G��-#�����Ծ��3@�U���pu;�2�V9R�@�|�RE���������r�=I� &�6��`){�K�j%����b'�+f�.�,r�1��~�垰�{y}��"�(E��|�?7ȫV(��TZ��5���6�ڸ�/�mNC��y�������^�����p�;*�ۿv���Ї»�n�;������k��;��q����r���Y�$�Ǩ�����L�A��f
V6�J��D|��Q���y&YP+����.%PE%��:��t��G}�C�Ya6� 
���T��khؘ�D`�Bv$ �������F������������7��4ۥVQ�R;����Jl5��,Q����3��a�*��"�Wt�������:����W�<;P�	u.�P}���_
���x m��q29$�lQ����:=J���6/�0*��Z%xh������6�5u���2���If�2�w�zH�0�8J�&�p���e��=�7Iq�-�0�5�IϪY���S�i�WWQH/	gzr*��['a��mgӝl�M}�Q�/6x�#�bX�O�8��F[C��鸰| y�<�;P
�8��ɶ��qU��Ehk?$k��eD�/g�`a��uaۅS&l�6 $����}D�9�f"Z�jP[,gz7�w�����]!oug;�����Mb�X��-���lU�?�i7�qP��e���x�ǋiB����O1	ˬ�Ȳ)ᲊ�����V�0l���}��YXS���ެ��	��{F�2.���V,@M���Q��R�+|��QоT]�H{��&I���:*��- l��+Io��P��T��ڧ���:���k��2v�"�dX�m�� �������Y���s+a��	����I��Ji����Ȕ��%���H�V����Y�mj�k�4S/g�
�.a��hg=|Y�*m^4�S�*���7����h��,�3/���L�HnF����8"R�虱r[H���*���)0O¡���!�L*Rg�k�i"���T8~�����B5�F��^6eS9�7�hЀ7��Q�Ҝծܞt=àu��D��0e���\��K*���Y�u���P�$DLJ}y�+��P7R�
{'K���
�����$�f��l��6���D��k��������7wLhE�|�8w�hfR��%*�N\;��7�r�A�ٰ�а��ŦM7����j6��}
?vi��)�A}9�i hY׎����*������Y��v�g?*�����H��?�ݿT N���
���8숥�mc��0fj���k�C !4��TvE�>?��+p-(I�=� �?�����=�L[� �`e�(�b4ڿ�M�륁 (A���v�n�/wg;�GR���x�g%~^��-P�هӧD��[�H�xno�x�R:�i�P��&:RΔqޔ]��ʕ�J��cƽ|7�����=����Q���m���d��H�Tڢh��8�Ѿ�R&%�co�D�A�Cj�Q�0P�J�r�G3�1!��i�����,���&-�K91kNg7�$�?�o瘲�L%1M���J��w��.ɏ��(悴�#�g�6���P�4�"��AP[Ms�#�����*��D�Ԥ�J�p���0(-h�	��)�zq'cb�K�K�r���@aY��\.��'���j@�o�i�2 @U�C�l�7�#�*�����H>eD�m:S�����P"�E�#�5)Ŧ��,X�y[�Ìt0X�%Aw���#�w,+�tJ8��Z��3��W)�\.	�B��m��|��v`X�u6�(iNGVx���<H*h<��=�~� �����a�v��qQ���6=�ϓ�ژ8'v���~�,齔ΙM�}���KzͿ���ɚ	�.����t��C�d��3��7Y��~���<<�vޮ��P j\��H�׋���M���x���v&��@��x�TU+ =s��o�d�ۛo��s�9��nv(����Y�_酱�t0�V�;f󖕺��u��>�Cmr�����%��N��p����Pr�W��{w�L�oaM�9���=��p\ͯ!��߆F�z
R0�y`��MӺ�"�Hc���L~J,�N��@�xlv����Z����ə���w����\'ޛζ��[hL=5�B8�;���i�5؏�!���6`~�~�^�Y8�Gt:�>d��f�ИP�mU��O�p���ev/�#���EBɴ�>���R�(�^y<�������Z����Y��CG�疹�������x�~�}����VcG75��i�A5��Ф���.��e��a��'88��SEZ���e�F�DV%������r�fi}����}�c/j[�6�yb�`��`���s�8���$T�A����S/�B>X��l�06]vyY����%狝��!,�/tBP�M�,��'��Q�"mN�T�������GT(S|����񞧒�o���a�A\�	T�3��F5.��~fqp�.���i	^F���Y��Aƍ8�l#l�lf�����e�t$45�i'��r#^�F�g-���!�s��U|'�D���?հN3���-	y�V��Z�|�j8�)�Q��!F�r�Pǆ퇽_	�𘴥˽9Ꚃ�Q@-ܿ�w��+lh���_�`��+�I�1�m���u��G�{jMK�E��95�)�D�{C���+�~u6<KËx8]���k8BH�S��K��Ο��S!�zۏ�R��gF�FG��8K��݋0�l�s�S�Ff��N����P]}��=���>�=u#��D9��>����-�Bruͨ#m��	�c��y�D4sf����
eZ��*���tŏVN�zFL�-=@��O�)X��3K�+���Nl�mn�L����2UR�K��?�C���q	��_.�gMbc��y�^�R���fIՋI��S�����E��w�,�V�Õ*W�4n�j-Q}�l����&,{F�O-E�)�֓�h��U��w��e�j�XU�5�S�3&�Yu�[�������-!��+��l�c���\���Z3`踷�-�����d��2l�LH5�Hx�s��v�����d�[�q����"��b� �`&�V��]���'8vZ^_��V��/�yn4�x�y*���w�u�c�6N�%���Y�ZU�YI�{��qޛ
��u�K���q��%�����7&bi���P����9�Rl�0�2D-�+���p��3��ję�њ�
�GuN3��(��������$�O�`�^qYGG(sP��3_R�E�Y�����e,ܥ���=�������vu�3�Ğ�0h~��	�g�,eA���/z��h�w�����H��_۾�O�o����u����H��j�����Je��'u����&Jb��E��}+0ݥ����b�t\W�$���
H�HU��Y&���B�ǟ���A���ݍ�5{.�C�FI�dn��F ۦ :g������ٞ�#� ��[9�W̃A�k�'����f�9Zly����7s'��T��9!C5w�<� )n����;�#>�RM�Ǡˑ���Z���S=$����<��F���XY��.�Wu������$�%��e��_7~z�@� $Pm�;;TT�`{��O��A
(_3�
�Y�c��q�,���N1���p�]����+w��կlZ�	��k���j�m� .����M$�e54d�6���]j���Bx-
3V��Z��Ne�8m���B�+�,�M]�6�|(!h��;�f��~�.�;��uà� r�B���P9wjF楱�\�Ѯ9�J��ѻ=��U�ϼ�fm��gj��@���հ�u1ļ�����׶�ڌ��3ޡ�p���BO]A�G׿�1@������;|i�3��+��`�q�{x�X;���.��O�ҡ�OZ��!�����6��_1o�j��_Z�G�X�E9�J7Pb���:���������2�%�qgUPD�
��5�fz���%�%��=�=lhIm����0h%m[Hσ9��9�]�,~OAv�DE�3�O�:6�3}��%�v�^��1~`�8��z�K�U\�'��@`q�\%i�K�#��=����Oo�4��&���D�2y�iq.��@gz�L��r��4	�[v��Ce�XH)9��4�����du\Z�n��~m��J���~)(�=6똔��L\�KiHt��*���*��i���+�ً�4�~w~
Ӱm�f��|����f���`�}h��A(ٺXҭ��y]�D������ݢ���9�dSL�w0��+8Ǡ�I�h4�Դ��ՠ_ �> b>�-�M$T�s/��͜M�N^dS�AI��o���x$�6K�1��"��%|��1�����	�~ʁj;�
�a��`bat�na�K���h��Ř����}[�-bl��P<=�:Б�_q>@f�B����q���r\^�=��o�$�]�?b�bu��v�)�����H�z��qAM�)�-�'W�q�C|�}T4���qO��lnQ׸qQ[�p�N��o���(���{|��g�����[�X������ɽǅi1����@�M���2�ѵ�q_�X����>5���-m�EG��Bx'_��1�G�{,Lؾ�p
3����W��j�L�R"���/��i߉+$�AR��,�	'�z�d"�GX��#H�zL���W�`��٬��`7j{���Q�#�[У�W����F��و���ʁ�}cb����$��!�Lx����9�(�.��D�� �0t�q/ْ�k�aF�-7�K��� e�J��z�����Yd2�)aq[�XRm �>_zNٞ���bZp�����d;n�d��{�A����h
��Y�A.^.�&u�{Kc����i���n� �}�]'�=�r�H�`ET�X�C<=]z�*�t�>@5��"(�t�+�72���Kǖ�ׂX��
+	G��Y�6-v�2%��!�VH�ٽ�t�܋|���+���;Z:{�,��?6�.�m��)���L���d(p�Yd�q(ZnΓ.��*Z1�u���t�IҬ:ξ�MNv��70����Z��&m�L�������wi�gsΜ�I\|��Z�5��pn�l �X������{��J���R���Hf��g�#��>W�bXɄ�z|�����r��nuK\���>W�B���9T�.�w���*~��`h^׻�W�b�ۺp��+��=d�l��V*p.�������3��jTW����	�o>���d$�jQ�MY����~��G����]�T�#���Y���)g+~�Yo,�{˾��ܫィ�b)n@���]0�X��z��! [d6�������?�dE e=����Z��V���+,�.v�,w��\��1���<���J)E�Eb��^�<�E=�.Rhza����*+8��C���S�*Rr�
i.��w��}�@L;�����-s���t^��bnJZ�?*�,��cAs�z	��G�Z�v�աq
��L$�,3u�v�	��P�_:��Ԧ(~��Ï�����X�ݣ������y�+����&��
=��#go��y��Y]Il,Sԏ���8���;<�O)w��h�ڽ�H����(a#z��(Ւ$�������u�E��倂�z�x�x��<����伔�p�<�w��\�Ǐ|��B%��Z�V��R`���<�n<�+�ۋ�j�S�Cg8$�������KƠvnT7E�E8hS����-T��c���N�?�!H,Č��"������Z@
�Nm�s@֭�-*t'U�8v���6��x��gޝf��������_M!A;���V�x��3e�:�U;���퀯}���h�۬�|�1ۡ��9��G����R1�M�6S�'������[��v��pp���N`4�l�������ڍ���6:��cW��f��u���.��7�,�ɍ�9������f��}@�H@�w;/*1K�ڤe�Y^���d�bx%���蟑��/��0XDR��q�+1��D������u���
;��p��xO���u�b����r�0��X�jrc�<�Ύ¤"�INmR�0l�?�N�L��>{�4�� �b��g��n�����bB5�8��1�@�a�\��	����*H�=_�s�e��nQp���˯���ʈ#2r�=�����様-��EZ�%��N�mԊ�i��@B|������$���Js-.XΈG������<N��kb�2eݠ�s�}�x,������wl%�5l��|����HG��Cb��]ȊF07����셵��'[�'Q��y����S4���0��&KϾ��[�
:�1�AҠ��E-]%���;�H�>�M�A��#��[!��|�P7Q&$�� �o3�ih�9TPT�k'oNr�v �I��Q[��e��Y���Z�DK�چ���E��.� @���$&v-JAрo��^~��l,�!a�3=� Y�A�<�k訶8��K"�G�;���H����n:?�C;�����s�����c��6�qƒ
|B�&h�.]&ݗ!��ܻg�
Yw<�����(L���o���\�&���a�k������-�wJ���� (|f�'��z����@@%Z`�I�(���Wf�Eb��`?K5��_�-f����㰞ͽ�EU�k�#�̡ /s�(���F^����~O�8��_�ԍ�7Dx}3�f��v��6�N�?�ap07r�����)6�7�n���7�c�H�����rW?l��J΀�8���ਜ�" t"k�)��lޚ�w�����"�t�Y�K<� C�ՏP4$�hv�O.V�Z��1��{^�	�#��ũQ��B��q/X�?�<ExG59�4��=�<�2�?��8�Ð���%�=t��wq��Y�IM��#"��bܘ!���3@;ἄ4]Mn����lKq5��ӊ��9Ѣb��KKZ��!�����H��W
	�����r���.���k�8�޵E.S��d�a�B��L*�"SJ�~���WĆ��LK-wц�Y*G��;.���9��WPrn-���9�+@��c9 ��+�O"�z=~"�F�:��~�������MO���hT4��� mػ�@��3EU���D���v�R��'���ц�;�E�;51��0�Iܸ��ѯ�~����g�pcMd��\7N��)8�`;��� ѫ�.b�����+e�j���M�13�:�!�e*�N�͒� c�<�]��(�+K�����*Bj��>�A7�۽�r�I��&��&x�Q\sA���;|iuϝI��? ���^kM�`��.���7��K99o��Fq*�c2��q��yA�
#�p
1���PoţbĞ��S-ʜB�h-y���J �͠!��b3��}���C�a^Y���q�p�����H�C�
 �i>���2�RRT�Q+t�K4�h�z)A!�z,���Whܸ\OKΧ"x�?w�:z��6�Z����Q`�+U���R��'��i��|W�kr�!F~�Щ���,xm�����E; 
�އ�_9���?�	���g�2bR,u�n�ؐ��H�MǄ�O"����k�ח0#�`iq�7�AcD�A[���M��Z:�_<^#���^��B ������!��I�"���5�}��6���> M�����}fr�$�a����6������ո�q�GŹ�l')���M�솆���GL\�k��x]�p�*��$�9����"�2����k#�3r��J�\����?�7dZz%��h�m��V94���L���=LC��"F+�� �}��U�PK��rk���#��ޟ�dGqKh��5E�+���94�AM7�+���'�m��F��|+mL{��M¡oe���Xr�O9��M�X�},����q�I���R�ҵB0F�F�d_��φ!�6ϭ4�X�����K��hu�����N\�Va���n����f���`9��7�������n��PԜ�is츧 �a�l$�,[4��/���ڀ�-S���w�M�eTp��rg�8ԯG�~�v���8�%PAd�|�f�z
h������7�h��y��u+x�~�J	q_{J�H���#�B��i��l�Oj�_�J�Oc:��豈���6��� t5Ń
 =���i�����Ӻ��Q�k؟a�%-�����*]Ru����՟�DpV؇z>_��	��O��_#-��f�,k��̓Yc$����,�j��yH��KF*�aG�F���oSW�ȌC���M#���� M�y��u�҂����8s�=��<�`����m?c��0lS��=�?I�����Tvh�1�?M����_�+H�%v�A�����:����tq-�����ц���'�>�<�!��{�z��4?G��ӌii��Yr��>�s�U��񋢂%.�l�����c��#��.&�33�'r2��w�<y�8����7�綐n-��"����W���<��>
��?LR�'RT4�+��.eG�:��F�j�t�B`��C�̝IU���C._bVO	���B���?+��D�������	���xZ�RfO��|)و�~
;����iD��>���,���|@�=�I�`~v�����rN{���G�/����/��8O�{.S���?
�TƷ^�h��b��𤶼n^$�Ė�LO�9�����>e��n~9������4�/Bz�lRT��Ip�:Q�R~B]98�i7�����VgO�$����u�3��}TJ6.�I��\I�B��}Ҳ�$�Pv�3�% ��|6�2ҙ��Lg��*��Q'6���3����Ph1o!�/�M/���w6�^�VD[���qD��.U����("�1?C��"��a��[q[�,�F�c����>ȚQ�!;Y�" Bl��ٝt�P�2qykV�m�ld��D��9zNI� %�r�H����(�mm�Z����AN=�z*�f3�1��̛�pW��� ��3��K/I^t#]b�oJ�^�b���t$��D>C�W�|D��C26MS��F�B3gNZG�eS�,���t�m��v��fZ g:�t���l��L��=|x
�Zf�.�i�7oBl3<Ӵz��إbF�ίO�&����c�L,�&�=]��&6�/5^�b��Ǖ�������{x1V�%L2_�e�7 ,��pZ<���t���c'B�;lGIT��X�oO����J$�5�_����=450^f�J��������Z���Oخ3LN�vƎ���X|�x `� 6o������5�:�D �}����4P=�q�xYGꕰ���+
�36�h!;�5����u�g\�4ј}��� �����9���<������u��4��,�f2� �$ѳto���6��
����*œu�=([͸�����F�@�q�PvH�0��OE���k�6a����ǵh,��� �ʗz�:��2�]L�AAR���$���f��<��8ӆ?����&�X0�FAN|>���#oqW��L�3���,wL�cw[o��{]�y?rm)cw��Y�D��?W�.0���X�Cpр�]��$(fk������Za�ۋJ�^�kp� p#�Ȼ�0����gW�uq��Z1�FK����*�6�P�'���e]�ISY��òW�ޫ�����:R��|E2���x_�z���5�v4*�2�[j�����y��9:���,��Wx�ba	�}:>i�)�(�R�ڛ*�z@���U𬭔�W��k��bL�c��P@��pQ�>њ|��A[������Jt�7���Ĝ��5X!�'`��nB��µ�:�j�W;G��]�ث/�����Z�=+X��+�K.���p��b�)1aa��pJ\k�����1;��iF�+�u��� ��ߍ����dS���Tr���n�4���%�rAd��7԰��SYTn�jn� ��[`%%)$�<��u�SG���w�vs������� o��@�C�5[��Q���J/��)����/�å���l�
�\BKEN<�caAAq�P��wm��vS�<ݵ�+��g� �h��!�~Q��*ȭ��A��d��iR^ׄU	�����m�Q�g��F�_��Ӵv��vH,zS��(1�\x���4�e� ����"�[�[���$P���� �"nS�q�f���$��������+L�ɘ�{�R�񺑀�dL� i��! �\����bF���D�=K&�L[�L��wo�▊�;K���Br��*�A��G����ُ�~�ܠ�w�^(D��22������d�ݲǄi�i"�,��3�b�r$�ng&��k{ܜ����#����u�G����2�2C���F��m,p�fH�ϡ?T�E�&�^���Dcɭ��I�A�A�G�w]Hvb��
�g�d�����Np.v2y�_�쓩���,�_q�[��Ad��cB���w�����Љ��>`�G�s*䤐��8Ɏ�vp�б.���|1-�� ����ݦ�qw1�� Q����?�m���M����\�1;>J�G�lFL�z_Ԓ���I�)d/Οr������0Gԡ���J*vU����$��OQZ�����l4�	J_���o��g��)��x͝ϸr��P��S��U`�,��,�vtQ�5 A�k�bE;ϫ��9s�4Ϸ��TDbψ���\�۴�ߴ��`r�ETh��ϲs��*n�R����H5���>��`t�8r4?�-��]����gV/��x���"��F��.��$\���0>�ɘH#L���q�̳M��GV��Q��cUg
�w�1�\L3,K�N?�Ys�ɿj���J�!f�t��~���z�tr3�n.��M����0����q����z�9��0{������j�y��JŠ�AYE��1l��/&����L3��y��v����5yw����{���Ev
�b����Ȗ�$�T�����v�8�+n���$
<)5R�Џ!���i.3�W0�Q�}����C ��'Bс;�� ��W��*��2����7��=��{Tԏ		�9��m\6/�g@��QZK ��y����i���Z�jHΑk�����L.�9�ű=�O__t���mN?	F�G�y��z���΢D�����	�YҔ����Y�+������l�t���c����+�&�t��j�V5��jù�ؼ����]�>� K��N��?�)Z���P�:�|�׼Y%�p��g��!k��(��=��|z�4�R]Үfv���!����7K��'��nBJ�~S�Zܯ7����!c ��6t a�vH��+=GSS�
L�ڲ�s��Ŷ��KΤ�A�)f��f��S,�R��Q��oƌ9�a��1ȶ�3,1V~Y{ң6]��/&�8��6?��-���P�7�����+>P����[�xF��n�
����&��ZX/cn�\Mϒ�7���xI?�G�Q����*��iV�3O���J�߲NGߙ
�(?b��Za�FS�w�3��h�6��ց�26�ͮ����Zu=?)J�r1�Y_�/�D���&��CW`c�K�d����C��9��z�̊�8726�&��{�:��+b�U�2f��$�  j>Ҹ�ʮ>��A�|�v��&Ô&�� i�̍Y�a�,J�����Yˆ���5,��H�lP,���b��Vݛr�b������bͧ2f#��ea�CT��Ы����dz⭐�>?gIeCt}�o��nV��ܗ���F�;F���xL\�yIHEȘ
�������r&��ii�l�a��|�M���5�i��W�,�2Ys^���f� #�Іj{�s�OޗT]WZ^��2v�>�Ss���I5�0�5�.���N$Et=�Z���YC��"�7���c��84NU�&�9�%�s�;��*	Et勚�2�_\��	L�M;]�hg{��_��+_=ę
>M����T��s���?�O=)y�9�d�9Z�8|�{r���Xq�R�K8�7+v�+y�l�i�9��'�g���n�x�Nv���m��5���۽�f����S?���j�!(��ck��y_ף�.��1g�g�wo�T@0��H��u�`�!ynt���U�����i�y��Sdr�kR����ep��+$_����2�cr8hM��_�9�kP�t|�Zo��ZL:�h�RYC�k��:[)�m����Eˤ�Yџ���0ؒ�SZ� xf<X�ʩ5����v���^>�T�F0W�8!���#'r�Z��U�T�
!+˥H��f���!���b%L1i@EkhZ\
+x���A9������H��j���}�PF���Dc���ՎL!X�o��)jv.It�gw�3�A8�!���җs���q ��;��~-��U�3,��b$b��cp�qS����uc�NY7�;��RKV&R�i�͍�q���=����mC�?���K��0)?��0'
��'9m���ӴXli�:F�c�rV�p�[Fc�����N��zVlRy�*�̟���*1M�σ�1�������G^�b��`V�l��������fZg(��&ϣ6'���P�I�*����i/�I�����	�ǽg��ˣ�77���;�\�;�OH�1Q~���cK��CNm	����|_R}��O
��&h���Ye����|���<�-�8����4���⵰�p�����8T�Q�d�lL����c�@�g�4�긟�~iצ�&�d�vc2js�w��?�-�Enm	����B�SƓi53��u�3b� �&D�V&�:ӆQ����|�W���J|��[����9Y�Ѷ�A��É�=7T�t��;܃3'%��f�)-�UN6�����ٙt�y��1�V(��+��(v���gI9���,I�C���vǲ0�O������<{	�K?P�KKb���TS��k�l�g�ꦠ�׿�� m���4L�fe��0���$2�����%e��SD�i>q��wk��E�?^�,|�oJ�CA�0��D�T;�i*PEx��h9�\5z@���Z+S|�����|�@��D�%��5�(�3/v��,�:��*_/���u��c}oS�bN�����#���	�)_��Z�&��3�T��F4��@�7��17ʾBu��$�#���ń�IM��1ރ;^�8?�$B��ijz�Vځ5R����yx�T�K>VD�'��%Mj���i%9�~�aA��:��;���ӇCXR%�-�y�;�K��Xl>�bR���	�U��;��&i ��\�RT��Kuo ���}�h'?⻒�Gէ×^�ЎN�� �Ԏ����5&9�����O~��\�3\k�h�w�����Q��S�����$��0Ob��:6D�9�7|�#���j��cM7�<oső�W*�$1�7������B�\�u�XY4�X M,�x|L#��Զ~tr��=��h����H�E$n"e� pc����XA,B��f��k�7�uk�v��*r$�."T��HOy�aȒ�y��i�:[�;�v�>J�&Q����`B�o�P�����/$]5�f�-����[I���J;D��N��X�g�!f+�v��&�'���r�Au_Т-�?�����;���\MƸ*�/��2\+H"�ԭ��:bG�;�!��>5�IS�'qzFY�i�Op�&���/
������A�wJtD_�t�Kq�>rH�3��Q�@5�n\K?����=�p*��4�9�ޝ��u9��y�oO�c���`�