// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:10 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JW4ohLxAhFdKn9olhEO4anyvOY3zXwqB1KAYuySF8z+/kLJFfjhsmUSH0Jny4lKF
oPTy9H7u00oWUJh4HF/EULyyDoqu8sUul//vUF7eAoZyxHO4j19H7BrUDTeYk0lR
V5F0zg2WAhKLyrpdV0BCClSOj1dK2LrSOeU2t32T9bk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 214528)
0afXTbX44QfnQ+nLzzERuTHMI3G58T3RAJN86xKQ7yM188ruAmzGvPrLjmeIvChU
bBV0rETenB/rMQjLmhk+bWb+MloXcAaGK6aw6RDP+eDvt/brv16GtnxZNCDe8TFD
R95rBDrwi7G4m5cT+AYSOnRA0KKJTDtwBpOHJ4berprRlhrXQh8FxgI6ZaYx5gJY
v/aMrvX41f7Zbp6ODbPlpGBsaOhuEANRRom/zxvbVZArkqdXpsrNIry/qvQt8rK+
B5x3ZnAxAdWDPnuvrSVFwkVSS+1GYonBACDwxJ99Du4KvdLZ5MZI5zHn03dGxzOA
731YPan5YqidxYT+rM1tfIAGbonlpPoJlLU+3XzDgrpO835gMg8sP1I085sM0Rgy
jMUJFtEaVDZLe1ltNgLeqVzYG8WkzIiLTdk+Ddz9OPkrg9perPtFS4VlP2d8w5wv
ykYSjwWPG4ZmLawjD28e7Y4/Pwlt03fjvGZAUmeCuEbQlgnClYjjKtV57i2lHK+c
K8NLVG1qZXVlUb4UylXLoIHZpLXGIUNYRAFHgpiAEo8kQ3okOyQ5NqREh3aD+pIX
7vLtfDNEb4oVE/msB1JkT+ryOu7An2AkvwKc4XgAsy4HsdsRglN0JyDGko/znc6a
3UUNbrpv/q7LjA07tboeb34dgv77PR4T+Pos8IkEa+5Bm4rPSa4PZ+K24d9h8IJz
xO/n64iEvYH/j4v2omMhmo7vGWD+z/SI+R3w6uoTiJeLMkvxfk37/bC4xXYsvE2/
/1Ly6vTqDCWhaka7PGrWIc8CjbQHfE05TVm4Nmo60VZMxHa/fqrj5Fon0ZJlexqM
CLnrOTiYngjWl+Was1QSYE+o2W4QIVKCwJxZqRrDHtjQE12iXTrh1SLxnJQ9h5FL
/T9erTluY9suoKz9gMmFeUfJW2Ddw1dEErLW+wO6ueuEp77NRBOl9fBsBYqn4pLk
6e4fOgdwu4iB58MmzqQZBK6cXLoeOrkd2rVvOBlEYK8SanHfqkwJCcOxgYNf3R8q
DkxSwDHwe96Iwsu9vm7HxrDh3cl2swEBCsP40Pa/k3zTYwhCh6gc8Ex8DKxCDMUl
HFqi1iyQDTvwwSCvGxJkwBjOyQycM6yMqsO6c3nVmxhvoLfqtMtvoZBvBCOV4RO+
YMsyzftmuGds1PETIvuFV1IsgffR7589NqdOwiZylUqVYhegS+vxl+gTIuQA9gt9
tkoocMGAAJrgfvM0Ep0y9KIKL34nLXn0tDsgKFO18R9QY5Vyc1ilnBA7bMfnk5nj
EraD5J/s5j9j2zAjrF9K6uNxfKF117vw/2IdJM+AubVReMTGQ9RPzMNIlBmbOGAs
Hlg/m2jPVUcGmeO7QrS9dcTXeY7mUwvebFvOPCa7j/5fiW+GKnZer3R5bnabphMR
Dmu4UEvxcJPNYN09zHhFaC41cCkDYYvkgcMH5ZQIFBe6LljkqXvz5cv1aLGkOqVO
zaboAFpO5+VEoSRUy8q0iipqUnhbK0KB/YPMSS6MBR5qGmK2GJWVpE3Me9sJLfqR
U3ZsVVRIDiNybzJtIS3oLQqmQrVe3UQQJhFFFfu2ZOFYQB3JZbS7fgJmGKtpVmEk
Koo1j44ZRrSXvL4O/OhtNorAdfGuxedaQ9R8MK/CMBtyaU83ajj/GFOc7sTfSsJx
xVSi7hKKxW+lCtWTqyZx23n3q+gruWCqJVPILY+UMGrnBYd3YExXjNak8+QLmUq0
mNQWfLdLcBemQ3OZclgYMcK51JTx8CKa4d14XNoOyLL7AYwvCIUVX4AlULi1A80T
tY4p94LLz/q7oxS/580myWlJ5JR68tpGII2bpk8z1v2IY4t2xJboepHHrc4clYlN
g9yj9EiTav2wq7pfgl7OzCyTRKq6N1ERaAl+K2EtPPYu3LdZDw1QTPwYzcj9eeRc
2tYo38h6U6p4C1Mylx0CF+XZMqRInfqTzqdpiAKcTQKoL7dNo8Xjq2aAcqdoUm6d
NN5xyR8qvW3f9MOipTBPTUCtj3Ij6C4d85qabPJG73Gnm0aSvb8m7gZBju5laCeA
xcntBPaSrfo2JHalHU+Q7jc/yKQuWCiFeB+GCzf3BntKrJEE9rxbX4DA6hSGv/l+
rqOUcf0O3TwLIwCAncZ/nRRofiwftbG4QO/8Npc4InOqbRSyvTHmiC0ZLamCgYq3
kVi0setxxA/dKYGsiwwiVpOI7gWmkGzmGthWbyd7+zKZ02++8EpF3LFibYN9wq4i
us2iEPwom1CwaEwU/DYpOs/9eK6kZ7jf4nyIG2LIRo2onjoDje/wbow4QXPlMnId
n9VUcRWyWjb2aS709lxE0whFlNrqrzlBxy/nHOeqWfJwwUnfwHxUT8Gbpr/hBvL5
WAmghOpj9JVQSL8n7+niPGON0Rx3OeV+xpV7HN9vMefO0f3ceskiwkpXEsnosnLi
aoW2ytx73f9LC9zWc88bZXNlF3U3nyB2GlSxmIk5fVzwPz0dD3mudTrZuDepGBFA
Wylr/RAX7cHyPFo7sOQNawGkB02lDYnvWiJnjX4TFanIYzHbX53d6ackxMlhBf9N
6BdUfndx96EKGcaws1O8JRZUD5SSPIWts+2ZNAxZMcz2DaQmryKgWCYFYWys8lsk
zAaRs/1Nv2nF1WtnV5aUJQ8IKLQeTEN4zIPNArllX0Rxa/7bE/IaVBZiKDiHgHQw
R3Dm7IR7IX2V1i4WyYd7l8tkrNyXl4g0cJEkjvDGY4+KJ3p2BYbVPQNk1n5BOkmB
HBHru0CxhglfgJ0hQPAcrvnHLVNrcyjUL+c1uoy28pZmSjhxNu/U4vMlQwP3+pW9
nHKEgsD5MnRQX2WwL9faU93hUJh0X4StvxxGVksIgtrHJE/5P5G8QxOYqeU/VEuC
mYsWzm++3HhqLPgydd553lsQ0o2Z6yJMNRJRmSXE/oNscSuZK4gVRbMfIAzQMsRh
N1EH4QY/WRzAnCUGhjHfnHX/R1mEby1Rnl5WglxvN9IkzhHKNdCsjbGSUni89StV
Ur2sbH8NJhmBJVlQB5vW5B5SdjDI/etiqSC8orGz2I/B5bR3ethZaFF0RLQRz5VN
kFZeYfa873lbXUM7Ni6STuRmXCQ+gi2JQfD2teYEBblIiuCkSGpBuQlM7rsoC1ul
Pv5nVXcqtSrWaZf7O28FGcm8Zp76Dkl83Mf7PRmfeJWhGawJxhZwRoNaE1IO9ziN
eaoxuJ7azbRSGUzU9aDrYNBYH9GYqFt9yTbSq0f+Q9muzxirHn1Vwnv03QxZcLw7
jG2AaM+wB6jd2rCASAmLxshIDORI6485AxncNVFwFrzkKsND8Ni2uaPfbP0OWMjR
wDuSuuOR5kFQdnl2EOM53fgzryajhzgVKdPJ2OAaj2M7k5WPz9T8TcxoO7LxwUXW
D9lLSgxKqbOYxR76DyZU19GsKFLTuZwWDK18Zhyais4iGJuzkG5mwh+fRiA1M4bC
kPSfYJZIMhDNIMwLe2fv0bJ37vx9oU0NWNrYPzeqETK4aqVMA01p5ozWjTPCnR+V
GJRcZbwLIFGnCx5s3hGeiVgZe1thMOSr2XQ3q5bUoQKgUDMZ3KzaMBBG5kqXuxbs
DkFUt00BOs2wLiqyAgu71H20q+3kZ8LewLqJazzrv6ZCZWmPjp3Gp5oCKS+Myrhf
2/Jp/pWvX+GwlORa1PqowDyer6RME019cudfhx4WD9m9Nd56Q/3fSh6wbVkoJdr9
FxtUNASVA4iFfN44QsTbKgcVQRB8WSG0SnDAF/DawIs4zSewYNTdtzsOr6iEQJz0
g2GBMdBUvDAkpIqTALLg+S5eQbn1p64ixwIGsj+BOCmCTSGAWWiI/Xq8YfMnmR/o
QhfuuZ2gGdBZdxOTTP4T35pZPiV/QrkTJLif0DNsjKJQtwwffn1bcWSmVKpBDxZy
Yug7SqTp/bzAqfgXrNIlP2Q/y9Bvg/Fk6cVbw82zpnNCaJSQ4bT3w9oaK5I2xOaB
fjSkBaDLVOni87qmPhevwlvKmKk8S5az7zokIkkg17pysR+AZswr1orCUBkxB3x5
LTwr0QJgJqhW0ERK2GfI/1cWtgdS1YwJ0LuXA39vROK7SEhpVWEJ456uCMxSQAWe
B8In+84NygUTzp4bz/OpXx4Uo7iT4Fv/44thN9m//OPYZaRtkc7MuoiPGNEEu5QF
DkEkhzhmt3xxQlGSFA1gjt39VPv6VXsZU9tsOLNXodCnxvlqaOdZU+LtAfZn/IQM
7MINFvHMnkULUw3Py2VGqO1X7gq4V8ZDuLtRHDFL66H9e2dGTkfBLE2fu3n/1L6L
/fO+vkZIoV2qdHppr/Ickq7hAPWQAuVOgnCnQ5Nxogh/CnloPIfhrrCyABAjYLzX
FXkW7mxkE1Iq0MMv6/wO0/KmwU2DjmvitbynDQn62LtomfiHvIxmsSMhW9Sa6xnA
270hTIN0hO8DGagQbbCIrHmHTfX827Kqd8mDI0TdXhCGOVKRnMQ6xlXJQh35G7JS
lnbPXRMljvG2NZOdUssCWYT5KKHYlpePb6RSdYm95prd+Mi2IR5LklZjY3lT2QNm
ScB7jcKJBCM7EsSi4uoLcKMRNnqMJ2PbTGlUOviLrCAuG2bnZKDe2AECab5hicx5
XGIEia7TmDR4GsHgffIOc/2i6NDFQljMBQCiUrQXdEXW4LdZbNr1fuJQ4n9ckDT7
Jh2S8z4x4KLLMoV/zLhOwLvJ6t5O3ZFHSIvj1vqKVYxTWWi9Aj7V4MExqPrsGoPB
TBJD0lOps3grlmQ2gu0aaJutSJc3cCeNwolq24PrAjfLt+VpccrFB2h8hOnXwLXU
pu2WvNo4bHJNwPXMUqlUNZ4PFjcGQa8U8nrupIkg66G/gHlYDmGfAIY4gYbDIcEG
aVVc8gryV1kYMxocscc1Zijc4jCMxf3D4j/w/H7s8TTEiaFt3Rs/2pAJPUjzn9f1
FTKJaUImLrIrm+EO3DVaYTFHSgVC0cSM/I+3a7xiq38q9uXJ4KaWRZaw3fVhWeS9
y3KwB/x6z3wpKCfz1TQVQnEp5fAqo+DxXrsQ0MV8SIY5gauOQnSVgeHHccgjLbUp
KiUGRNjTWOlwJPF8Q0qu0wZO6yDD2QZkNgQ3eRo1n46vEsqh5Ombl9S6jZ47tb2O
1NJxSCjit5NTpV3TU8iDsXt8AWm0Zm5cOsu/fyJOfasCnvzOqDwAcAnsfRS+oCzg
byIhD/AouixqXLHFf1lCiv6p/qjht5YrysFXiiXTP5Rstl3tTQI9N+KA0Xf9vpK7
gfoWY8CBxUfAm1CYtjA5FxKM7v88muq+j7vAAAg6V4HBPFivgI5JY9p9gRx/g6QN
oHiiK6yeWC9bsyzi/IkLUxBZ8ygUB6MEwwAxoXmPXEHvHiSa8nVYaMjqYacKtMTG
pIJN9nqPhkylLW8Ya1r/wwUJuIfHuYUgobMizC8vCIkbCzgh+CfC4Pkmqjd35hTp
MNOyNfiW2rMjbOSlnGPLmmU5jzMBxj/uifGPPM9PmLBWaJBIayJPULoGPb6YK8sI
aGoHnN/x8nhUTw4OXYIOd+ahs/YaisYKCqgif3qRilPMg1gufxgo0aGdEIAuWxKn
n8s0Qwz7+xnmD3+C6FE5het8jR7S/X4xRPU2wh/bSwLZI5mirFa2o3YQg2kLQb6d
RXGjwEPwRdbBPGac4dfgezNAqXHA0GBq3gfub3JV6ohS0FPwIM/xQA5nvAZfQrEU
W+roOIrMKpnR3X3Cv4Qp+2R9/qjXm7SaqnFEq5wyJMaEQoXd2j7/vY2W3/B05Lbn
Q9xe+Z7jpooH1pQWVX1AC9n4Tn/yqt4WgXWGt2Y5g20K0SNCJhQ5IbsWI1CYPQyq
96UzzZrikMlbHYo2eYz1RjV+p3OlcnL+gesdWgQDWMjhHehPCJQvOTuG42FNo1pr
pMXzrkCJ/KpeYu4kqZfl5/qkNJvK2G0FNPTsfN+wbDea9cHl4KpeUFtq9iXdnhJ8
iWPvKnMSSW2ZtI+Reqwz58UONss9B0PsU5pqwjzoeIuFthg6yDuyj2ez0YqKp6lf
zeY8JMgmoBEfs55xOIFJqUAAw/6nA8SMdNZyt7UbiE+iXAPTu61jSdywbRNsfNL1
3yryU7uIWjQuDi/DR/aibBwmCl2j+o3Cdb/LziqpvTeH7WAHFKwv+rSthjrM6G3/
2ECcyJZ5tXcoCdq25PJeuz7a3bi+9W44Jk9JMFIAH/lvzzpelQgI78JuePvp8cPM
9Q22hsb5yx1nAKbVsgdmX1QmbToto4pXH/Rw2vDzkT8uwdL9b9wuLObiWPBtDU9G
k8aMbFBqN5opt43Owi4HdHFuxbDPmcAZc4vq9NqvK+Ehd2DRT6JdknEJDcICLdo+
IvptUbgLVcDr+dMrYwb6Pae69LmbltsXYJ/kF4U9T5pglpYipNMN7+xPnxKaQoeJ
sKWHHkgyYwHLSZeyeGCU73A0flrxdClbdhMhdnMbTILR029r+4lROCUT0/ZT3PgW
fe5tO0Knhvr96pBkHgfqQFMXE2PiclTg/D44n6TefsK+g1w6yYZRGCr35JmLbr3g
taVtE1D3/yImAig9+sEStBfW/xPWQZK7LxBJ/Ypm0OI0XAgJYh4d0uresJqQnhnw
0PswAAQGwpvvGFPRuwpxQe3JcSBwssS1VuZ7h9kMjPlbhFFP5/7qOAj6eqmfSuYf
b89ln8WMtetrZEmkS8GRVS3Enk++oP9Gf0OXRThwekDOnNkTYvoAKbGkwuHReSiA
lSh5HlLpJYShayTAEwJFIZ35lLMNFvY4OYDgJImAF11N4MaLJ/auaXszC6rl2J2F
1avBR/HX8XuNUstVhIpZmplEvyIr1NFrsd+u+f7+7Aw5thw7XWBsid69wqiqKfdn
LQ2BB/OhY1PG1Uu3EZPW+rRYMztpzXPL8yi/DK6y0g+XAlRAJLzQTZhCRc5LE5ku
blAS3R115qyWvuz/Bd3yDj4E79Kwtw8ppPflof+3oPzi/pkmgaP/gp62R/cORJD2
26KOT5bbhD7p6UMf7U0nVy7p6bsQSSh4B1t7sCCax38B2bjjg2WLji4mt5AB/Reb
YEB7885Hf803KHWo31dZXo1xMnMbDOneFCqlZbXm+FtymBswvlLPz2Fi2EXy/I2y
bc23QLLSKKZ7JbJ8PZEaXDPX5RRUx2ze4dJyTid7yuKXklwCynGYay1jp6eVFb+y
DXL3/JxKOGHr1ezbaAQiUq4CcRS6F7DRwCb/15vCOa7GkWI5oEXSOFnjo9zxx/A0
feBwsDvCmv8fGd0V9xxhSiVovgLdVL4ix018hpLUhAy0QfTIBL+flhtvg2IuRkNA
VAHbNNWWDORigcXGmZT2P1EsOrN2q1vnYDT1kptQ9kqLM3eNgi1s/2w20IwYOVAF
8qGK2M7F2a4AmhNYKf+9n0/Usyc4G+5MHcReCo6RKA+nD9Kp6ABLQjpe8h9VoIpn
XRn7zjyQNuVu2xJHvXzy50MYjvFJ1argvGJqvcAc2D/ZpVJ0a7NmerrjPEtbLJys
P2R/PwcbttiLGSoXHSruxKQmq6Nlw9dCKAaxqzrEw8DeXdM7dRk8GHD//fx3wQIM
TSaeUNX6kYO/RMEWp2AZ0ChuIuqkuivEurZTCasi7qid+4VFE47WBdYWlpcx5I14
gOjAsBui6kZrDqHxEDlvurX2JG1N8A/Lmm5RBqHEdoAUMiIY/rhqPJBn7scNPC8e
4x+AQW/EZMLz9JIs1uS4ipKFNUe7YNsNF5tzKGiv8wtaY7pzsZU3F2If+PVf4I+q
MJ4nayMMNJSudBBlWUmZeiSkjWnK7SB9W0WiH0gbj90kzUMGdQ2deB+1NQnweQWf
a9sRuXWBKkETd3JKBUWX1RH0Nek4ntHM8sQbxzope6GfyQMqHPLUEmxax2sGG1AY
UzBDhvWVu9lK5howzc2cZtEQIunTzndOMc7nGrClVo9e8ngHxFkI2NZcFlMmyzAS
0nyod/+A5UEvmAUXKeWcLAf+C8NdDK3VKDyiOHioIoTBa/FNOfxW2gRHhkq0Ai2x
tAEUmQ4DD6D8AK9gN+ZTfYlrMF5gfCF14OLfynJEiLG04YQH5ga+narmP75LeMJ9
cYFGZ/FbDrwds+rOmCUCHbvXO+/8KMYq9L6rJl2oBgb6aHzkyByiKTwK1OKP+kGK
/EjHJEuGNzRH8wH6hUfzec/p1j7+3UBtt0BIq2JXj0thh4Gmyg3EJ62IfC5jkxHH
BBnmfRqh1r04jj33hTTLysWcCpDTG7mx1ldOv0SIk2+slGx06y5BalqK+xfjLhJS
+8O1cY+hjnmYLir9mmApi1fQjwbnAQ9W6J+1aa1i2oYl90pBn4L3tNtL73qvDFdg
8N0rRCJAkR84KrCztv1Ogeq73men37BbAW9sEgqxGdfJVcuIGFmJALlfALSeNYM2
8Anx7f/64V98e4L1nYhBfxSrTe79rmf2oTdOA1Wnp+r0+8Np8NZrWgNzqD/0xaT2
JSGpvuLefbQKNHPeBi7vLLO4c0xDEzOoJ1oBCzGVpauqDBycOcMm8D2k5gYuslO5
R5zLX4hsgnOhYXAEhSQQ6mm8xMBbv+U9+XJwnDhqBsgwa24XqUaVySr4kV1MsZGK
lQ+b33PgIU9Ptckn79XjLT50jimc8AUjGX/h/f/QvGN1s3Z+8sZrGKqJvWyC5Mq2
xRgqZwT/BbURJcA1UYfZN/LXF5nTOXJ3FB0UxphbKvVJaVC1faIcD1ZZLfPQIeL5
+n9iHs08/h/7fdYCa1erq5OmVLrM8634ST6fzSLXEg1dbRSUHPeWqbVI5X0QP07t
p7mZqW8jBLI7dD9KoGCChlFbgnpNSbAppb5V5uNwhJHx3r1351FR3A700ICZ4bGV
q2hOYeBWTwjbGXOhgT8q//+jHS+28I/C8I6HlCapS2qXFNKCOfJiQusyVoMsLMAA
4d2nj6ejsNGqQxYxsRB59Ps8cEwcFx5ujNHX3QBN8xarmJ6rBT6hrEJQzwWLgWsG
hO6iQ2CMrjW8fkM91JLrRFIu01Ex12oripJvrkZONIoN9H1AbOjhxzL2jIQ6N3eK
KipQ3FrDXB6by6aJfPqEqGFkL8emkflarsoa85B5gaII6a/2zZQmIIlXNfSpAbcU
+ZQRW8YDWWW3LZZX9oNJzDpVDBn9DfV9qvRfoJc1GvUTX/2V2igASfjD2n15HBv3
KF8L8Vkw+811zHnoxKWKE8Q3q9Q6Lli1fDOy0YYI9VemlbjfWFNJaf99T0kqqTip
JnH1DDWl29LADydFJrkbFa608Nd9E0cxb92UsjVzSWQrmgkunxpICBQFO97QCw1K
QG6vmrs40NepW0KEsyV4bstHJpxECSivCWNYwGS0LaM8n+tMSf3B31LeuvUcgu29
TID4cMaPGjc7z7mkH5xq/clENDu0G2XSbo5eClyLQjjuIze2s7LXW1m6uRr/YUaG
pnZvi48xWE4Wj7L7RwyPOxhDVhHEbntXyxaM2I9A2/uuHcqxVx0xnzPt2UnaTJBX
sm+Mr6Uo8RbESbWRtTxyDx0WvtbgQjxYTyOTWf9G5yqqVa4X8Ada5ytFLOJfA7NU
+hokqJ2Br1lOt8wcoiocbgP/SPiqvJn1kP307yYvE4wMy0u6PeSqfVSEhvMSWgjj
k/+iT9sv7rQjv4soEVC2sNMsVU0p1ZdSklhkJCENX3ItEUIFTJMw+l48XSy2HWcs
+2PwMAoynzER4SIwQzDHQyJ9WKT+SlzVcybDftAFt2GSYbKr9M/ii5rJ8nVpEQbx
yPnWBV//BkCUmZOYU7O3Gc9mobH2rDBWMRURWVyAylClnH9CmT2eRlAdlIe15FKC
CxZfTe/eiBFkBW42c6KN5W3LQ5TV9lutxPrlmwMl8rB4sC+ROacatzz3mPSb2FT6
2Zd9bmR027dZWAlRITg6UP4qsKxv13LQOhaTWyc581/uL8MCZaAbVUi6G66Un+UI
viuBe9cOy8CGs9heraxLVnlU4pYmIYX6qbpX4eAp0PqsUJL2D/pQKniYBDe0PSCu
D2fL9aiGOabjuFiilrqqqlUBAiBHaVTjBs5nBWyfFqAocG5LZavsmampNtKDsz1n
JbBnd+3hTB3QLoFykTqup4QJYwamoYKi3pInUs4C1Th0hBQR1V9fJQMZDJxtamQE
tKFFgLgWwFOtUdLA8ZkRBaUHwK+O4DbKpyrwMJo8TCvNTWHOMBNQQx+10qr5wlj/
p8kNrJ4qPqR1T17i7HblWNEmuRPXEol4rnR6vibnw1Yr4maYy1FYzcoYJnQPv1SO
Le3tcsvTl54I63R36lxKtflKORyAlN2x3jS/8OItz4eitTYIsmTTfAQf7djPVSst
g22E/Y+eOqtK/SkqsfGyUolE2intcMyL4N5NWnEX9epnC2V+gB7DOUTspNIjKbOQ
TCJ+DdHXiTagp221QVTkcKU+E5xTZyhFURRPy3LFa1LpwTSqxYEcHNWP5T07eCl5
KFVMtHTRtyBMBOeviKvesz8TcSfRfeU0AJ1ITOd8MX1ul5L7kZUZZHIyY4Pw9nEH
sIDz7mlKyFCAOjfo23zNOLV++mE1O0qU66FBM0H+vA0B1DtyNlbbIlLOFK39aQOu
w7OvcWMXW9A/nlgoBhj4Dt8FFtoAfifEXT/2qVk0AQPpHM/LbO4q4Irl0kRIexy2
c4M5oxFddCc1UEzNWhm0qrh9Sd/A6qccyxJZwrSOWyGfl2bT6RTDKtH4L/cXmzRi
rOBM1M2k5r4g0aYYlDAroR1bMXxbDY9T5cl1onT00G5fSYpT0TmzSB//gj/GZb8C
n2slZqxHwjVrBRUZA92yb3+Cx3E40T2hMhVygtOT0go87jJ2UcD6d16x1Y0pMUaS
lJmHpV7sLZFKIss+zopqWndbvgixSljSm4tL0aJTF0Ambj0RMyMrPwC31QRZJdaM
VTK0i29IgqZC88PchIXZKT5sWxMUKUf5FG6LZn0UTkuhOvnnlANi1jnYUH5njxUV
Ks0Zx6jsxMts9/B0QE0tNhdQ4Yrl16R4/TWu6mko1Y/g8JX3tdnTbupNcDxW7Lbb
21ZgIMWe8SsgxCYss2fN/Os06oJaUhRcqGocFAvl6hgGKBmhsu3f+X337AI0rYqP
+lEXvIVBShybkdgsRLGDkeadBYieO0fZHXHRwjIVEtnMwrW6+JeouX16x1XQQ9hF
zW+P7Xe5irH1NqPlYuXV376CQsxa+sN045LFzSDyXmJJogpsJ7uwvHCHfmeINm9s
eHlfP1np6A6CV8Vpzu3qJpTyBMzXdWm5UOYPoFbAf/nHITcUaRMMRitTfRUicFQ8
e15KtKCXdhwcLSuI+oBfhb75H/n/bQ/AbJc02ep+S6s49mCUL4CqOHOB+tTK/A+a
pkQzZRniAXeVxIByqDm/SnCo3hPNSJAUi8fLSIDq66w8SKROEkAVDMsoTWEWzr2x
MtmjPpW4oKzUIhHtDKQqMzKFO9H36+WJW23xAtjwQkd4uSUT1fO5SQPTpe3qQ+GM
/zxg+5flHh8y8AIK1YJ//lL5mXp5+My2fLiVUTJwyPTQQorgDknyYVd19g7XA/Mi
HdKLT0DDIJRchXn/5chZilLI8N/esURRs85QQRSPsZ1uQG+fqB8kV9/1yPr935RO
0Upr/XvLXOwj+w3DpUkhP7agoEX5YrRc1mAC+aTBYeqwVQZjuwV+cSMRDULr/WOv
TH2uEqohouShll4PpWritMknAMdj4+oTDxW86CdqveSWU8Sw8VprclyJ9r8Fl72A
CbTE4+cMYXgv4qq6+lftimzpwtfusnd4DC98PN9VpiJ+pcj9ke3XnS0o+TfZgm/Z
iGmeEsmiBGa3QSMnDCYW2aHy9dRmHx8m6714sOF81IT5yNzKZXgsEJXsEb8485eP
16Ohox/2EN0mg0kwpGI9bWksnDgeKmwGxYKepmIuMe//C8XiJaG2bJ/vGFfIrXT4
CODvLur+1Xk7hNVf4FNg1v7bDbtbu7pbUw4N4VQu1eZDl/Gj0zT8Iv69ydmfaN5A
k+aYFfxkHybY7NRwkfQOYYRCg7rolHZ4odS5ZQ1GMlogenEhI7V13c/0WyFwbP6C
dwyFGJ0Pj1A86BF0Hf+DsQ9U0Mqk1/dBpNb2uMGHixecBQ9knkAQnW9EFGewYo9p
H6Q957ZOAecxgSstDhXvdG68BlEuX4R0rTIk0eq3aL3qVsGxfiVylD07tlwY9l4t
kdpOqW95gfD0GkRkH5w+bjKb3MSh7m5AtZ2GRT2TPzHEg8R7o/jlHpBdM7XQMNVp
M8YmYstLxgV0vDx9cSwEhlKC6/WoSoA0QJP/tUdVvaCCU0eyhOjdXHidpUAUGny7
gEKA5sCQAik/pP9V1fUKGWjvO2XBeEtbLnaun2QexTW7g0AyNcJOJ3kSj7neH7C6
ssOskgg8KUQwtv5AzO9bIno2tShlA5jtmeZI6e8O3FXgQq+Q31VMm1i2rWEbUqQz
eLMu0QfolWUs6ASISwnBLC6bUxyETrkngsap3ARIgARQd07826FHQvb1GXNGLVt/
2jM+pjCAHsyNitUMspbndSqkjeyZfx1/8WaRgtwKJqGC6K24DdF40K8ngnGRFv3+
hKGxUKiA0lYHidQ9SEfqpYv8scsYyTbqv6Or/EpdofMWCDUl2cLADbDqmxrcasIQ
xc6eVDrxw/nMXcWjb2WsgOM+Jca0fzUHD4maxnHcVGuPnZRmRYIniNr9cg1r9OjT
hkWwt8ufFa7dUiCaSckYRuIIxSB9iiSc63we9x7Tu7ULcFHLj9N1We4UpVjwV7AO
pNQMTzTN635DWyMynKg2n467lJY6ki8CJHtFhpkSXaBUfFrmsw5DOqAYuzwCMvwM
AtBPW+a2z1k6XAU+W7Dx91n9sHpybzBomaKHVDVW31sGZGUzOUGPkqX1R+hb6/8w
+Mxs9nJreu8ENKuX12znAJgr3WGRw2bvhmOfp3gOiGxBYy7M8MaCsTIiMos99XG1
dJyVJtXm0HK2eLJzeqfAzh0fhl3ejLxd8w4+XjM7ItlQv+wNgh1NLdV3R0vFw5Qn
UUBvReCDqfmkkC19QwA6OdQSSC2r3tOBtn3+q1wAUZbktTD5F3hhh5xczU57AjyY
sQZmI9cK5/JkNTIYZH7ZILyfrMYFBbPKmxhT+FyESaRpu8iACCn1i4t5SJkaCvBC
swpx6sAjsjHWJcbmM0p5H2+lseJ5k8VNjHTIie4ftwYbJJO+832Qy9MlzRqZ3Ivb
xmEgg/EUFSaLM9V+yjnryBxltlKesUnSpmX5MUGg5S9hS2D5Jmrvk+vIpMjOJSxR
pEFVyvFtY0jYrH5H87jG4j73sZXA0ROrCtZWyjFGOEA9yOeN/modYqYnHE5Q8cfV
LX47lcrexnZh85L8iWnVkct0KK0+bN3R1IURF1hBqTCvW+sfC07Qqf7VVdGDngnr
0Y3apNXF66Rk5ynVvJSnb2iSK7hVo+N21+YlqSL1WmI8Un6NS8btTMr1znpLZnY/
YtMbWR3QPUJsjA//B48p9jHBMwQOX+cJkpS+LU8gjtxOgk9heysuD1P/Ywr7lGqb
OJofbUAU9AhYBH4X8MZ9nNe88KkxK6driyp1obvz5F8rH/58puHoP6VEddcBVyqS
VrpJuy654QcmdiIVGm6q81BlYykQFCvWEt5pLx8wuFiQ7c7zHIM4GVbXt6k2zau0
qAIS0sZKHDa4P1wpxiK4caSm/36pt34hq3eAg/Vac7rLI3bxrS4/t4zBj0mN93q5
ildWakhxyjRzfamWowohKV/j8XMAOPCn5YHQIfruVQDrNVkspdYe2A6+QZh1rpqM
r0WDI4WfvYHyRbFvM0L/nCZKkuxRN4sstWbQLHjsr3xnZQrGTntLi/kcsgfduz2x
8exypQE3IS9mAio6bDwDJh1gqB/l38P/CEbJAux3KmLBrmJnFlR8zBKssBjPT52p
sKw56je3LDP5vg3eEXVclTz3i4CV9p7n/2gqvL3CcJMKC6mlOvfb0wrIo058dPdi
Ny6/iVhlACtHxFJ+vuET1MITTlgTQ+UczJQu0RX4uxS4gg0AaZZbLb8qXnj5RxM8
sqEZWtZaZdduNmTaMhX1SlRSLJ93aCzEXCGD79fUAD6MMOQWgrIwWRTPET5MPhct
ULlCEbtPKs35DdEE7zIg62n1LjQE2a2BtMZ+mWxSXSFPPorQpWwChcm/LGNbD4wV
oQv1xLDD4/tjatR80zW0z1o/vgh2oTACpBEQW4QLES5eu1mYNQf8ftyZDvNb3QgZ
EgAQKjsk+RlwD5GIdXo+ozuvUw4KWEe6EqaFZxU4ZeKc+UZkQiWGqoZbqbjbltzT
2b/4y70dNxlUcOak2vPxxWZFtRkomzVS8xpyndQeD4Am5DQb8SUAjlXJNptPqm4w
nPwD47nuI6nm1thPC/dXGbrrUe7fTfR9a0Ba4BO4U42RR2T3rxC3bFx6hzQLwlR/
vqSn89keSN0Nl8ZgZoABBl1GGY17jp3rjziCo5d0gFaqQuvdRJ3FioQyxaLiaUsf
1GMkQOimShgolN7S7H4rtjfvhLnM5B28m/putM/v8fiQV+rqAn7uvrBAv19V8aAb
vVm7k97B+FQ/ZzK8Ebws0Olrfrl69y+qgX9RAjN2qYCnmT9QWPaVONIVHMp4PWLi
OIhc/DnkOONCywTBkISb1NKjdnV1ysmiMZO2rCeeYB4UyHz8p+H/AgfUanVdOk0s
aIXXOOYj43BNJgyUkl5/I5MvRv4PIUhslgoOvmVZvY+8e/PkkUNn7FXWd/c5cpFg
R96oTpI5DceZpkNA4uyCe1M16CQT6IddhZu8ZBk+a5yRf5IcsFhGzYDJpf0As88J
vcPhj4Vh/wudts1ILMe2JiBE542B5eMNkk0lueEfBuUUCmzHi103hnOzn6s9n4Nk
0NFQu5la1P8MOUtheH6x4agI7lJJrSqFRV8oTQzEnlM0tzWB8xYgce4CvQlwKauM
Vnr0aeBC6h6Y5dwWLOJJKOlUrklPbHwISZzLNY9BRuxKmyy9Ave0U6ECPREg1xIs
E3oBP1PumZ+R5x0nXcPOqx/PmuWhqvsbzSyZly/lDmV8noebmkOVy6+7vL0TTZd/
Ic/M3Atmhlk/z/uB1whVRPMUbdjV9U2/9oNUWIHW3nucVMyXK5yldP28fWkdwl+D
yMmk0F18lZFGW59mJvgLvS8h9ByX3k3dsbxTmdpJtFgTCfHKBhGdCjbQ9zdt+YJM
NYqx8QFIK8fXAsOmmu/kPYxWvxsNxOYKaZ47qiuJy56WVUq7O9ZE3WVGCK+BGiAT
VEoqc/h8kfJV3Hyd4FqVZrZUYjmNq1Ze6T96SnI8iM0SMWUMwl/UfJWPnRqMQjMt
CvPSY94vb4q5cNTPP55pUkTx6hjUn23LEzq6c4dJMEDLIACSNgjEu4BK92w8vubd
QiYHyapJsyIDjHDmbtCX24f3q+gyXP2jXsso8iPOkRWKEOb+y86wO2A2BHQYV/ox
vHxj5FDXAWbgOz2k9VdyOJ4pfPHbMecbAYnTHbvWniv9STMvHCjxvTffp2fHJ0t4
9gQ3F7LbyUPkOOMGIO1hRkACXMP6ZMT79D8gpVBDNHDsMcasP2lqYaV3T1q3x0uu
7FA1aNqF4yjJQx6YmRscnNrGHjur28GkvLn21K6ZjiKF3JN+MlFh+hrq21pZXUC5
6SxdkFHJTFMXQzc0r9Ps8xQHJPlBVvlQlyIdkyNGrhPpjQSd+S3i6BUcLqGoEe1i
LdymX+vWUY/Dqm0PikxDYPDisEtLeNex0bkYgoZ60gs2HtY6mlzJ0NFLdhsn+R09
eE0iJmB7CXIVP8Za8CUOz38q4LB5sUJt0iAMvGcuzMc9Dd7hPDuNv+nIpdNdbjnE
icw7AbJOjrLV0Z2fDYwPU7wii/oeEu0Xcb7MR/Q6cb1VpH3WPzOu+uJpMvlzG7AP
m0MobQIP0qLGvm454wUJwDp9mzAzt1d5S3WYJkCfsCV4nE3QhTxznujiYEODLok9
uZkKTwBgPL0gt2ysVFRkSdLyR+VzB+THHHDB2LQwP0aMWky9SEsEYyAYz+iQNd75
EihVZpMJ/pgCoUT4cpcvWTpMAVnqBSKs+fUtcy+VP4REwKcvidUOErsHO6T1LZeW
dXA2qc0ZQKnkIcS6cKd4zpim2hz3fIauOQuYN3bYhX7C10bMESWQmiYcA+Mq6Ku/
IBSPgBFdes+FAvv36C4OvR70fEWVWUTVdNxIcbEDWjK3fWg84JKtxis79M9EDxap
rVio2v2xbQdvF7ZYL67mxq8/r96EtE58Hnjex0Sv1lte8Mrnujnc3Oc+/FyeMuZy
by3PZEETdUxhtJLVtXtPaRTXeetWYNrbFCIAcyyIXoUN/NeZZQmKrzR+S/r4pvbg
XAEe8uPvOx/maB1G0y3Lfu4ENv4VJULA3oP+2I9eB8lJQcS+TRHu3Q3WT86JcgY4
yN/qeopNUdQwTOf5Z8i5hh49UXyPcOtWrQ4PlDj0buPiRagiLyXYqDHlo1U02PRT
0wOlA2yErJJM7WD8b7pbMBOuDwcI/HsMF3P7tS3PCGszGDiEaPmOzlX8DmKd2p7N
SIN9M4mdCIDxwo5Fb4O28boeGV7kahCbWQJMrhyns00mO1oWAolFL2xH/d/n6zkk
MUugCbdRcFFMG9MRWVfhK8Em4h+oA4Awtt8fsPO8n5ZAnMcmnDXtkAGmoerbIq+H
AZywAJWDn5lddEVstjMN+q3edT73udRn6Xuywm7wpJKZqP3rqmdbfO9qdJHCIcjM
qoGZXnk7rNQs8LLbKaNWHjDaF0phMgp7jJ6dFMR5Qsy/5PiV8EM+TflrOotSoTJl
h+3hEA40KH5BqnSaj4SukHWa7TETwgAJwBfQ5L9fUzveAFpu3OR+K2Avtwdx5Y2Y
STXvKwPiqiWFJJS46kci6PiXiw8+4Cxhe71xq0laznvsYniNJMZV63XW6JKg4zKo
oSeb8Tkj+GGYcxzsccH4n+kzEf7BL+XOXr0S2TFi75Eb6LcxFE86m0IS5lRuVL0k
GbFka5hpOhTNVe/hJ3Z9yOHLzvgToVHjTbDDUn2VAdXTaUbR8Xiw8jIko2SUPzhz
h3oXAQly2B4f5ohjgpkgHNjVtKdLBWtKyeaC3oR/ujbGvLPfKQN/HPBhio1gbDmt
2IJ2cIbd6RUUsNVZrMRXooIetjzbkoCWwf5exwzN0m9f2En22jLk5v+56r7lKovH
aix43vpS/Py3FQEvPXr3kb/fe8KEiDJNDzt1J1n4I0sco2mBIRawK7iBdcUOEehp
VGSNKbJ0vI7CB70gfGZ1lXms3QlLc+HkDIcb4s6TfR7oDv7Da17hE0Ha9tdI1ZIm
r6LeCBv2HO05lqVfJhHHSaLs8mKPP7647ZAostQWpJAoFK44W9HFiUkJSX8PXTEV
w8aXbcEFrkntOvdaqmSk9aeZ7s4bTPzyLAk6leihnMRaCFAd8UhjopPToBWtbRAw
gTD8sOkDAewP0i5MzQaRuAOYvMzio0tG9iqrLbmUTQQm+b2fHKRo8arJUm8wI1pu
PDayu3pY5qYTOHNM++5sDjah+XwvmfNwL0Yf+TxsZgFwY21AhQYS41W2iWkfDQO4
91zLk8OLpJDbIToffM2b4sAaN+hmnUYZpdPt9GrXpFlpPWD80Tasa/Nss54VzRdN
xpQNa2VtG0k6cKgq1l1316u/xAvoR5BVZyJyrkJPw4UmzbXUEoK9pnljWSHw1Nl/
kgNEDs7KL69VwF8TSP0qN+8/H51f0Q9G0hAriBklIrItt/vjhHlQnmOt7NvglIad
exijxFwODxm4BbxQVMUmiDZcCeMFSF0R3Gs3H6nV5nOKcQy3JqcKMEPfv8g1jDvu
wesOLS35NJ6oreQejF2Jtn1JC9M9+9TDGmegLBekLR69SUk/wCm+wKg+2nYdi5lm
dlbGYd964fJZUaGfr7PgDB1m2kgaQ0XvDeSw/kO5jHD47qFH7Zh2xFD2MA5iLdsB
TXmiZSKjjzJuAgBGCzmN7pzz7xy/DAf7VThcGdQWw8zezee9MUN/UHa8qsS1jBw1
n/BgpnTM6GPzW5P0jGFr0mrFT1RnO9wcYOcwR2NRjOHXWJZhAGaPvWjbqj4IXNVF
yXxB0inoWV3RpLgeendxlSl5JIWTVNfTTAZTUBrwa4CdbsCEPPNPyEIRL78P2SDj
MZJtrqo9fj+ZpqV5tgXpCTKE4z6lKCjH5e4XH4BxovUP/ob/bGk50+WCkDiVq+XR
N0n/ZT5NJHP9VAIzdE9By4idDjT9ISj0GtxGziQNJ6K8Ql0czhUQEI9BHuv+wyN5
U4nBqgrqBmp/FIYNuQGmvTiYwKJB8XG/XP3R8A+P0bM3QUlwSvnN+KqV/wkdxw/w
jCe+p5o0jPNSJNm/2EXnHWdxe8S/gjBDpcbvjQTfitVWZStleFAKSZdtuOZWnWwY
H6kA6avDLVI+vN/bwi89v7cUodv5w9uAJ3vRr1rMivFzCjYMBC/eG7vTw+It7uCq
h4TIwM+1eRQnWSy9j7sVy/O3h3vb0qEs72Xsor5tdWs17HrNIQaW2o06CwYMUeDb
pOQfRG2uDNq6jMxrKfsi00nRYMvCODXev4qFPOdSlrm94pjGDKcQfSpbVyo1zCnh
vB6c9aTJ/OXAGeTF3X7gesqeep4FQh3rlZJkiln5B//ukbqNjQwVXLJs95aYHbMA
yvaMcJWzBaJ70PyJtA3vISxS6Am4FvuOCLHiFOWSf+Y8nhyf0x4fvNzV2x3S9ZxZ
I2sjKZFtaTL4fvjgvZTGlEryW+u3GFR8h4tJbBHFkitV8yZ8CIfYcFYBLMtKUlb9
wVP1ll+n88t2QrfmuwDEakw93uyWQKfEZEcgxmL15vhMlT45srndgHwP6bGTMtet
9pHQgop7AIKbLwDxrZ/SpW5qAx6zdKxVb+ab4ecPFRpNV7IRxYaJO6jGRXvwl6UE
DdeN3HKG0LIbefkfW/v+zlFz+2x0V1/4Nv5k9mHqhM8+0322kQZFzwzoqF7OMVHM
f0pICNH83WA1fdfmGNfXY1ZaV2k0UkNSfsMv3pF+SgVr62Ez7dQdJuPpQ9UycRgc
I+OnoHIEzcYnT2++RcCTVFG43elmirMBEmv5c5PujiElqXb5qtiIWlzm5GNaJow2
YFRUtd+9/kWqz9VEa6evdXcERF9KuRCu4qYziM9u7AKae8FDF+rSnmFUk5mgHQU0
UpWrSvN7WH9dWecVsif3GZfuRYSHCRCOcZccZvXSwzr325oq5MO6sjK0DIEt3Ejb
5YNi+Sa6s59DxRtQp22+g4ciy3jBfGgluN7MPh2jPcImj1B6jjZUErL8iDlloaQ4
vsdiYmxhav6V/z8Blx2WCPemvOp/3dJHdyrtJexfefVVty80npiaRjIeTI0idPCq
/SitlwZB3pxsnbA2o4xof8q6cRKzaT41Axa1TldWSjBCjh7K6/FXVr4aF0zL+jvg
Pb+Qb8WEBtE1aEG+AE9JxtjrKq5UHKj0azI68nMmaH7WW2/Sc79by7AJJvQOETB1
DXBxni/n3yjIoERcoRjikoGyk+rCRdVxvrKRc0L+8HBExilBEzM4Ht6mfJ6wcuee
7aQ03diXKVv25xac0y6HdqvZppoU7VQ+OEmtKDcr5kubJH4z5PhO+1pZmGCKhiVr
n+OP4JLFpKd+/FjxWYB7zgkcZ62Qd8xSdVltW3myDH6DPhlvip62WtrogNbuM5I2
eJDSbTAJCxhiPgJTHIQXdILsH6Q+jwaCjXFSVnfs6b+Ekt16jYXqezm8gWkZeoZV
8y1ZApc+tV+mEDn/UislRl9ldnsamx2dWW3lWAPZJj53zRoBlhsWXTUEcm750Bak
/HUNJvhkx0QGYceY9ODIYx+m6zrrqlGOVYTp1wJILaGnS0sqf72lpJ8dXFu6jhui
tR0ueN1ibrcAGheic/KP9rR5OkDywnMbhp7U5ZHATUsNiiQLwqBuxKoGaJJ8noVN
yMeDwd+PwDi89hxjVIS3wDy4ZyQrhfVxjws0PmxRAgeCB/Q0OTowHU3ChQ7/+ySu
sTPQ1ZQJYzTxIPrMPV+CAu1qwuDmI7EucloQsV4uFf/svn9+QyitW1HHGhco7x4M
3OtlekQ0kHXEQbsTNeCxuL59oTTraKQc2nZti21Icl6Sh/KtoTURq+wDspIq5Btc
odWXO5MEakmDEZD+Ir2cyi1bS/daB6EU7rnBXeXL5J8koU1hhvmkxjBrqhKQ0qLj
svi28iRv7L/btv4dHGVum/DKqI8mWlRwxLSSvJd+f489/Vhzl/W6S6wR3qxBXDmc
aOipahO6wNSatN9bpkbf4/JMzdvxKlfxYsoPkc/U1RyFyJEJT3P3ApH8OQGZ32Vs
OAYwS8QUJCt9TlphjPeQPBtAgqEOowTE6lolPz1kluFCME2hv6Eop+UDUEmtB1/j
FF3FRFR/OzHnUUF4Lw4KEr6mc6w+reLednXeVYIwSj4IfSEdTEMCPxVroSRgUoLB
rs7YbPzWfXb9dAw/Owd2I1wyu3nhXEf8/8M46tNR5Qqnb7dJRXBlpKlFKA1M6a5C
lC9xDBI094Vd58eLsHYUDc4kKolmT9n/p5IGzB9pI8kmx/hs/KujXse/lleNmUCd
Yc+/9wY9ot7dDXiZKhOzUrwHE3CfP1wJBk3rlIKN83uo6hSIpAwpgF17u4S7BrJY
yp95UDrOOaVa9xrXloRBctCHxUFyUKR5Z9Fka8jhiI92fSCBgrSOyGm6O/XT6Nqo
4HdKUECfeMP5cP9HpIYW8hm0jPM3PM9eykmL7FEONId3wkhJbIiVNLapq6hf1SD9
Dq8YsM/bI1hpdj9i1+UPHVHlelrus7SUgwb6D8WtcXwYONCWh4XbbQuNo2e4mEIW
mkmInRnrt/T3hzxcu4QhYd31asZ8O9cJ1Nw4HoZqrES+vTta6bxtUcqh3cSmWfFO
ChFDIJDyNVI6D6BgwOHS1f6SS8RY1VK1n6L8jDykeA+ChWSP4xr3rvn88ZaH2ADZ
pKnUuT0azsasyWhMz01BA2IrEdbD8KiC/cp0itw5yfmw0u1qjuMpha6DLVe51i38
80Tk2CjqgOokMx7Fc2X9bLub1agp9QYrCpWi1mqAruuPyeCIatCaGXMgFHbqaEHe
UwRr5ECzA7eG10C4skxS5BDhKQjUbymt8rvZ5cj1jhnvjR3q692wiczLR7WhH3d+
TjN+GOrMBFvfzjmhfcdlJw1WkA90J/YHwT+DTNF6f4X5FH3K/nCEZ7iPKedzZoHS
MxVBINpiNvX8hj+R8JQC0t8QWM48k+3waKph/JoVqZ81e7GSlBF0hupntlmRhw9G
M50R7+1SksMgYLOU9NdOPei3LI8PAEeC6SL4NdWCA50ZoQjr/tHNUr+j5JK24E0O
RaOpfgfqzL3NGzNqoUoIeYqezNeQzTbQl74ujpnk2pl9SHUyBoZKN4FY4t1wW06q
k4qefo5IQyONzCvhzi0RIOTj2diNoHk5qeaHrBc0sWW0fnyj+tdyc/DIHPfr4ALu
IuqoX8v2zpv+bOYPwbOhmGsSQqUUHraTnQz/Ny4O572zBWZIlY85VzgI0giZAdGy
/bk1x2NqbMvYYvhL7j3YcmbsUrXhZ5OzmFYmzTKOCr4KrP0rIsJSg/IooSRzSpD2
ZOPVeDovNS+GT4pG0py1pfhaS7KqGQ1+4jDY//I0z83LvqAwrn9vFVWVgYY7Kdl0
afxAREczHndpkQWjiBh3AmuNTKF9F04oEvyaDPQyK1myT8oA6jSy/4JfU4sSCVpw
HKtsTSYPW1Gsy7nDK53XmwlHb170owCm5gBq6U2CroYkK7CaDyQmXauqfFzlaQGn
zQkDLAt/reRKLEwqZQ4MO9oPyuqXfh4nukP9wVvp/1WjqixF3kjefhsiN1VLYSpv
apoN4krz1FS1qquGOJiPLLExnvBsHjOOpQAIZ0GdC4ihOQxCFAt91ra2HkVI540k
dZPEIUPkq82ws0zEa2/KS6umlXq2uZ47iwN0NFIxpxVCvFBgILWKFQV7UqMKq5z2
1gHI8ozXh9X3kteBgSjklB5dSa9W6QVcr1G7lo4db8WBgOgAkyXSJrbm+ySHEkNj
u4rBQcOf2YyEmo7264mWn7vFFIKoBSVHioX9r4o0+rg3E60Os01Hdew4WL8EI+b8
tM1fx/zIOKvAvRTgdITZhrHDMZB/Lg44w8k/vOqqeIei8W++u8frx074nNuXP4yB
0g048kw/0YoQD7HHxfg+qnrDJVIA5+HDVIdqjJY3n2EiwxXra7yvIuzSv6EuGtOb
0lrrPU3oKs9dGpXh0M7Yby/rFuKtJFN9hpaDd18TLQ7HINmx6xtT1s6fcX3vSU6i
5ansqt0dvnOALSSAUNggrgj5FT9gfn7VfLpIVYhoX2EE/G/GnjNEt/alf83nzsDh
DzjSHuWi8S/A98LYLU8I/BWd0anoh3l8N5FJkcWJf70Lcy7hExlqvplP+sUjeGaM
lvoXGjrxYsds5Bcmibzacnw2PbZc3K17+kineCi2nK/X90o6WlPj8jum4n9Vrbmb
bo8Wdh3Y/Mn0I4m/32kceP9hlAvC9WLig8z/8UADAKIzt/OW+ykE6qEgWQyBN/tE
EaKxehJFsAwppTEEepzlnXB0tWnHZd2H5YeQwpghWJ9C7GRnGLfbp6s/+SY8XBfh
MjnfefC5wbEEJxAc8K2bqdRtVoCdPUDRJEm48FTcKDt3ttjeWNc1Qm+VW1T5+0lc
W/omq+9o9Mt3wuYp9o28/Md0LBytGkNOxnInaCvT96786+py3PiYyIOQuxkdRL4M
O63A2Zwy0VtA8V415G/NYQKm/vvNdAKHFNrsrqE0r6elCC41y2PnUP9X8QNGmefs
YoHeXxMSdGKySX5YC5JcqC4ePc9e+W+AWjPTk68qo8dfNOEtW3+CqGKd0M4Mihva
gO6araBBDT91w7MG+4tXC2Xe5bfjLZlUxx/dR+XDEDroTtM5nErcySabqqWCRLFk
E9fWwkIcBCgDaBMCJPKrQv0o6I27iOCzqMGvGb7Q6QwJuj1c/+rQAXZUW6VJEvn9
zvFlOHlcI6T2Z2E/9HEbRobHNNIA00bfUkbQCtqfpJ78A3EsDQxkQ88CjskA9Hf3
WNY9mxdlmH2wD07h5P+yntsDW1sPlHCBBvefGN3GumAPI4++TeLvAfBJqZIMi8Wb
sUiZkiOjEQYRyz9CjvnFfFnqrs/LEXSu1ASRV8VsjfmIBHAUUivFtq1U9RWBglip
Ab1XCfW4e25WaVWyD8Y0OFRvGO5A31AQlgE4VHNoWJIwaDglVqcY0MBIf87V0Hde
gqSwQbQEbus2ZWAa+/7AHy1i7DE9iH2orxhvJWJuYcndt9sW8IYKX9HRDUaGpRoJ
iMdEc+ySAFnKRmIZN8mUAXBTesLwbFaBJtr/5EXWrwIOm2T1lzxlSQMg9/DmRUSQ
CHv/DNJHozIkdhWiodIfG2G3PkdskiZ9N9rrndVqiGpqwtI5irnKk3TZi5MJ/kkf
kblv1j3yOmXsU3WK8kbkl3/kbejGSBYt0HeFGgCapJcpOaJNSCHbh7h/djgIRKuy
k/3PzYDUc00XGW2RLNvstP4UBQUA+j/B8sLvLsu+qDLg/b9TKGA5oM08S/Hy9TSn
SurRjLrqKCDDz7nrPnpyFLKSAIpBQfQ4shiXnHH+S/PFdOiZDbHt3xABzUM+Reo+
vp1Gp82cYFssOabzpE5SdNJLx/th0ZBtFrBoH7aRukppxZEddcSRNMP0GqdfUHAu
x8jqMX48xBrwDm/998J8RCSi82GMnE5DY8Xk4jLRaoZ7HoepkwyFFpvkl1s3wcMY
5tFgHIVJU7ylr7rQ8R2dgvVyYi4577SYpHvuWY2dH5JPinS247Yr+nibHkYmqT+d
u8zyIs44FWt2Kd6ZntGH4r/y6lvVBnMYEUl4ur0pO3mNWhEjX+DmctNnghsILmcy
JMlpbzF0M8RE1QHhdRfPCGD+d99oSSc8I98HWZJQAiU6sXjVYYnGk4TNRgSWgIni
mam8HCybwVQoB3BG3mN0HgvyRov2DmYQ7tU2yk0RJzLmbSZATU20pdpNj4LLkAYp
USMYGMu/rkeNivyIIqKXRHgMyCToQyqi9F5zt33YaP08uKcpn/cVkQWBrpEUgO6a
EsWlzg8xgJEvW+T6qRkxF2+6it4Wi5NmIHzoo/uwR2DWlEaSUm1XuB6yBAh3Y2Ci
ntypd4OMQtQEKaB+u4LYVe01yGh6DCGvQmmxVRjch6E1yR/Oe9lwrro2uAS0NXcp
WbgW+iiA7j6DF/Da1lJimgJOrhPpR2LPUtxsYW5tICIA4fliJbMam+yUHffCz3nJ
J1/yLc8sRu/mKKgLViHB3vhpT1giWTWdCP24vXrAQ/CmZW/ko5tS4gxy/aVKGKEj
XmjfUaV8Tq9K4ltXqYTwo3gDSduWK+62Dms1wuvLERzWeYO3eja7qLmTksmSVSiL
FcS+FgpEOJ8vKKV8hPLjK6DlVDCAQIsmmqN9LHAk93TL0NHzsP+Amyaf6QKo0Fuk
idCKEsxuczsBuIXMaWvY7VPJi7MzP5d45g81RmpkIQ45MOF1W+m5I1y3tkScv/Ei
4YclDNpxED0xfYZvMOB178D2Ilf1MiTTkpPe6fTtsZWhYZdHMihTf41vXuBTvcJc
YSMAR80q8yvsXcFcQs9VIIsp5KdUZANybJHpM7QU8HR0/yX+BVaBXGmPiQlfzxUv
4I6vf+aiU7mdUnGz/u57ZnrigDhg+ZOu5BTed2CgASmC2Qrv7hxI+H7EkzXZedmO
WbiCR8W3zynnNlenNa+9+3i6FEZylCeEihGMSeRNsUjcf6MgNtXOOjsy5deBT4RV
WzpCtntr+8+k6tyzZK1VXcymZiZXjWUw3/GvTtH9/u1sZ1DPxfCcpKPX9VBt4DUp
Oe+hYQtKfQWW9XJmQV/X7Ksz+GT84UBaVVjoBNHLUwpUThhbTGQ+VgcLiy5fPL8D
DCgMQ5w4HJtK8wJAMk8ypU+z9qtE1G+rjbt3h69coNrv5Ifo2Ch9gmvuO6xkRnjN
1uYFtNEdhgPfvPRmIeJ2a0yDnDUQwxoLLVEdFZ8BgXmyMKwjDPdF7AKFTU5RSKQa
+21P0K94L2zj5lRgOR0AfaY+mqTL5MXeVJ1Yvw4REOJDLrUnbyBYIezqf9V7Xhs+
oBAO17t5kuHwe67JXsVLw+J2PXAcU3RvKfAmWQ9+2s17NMpY26dBZ7kTCR0gpT90
giN7e276kqVaeFRDL6MSESoUNlc6Ya4rMcXp24i5hkIpuk7Kd6VIJyQplvBojTSg
85zO/8V5sQk/iJNlOFkPbPRFnXLyEPxDaro4yCwHz6nkRaIbqdQ4UQKgpOiNO/pN
olJnBVNOBRONE71tUL+OxBmdHtqErpzrXsOvesnkmhebGkdO9e+Mo28vJ5uy1oVa
en7AA/UKt2bhVLirOjtVp+lEtXJdn2bFusQkldNYWz5HDcnovSbC1+5awraEYSDS
Su9cuXH5zeq2/fj15YYOoJiZoDyLKjsU4p6DPcgku+wEWeYQQWfcOzJOZiFk2ewz
joTnoBbxw1ZTuLh7vrl/MJH7Fh81R8wgT9q/ImJ+TjXLaIQ0BgeafZgH6DNiHI0J
UDePuwLmm2SM0kUKvkQPfLMl3n057WNNlJfXfOZVR6Q3qn45MUk9+rBuJT78lAVp
nCTdVxWGEQzL8zNly8B3d3mojn4wgoOMaOh1YSOUDuSWUws+TBKSIYP4KYURLUI9
rxd03TofZdPxdye91spFEzjpTrXFGCRBMFLgECdyMlb70lDmalQKi4hBG+Np3xtO
J1gmn2NZTfEXdMcWnpEC4e8EvZfZ0fobXJoeyDQiWpv3MZkgOMa4V1Vqxd2ol3Kn
I4j7NDpUaaIM782q9mMtjH7bhZK42hwKalm0tcA/kdAW/TVRUNjhbrYK72guSfgj
xFiu+l7QWTNbWjqZDlWN7gfJH6OwowRVWZzCz89iHaPA0z8yXj9XVPiqza7JbLtZ
Ue6usfT7/kvgHYm3/wKq0+Qa7yO39Xl1H7l7xsVoGGITQ1rgaxqSADjnp0Nd7/aB
B+YXqUSRVR/2i2YQjtNAIxY2ffrYWGkvU+Ocx+AsWRc97a/rQ4xbpHW35/F+NbwC
kn2WNY6Ohx4DbOW4wiVFmqsHWmhRcRPCJ9GkL/ayIuzeMK7neAZBhd9k63cde8X1
RA+H0Y+kMWP5qZrPIBpd9vI5VBOuXiK/i2t5KKx9s8cbM0faJSEiSW4mYCOzkqkg
s1BazWGB0rjIxcODrjlUuozbuleAY318GZMIBqePD/3dEyMUTFqEEL6ru7qlgqhH
8v5vF22pJ8Nt8sAwXLMVSjVKlXVFW39Jwq4CXtAYBTNxfDSLA2ZEdw23Ak3cT1V8
Rn+0c80RJJT1TWrnxd/4nI5AeWS/9tz9A7bcKUkouw/aoyyB9tKHmAvGjsw9zCzT
aMAM6m6YKLB4U/jQLg4pMdIzAwSI4iljAN4xpZbHu3q6p3gamAQ377rB2pCLml0P
sdCCLyzZJOnmB6oCS38ovIoafcRNZo7Bqb6nusVdBwN4Cjd8GcVg64/dzRV56Bsi
A9qMAq+4PWouuvQbn4RumnmfSayEBagMp4myg2um771v3OWmsELui/t+pKHhrFUt
F0mazMtih8CVPSXVu/totaFhXn0icieQfQlLb3TCdidFLKilI33DEcVSMK499GmM
BZCZoEnlHRit2qG/m4aNY7E0gWJRMsYH7P6GhakXBgq/cEqEvoNFq6eonj+dn+aK
1iC75CHtSqg0M+AoNckn8OeJgAdvzpS2A+1GtEwfDdcPJUAfSnbBjT2ROggicto5
mkkBAfED4KFxKVqki9AsjusOqarJqeKgCE6tJrzGYVi20hPpqgt/QuyZGAUcX6X1
ERFiZxYG6gfsQmGVqWQu0Ln14zEv3gji0P9DTvPB+IxCKqrCJUKAPbNXWWmdH+MR
UsUmnLQyGU0JdJUVd1NtecyzPfusNSpQLDEhkOqcMXubMyjbiNXr1YJupC0C3yY0
UBsMd7gXCZGPzUP6vx5foJS0rNdpM5zgrew7vtijyAbo4lwiuLjdLZjkEUq5h7D8
J4BPlYwBb4bZkLE55JybUziD4vkqBGqquo1G8+GxRjNRVjYloSwknDRgiI4heFhU
GvFB822Z+YAmRx8lIvd7tG+X3osnbmkyFzEc2YopqejPvFtBB2qjSKTN6UTK6SoI
TBoIJxfUlmJjmd7TzZSBhF6A+0P8mjrvMK5qv6w6PsjAkLPGuDpt2aZwOO/M8LDO
VoVh4w6BJM/+Dxi67kPJVOHsZHLgFlTjjKxR1/2/sJiR6IecMXRtHijthuedsuK3
920TUpwjfxyFz1Wcj3M+a2qSdduBQEYe5Hx2dwyJ7h2XTBwiI1A1yl5H6/uDVaFG
AiUkCxntEds24V3WR3iZqSIBBAvMCDSbCNzNEQ8kkFkV57Tbja+eswAGWS7xvQt/
CtTkdOZojNUn8AXr/Lz4NZ7Ub8OXtDIZS3kA81f68wlnof2K1GUObMuHGZdIdGNi
IuYA5wIunMkjBLAllQWmoK3wwEWQiW8DTpphETaI32W9/D20gHsVDKIQtV4TVAU4
vtQMhpQ39jOaOeG+76ow9hPObzfAnusY5ji371ZffGbWyrIyH+MVTwtYOV7KJTpZ
R6dEDwOYyRxMi4f9iWEZRWxd2pramf+2AM3qyt1IP2DVxOdEALk0mCcQtvfWudtO
g/ZaWgDevXNzWxGg3ySPH2YhqyCcUDQqth53CXHwyjaLzGmmPaviAu/Iu+Jgq7Rb
ZQGbWPIC0rJh9OkCNs2MfqEwdxUPvhEkuKInK06/qnIHSYdvyXoceAyBYVw04OBQ
W1IZFda3ryWBuusTMOhqtQ6TJHa+iag4gvCyV7TMmZAMxxDo/0RXNlbIiLwtjuXI
bLLk6Hn8mLziER/9yjclWIKezw786ZjBBfgfiszFa6j+6XyANHsqS1lj9fLOIhsd
QAsGLqRDB/3k0xHpMgqiFgvvq+18Atqe9u9l370DlC1WDMrT2ttqlks1IDbOqJzd
XfZGfepF+dWTGOyL1U6RAf6OYILWQoMPeJehPtKDh7UkfkdxuRbwImxfJJMoSx9M
GyrHOe714tDgSSJtRTKiXTqPtn/j2ytlcxh82rPiWEOE/hDAuXd6cpKVRsYtQ7nu
fbmRJDq6AZcpJY/s23ASooBeCfWChd5hsYrXr5826xdJyI5fDKxmcGgqPCH3PTb4
TenI499G78+1vfJZZgIDNLuSMv3ayqgqsZTCVd1U/BBSjy9GiZEi6b9vJmZlkOk6
hVz7ylXNC7nukTCbH0Hg/+q1MO9VahP7dsNWCowX142Ol2+3gKzdrNR1HGAsbu/c
CeYI7DsXVgaMEIFz+wtzQ5HxpJm1HzLvPxU0mLlufNVidtoHSxMnssbNS2zemaCa
MnRwB7ShcTqi4SpPoa6JAGUXu2DIl6O/b6Thf+f/UdaB+ZmaYH2LzbvBTlA28M4G
PSbza7cXagwNOlL/JKsyKQbJ+krcZZKfaYLUIFhyE/hoc3OK6nsrupTOfWP4/w3O
Q+kjoOj2XGDvH1noFqvK0GXtpVguhtKUAA2zFYJNRzQHNgN8uhB3PZ2lH/8d0P07
wZagZTZEqiJ1ivbZneR01O+QNcJ1ovfX53qWZCJCSh0p8yhII/ZaffAKmqNIm+I5
OxnyWHL3uh3EVJh5BFZrv6REB/v05stg4QIKVO0xZs4unPW0k2/b1UaL/51J1qD/
bAXsAb+CQMB1/y0Rvch2Ff4PMuygonIZj3FBZsEA4KsYDmshMmeC70IXSVJNSRPf
WlKnswL/xZC1sz+S/JQ8TNGvZ7u0acP4fgCNpM5mRPDByf4hs2J+4EbTrwIOgVOx
6H0ydRM84LMs+abWahaapLARVdn1Cr85UMWEcwQIxtfSyeXAxtsKkLSt99MVnTCS
x5UU9m9hUCCgYLaqUYrP/7Bvmebj6IPfJ6sFf1fDZr/mvuFX2cu78wt20a6NQAQA
AGJWgK/PvipI+BbOol/5K40t/Elev3cXYYLzMvGHPEFx7C+WVv9JomNYEDG2KI3A
FjKH6NQzXEyN/3wb4mAqJMy6g7dBb6GQF7XMHi/JhThlse+pTyUztRD0VmFzlG1x
5gXXzVVAQyHQe/Q4gqJJufqMt40H5RqvxMr2cVgJNNPByyNnC6wDuuIzwOFGnTDh
DZKvF2aLO6nhCYBMPSsY6mrzpgPB+D4jQinNAz0k98t5jKJ0bcRfbWqfDTWOQyt9
+DX+FIWpLPmZNgarPHelhnPGkQ8JDJcWFefzZQsEvHeCl+dYqqmYx2LSdvDzr8RP
rxusx67VsRbt0plOkujI9r7cejvRde+YRm0oy1wDxNXREE+BSlby6DVy9bZVjG61
CDarM4Yz4oL1rsnOwNJaqJGgJGJhS/Bff6APhHxQ8P/E4nYe9+SklFIBraeMdacO
eD3n178MESuhU/SYL6mvcHTeXx6EzB7cfVFT4JSV3UVwLcTq9AeeKPCJnJ2l67on
H9e5VEMPz1CAo3W5Mg9Vw06pau8gz26eXA6ZVuREfGDNgVEgs0j5rDgNbTrvJ4nX
WDyaxSQJsJk9qbGid+zBmS+HtjQSwdWar+0bH/gzI4a8U1Waa6LXdBM8trhurjmK
53VwpUXhDJ7//ppZG0MaGNS1MNlEIPRShnob1/+uh9o/kmApm/z/fcEB3WjFrrOd
5I7QQ/2YRNJSuPJlG4aMJVL68crd+74LXDWilQ4Ht0p38AVf6YLGgBxDCEKSyeCi
LGg5n3bTVkkWT7s2ULGqvx8l46lIHv9EOPBJhELZG+XzsH064mZz1zTWi1MwdJ16
99bsByNMlf5mDHBRzwoTuXBZPRuWXNptXz1RktUxKGXHx2UnfK+I2hYZkHMF4Cfy
L1zWcVduYyVYnNfIaBS7S/GU+R6C9vbAwWj+PezBOFc9hMCqZGJ829dSpBpaCQbG
rOa8yyEA5vYD1FYw8DMoaaTssGSrxvlaeMDBbqsH2NoO8J1Di+l9Jcx9u5B5vT9n
ehsmUNBJtiN17MVzLtepSWcaCPVHtSZXFzDD9b8I/5JEEtR1dzCDmrG8+1D3kalt
gJmr6XAFg+LlOnjewXa6AsBn7/F+Y2JoH3MSCxv2Vy9ebqdFmOi9FYVKKfWCLHoq
jhHf4JEc6PN4WeCrJlPJlHJ1xh1UXGZAsyql6OzvWnzoom0KbSyXExJBWoEAnvQQ
2iZia326ZLleMzHQXMukGc2ToBF1v5xAJQIDxLXaZRURqFTvmqE1dfhE/aTCxEAG
K/MJMjvGNfuCDcownWb9ICms8tS3fhVaAxKXiegIC1O2PzsHyD8wzmA7xwwEGlTC
sqvotLsl1BtuT5vU48uFOHiFOxNE7Yeb+V94Eisba0NAlqR4JovymTaBlnHoQXY0
e29ZQys2jO3l6m7slOINN0MfwPNbhUnZFpU0muV2VSoBhtxGfcSB1zQjGyc35wnH
/vTmtxcso/TZVR7IYD4QMLDj8LNwEfDuS2rIrg02MFgtUGItfyzsWZU9bngRdhke
I8b4I0XHP5tr5HB65kcrthucH3Bm3bIj9IPaEZ/ClOXtLcBH3vueEshTQgcBJ6YP
wKxDE4WgbpFq3Cc82lwB0EhxG53g1F3XY4wnXSVBuBrLIrSs3+/qgyduPKQR/yiW
GsQJPBnuqKIt796GTjpVEngtbfWMwEl7cowKetOjfaVkFVH/uaqnIyNAgSJ26K0f
6KXXnHKKPuUSFgpHG3Le78ObLrNSx0E06tM2n4BBYhMikAnBDdnoTwemsXldzJK4
Qo3V4b4H/0cSwTVLbNHi/M0nUtcDsWJUIEoYSYF8anTvaV63IwM/qGC2Q1mMXxsu
fs3KlMvebVK0EPlt4Z57ddfYJleJfBEy+IUkeLlGDDAZZbyaYxbDn9Z/qV0FrHp/
mddwGbyIIjHrhfzNhaYPH7zn7PpWHJxyyK1WNfyz1kraMwt8MU2jwjE+BeXOtJZY
alhAO0AlbEwJ8uGdOa6DRPNKxeTQTJRfZYnFGlCmx6S8LRYRYRpNYF685qQ4Dnx5
sl6PNuwwDu72KCbf0AGjAD19GXp3RyUfIQ1Fwt7Zk1BmEWPctU/Q3P+c/n4ncGnO
HlQhVFCfcEXQER58FOM7fzsrDTfHYxElyXHhol+BQMh6EgugX+K8SoiCkR+Q7wnx
z8UU68dL/jPJsLPhxKV/PdthAmmvvc3zBAw+boR5lATjvEgDxjPosSDBnXBWeqVe
TNIGixyBWXYXYDOOn2WaFI2uXKiAO3x0uFEnrW8vvWUWmF3Ijro/XYZE4CjsvjBy
136pfzq4X9peJoueyXkHJdGXy2SGTiV7I575Oh4RPP3kpr/SWJTuXbRaMTK+K97w
4HxAu9fb2UuIupcgplzSmYMD7XRJwR78CDgtg0xtB+7XEHxPRP/OqoLHR/TEUYu0
jFZ+74iu1XqdBS+DIK1HEBh/PJBFKfm7ZJ4+RGWBkdYwfz9yRCh8kgCdkEWTLjmY
XxBjvX8jKURo2Sb6TE+sj7PZMjf0VInSEz3oAaxlnrA2l2ACnVVmYRLdYsqrFTzU
dwNjIn1tAVoJ4/oDdE9gKgNpWsdoGihNpkHnwY7MnQ1RSsNQw5/cNguX7xj1mooz
LUxq/0Nx1ShNEvbK0StsBhUv19tN1XdW3Fc+3V1i3TP/CHzgWMeKatIOXMWlQpKS
mAFCCJEpxri1y23Ohu1+Tygbo561vjQz9gy/MsrYCvMD4cn7vZJHgfiNvfT+/DGu
xuq1On6B/E9RSjICAETf7BbEZEEVR/QxKBGoU/8NduCQsTChWesw9EA3PR/2WIQt
UiFt2JfYD+YTpAcLSUCzbeLLpWultrVhRweDgb7yNIp+wo1FPJgacsWH5ElaFFRn
FhsLB8LOQoN20sf0sbHrOd/5XpIuPefFt+0ysHzgQ+WAKqbLb5vZMjrzAAIsuO1r
SbdIppzaO09kYxV/rllEhet8bWIIeinyJYHSLgtdVO9e3s2t7Sm0XUamBoMbr1HW
0o6LB/xv2ZvZSTX5+svCdeH6EXid5MLVKpBlaEVR2m5LGKBtw04izeaUOV3XXFeo
AidZKV8oYFzWCNxQAb02RCETEQaCtcYFrzweH0Ft/Sb7BH9wnSPgvYRZeMMH4IFA
6Vt/BJexLWdaFdv4XRPkVKe1YFyElcWp4V8zfNVVuisKPnqrVEv9potsnXqF5zsM
SZIesOq8VV/7XDudkOiByqDxGQ0WfJWfKQo3goboJBH9JbABLZMzUIowgrFzzJ/F
xvgCJlS0ArPpG91Ew96oFkJR8bbIqNy8+XOjizlsDmcXskK5u3+ZgTgA8FcBhcm9
SQ+Lk06nvGKWrOghzlAz1jOpIW+IE44l4ebC2uQCT9XXjsGzrqzVG20vKEqfDI0P
j/q7el8BOyDN5sgFBcxYsLLLhdiLZ4sxuIJElLr3NEarjEX+GlNaeHcXvLEnPSaq
gTwjQK8jOHWRUtEPFTvV/yZjWmO5uEJU+H1uTsz/zDysMt7Nn8t3LqQiDrd962++
izc5vU6HwGDCtfSUunwTtSuTJSfKFmnZ/WiwI2jMdU136RXFc6xp/XR82vy4Pmeh
51aUlIk1C7x3H8XaO6kbioxdRehfMQrEm3w3arFkyFzFXooTYYakTRP+o8hze91a
UTJqI0/4UwPEGNx6qoG8FMArT+nnorO48qQ52J9HlAWPD5H5eGmHMDVzmRKX2hsm
8MrUXcxLIZPJVCykkVZvHXMzM7wggNIrKBwNKt0+m+kDG1rIeidV0I2Fe6aaTN5u
MDoq8pWsn8pGF5I8OuhMpl1Esa2KfFiD2B96UMKp7Kt4M206Zbpm4VUItRbgbeYj
gxbcDGY1JHvr6uaah2K7xM0LuSZEuaCSi5lcQomnUXSxMD8W5JumAdoE8tZKByCN
WtCerFpC+OSlgTvhHH8DjLfB9oRljXeJNBaMgXM2gdv6qtf2zY+ZsfvfJAprdcA1
2RUvAviZrZK2s0j6pjgP68MYNGjf8HZf231d+RoCnQCB4muVGsIFH2i+oieIpuqI
8tfW7EEWirRsn52MEtt50b2mXgg2kCSJOLn/D6BBWEgFxfXXmAGq9PfYJ6yn3aVG
kUAcTk8SdKArmmbZ6W/qOhh3i2SX/YMvTTmERvGUkxZnwyn+1Q9BRj0y/4a4ErTY
jXcs5itTL70h9oDZixvkuRmNZwO4bHBiKlzRtkSi/4XbO7hXZ/466k6yxUwTWWQW
7bsM5zmLWsOAmv7MSyhU4tNuqqTCv3WSOWfSyDVqGq+tJcxppIp2aM2L9NyoE0Qf
SL68Dwuitmmp43VS5LIDF3uiJ8yvhM2wTjfrg2PrMErr++6H8hLEPMDn5vq+Jbzp
TgKtBwFeoN/kAkcMyQsHEQbYwiyBAOyZShqZXZk6qOhZaOrftojnPVw/9LElx8Zt
eBgR7uRTROKOFzJ2a/4iE4HdcFyeUKNzkV/7uPYwwD+Vkg97Sb6PtGrt4m2HLgKt
lLzgbBqU2lZ6iehAnuYgpJnp+GEa0Uw5emI8FBCL3tmU+hW+Hr5C0Lir4GnFxExo
OJNQlHWjGu4udTzEr4mQOTeYGdh8W3LTKaSKRbmc/A6BW0KL9Od8eIINw85gmx1/
gL8iOca4W7QJrM5cv7WNaGwXS1daXq/q//ipDqiWkLePEfO70pMaaCu53JcgyWr/
NT43UNv1IvIx4Z9UO8EXlvwZF8sbGIcO965iD/LVrcQmXXX6xyJPploVel/XM84F
JLI9rdyQ3wgmu8sjmkuliIMwwRQF1X6nNgx47+8JwXF+nq0GaiAu6g/yd9n9510O
ODfvZtWOrILpJ41OFyEa6CcX1tIMIk15FGIMF76pQWrt/gb5L/xKuoxUk8rWbNab
A1Dwkv9gdwfy1hEg0tNiUQna+YB/FpKe25PO8OlknXX8r9rTCKSRzyxNw22cyIOB
jZTPO1eIZXBBihhD8cNE4wgIcVNNL3nnYy4ObVwws+J1ubj7ubKh9BxWqbk52jMu
Zhz2xtA88BgKUUDuwJW25UUHE5iFoA/ENRlMtx6MDxBpoLaIVjk7mmSic7k3ctSr
RUncrut008LNPbwsWsNOkKVq2hZkheOaMGRcyloAxSNdLuE/jKrczcUrMgq0ibyD
5Gy57JolfWAZI9HHjKuBNzTcIhrReUkN/LF2utYEGf/r5YuqsiUIQlJp6YxH50Zz
RhhUc1udxbEBLcRST/4sEKvgP8ljysr7bX9rwwRxPRID8OLUd7FomwMZXeGwh0J9
m1bwYc4j2uesEPaEB90wkk18EbH/SbYlsQ1toXG2da2+a5L776bcki/5gFvfjol4
SRH3fCKINFR9UWz/ikeNSHnhT63ruYsk9r3KVYuBe3nJ68HOft9xL/Ej/LGHDc6b
HFItJc25g7xMvBNYdoZDFU5qMrJvjP1fM8OQARWvhNLc/o4wSWDfpYKiLQ+3aBcX
xp+1KFIu1OLY8pntfz5T4WiIU7tGP2t/AHZBIakWK2ZqU7pQsQiIzzByeCRAwwJA
Zc+Ctm1VJkeX82lwco4MUKGZNXqjhNyKL43DtCVDQ9Wdf/YWzzrYG9aPVxcvvpJJ
QBztWsTemWAzt7ynV21bXTrDd/uNPH5fwgA7ULiE4SVQysBVoByhqj5gBnD6LsQ5
6dMEK2YgINJlf7o23KLAgy9CdPFELfQ/0p5QaK85KY7hjDAqRb0s+3ywgijx4Pcz
SGuM2W+tIwMXrKIxbV3a2FLu26AoB1wBCJ6dfIqEVS4+uVmKEc+VQvOTc4UPRC23
b92G6udC4ItVETKI11amTuB1ehTtHgKLJL/ucImwk6TKAgm5+ps44eU3hjxQNAuL
2xGCP+NRRgN4nGxHvZ8uwsWkhnmQZD7rsDHLuhe6qMAzWjH9z+LywEbvlppaq9+6
TPdlaFaLq2iQVqli0UnOxblcalqxmiqP9jJFjxSJ6qczT96G2Mqps29xMVu4f8wA
9/5S8m4ALvg2+pmjA5M2jDa4t38NMWIpFYDaJGx8Ov0d0pZQuOm+gE4CsHSWFcEN
zmyUINfYmplPcaBe1SiY955jbv4ALphZ8wmPORdUrtCZLN3UvXbxTWw/QAq6HpUw
BbeF9JJ3RlHWiIKdSskXe2grlOxLfeaCxlTjqpcltlUnCmAKh+NUHqDPZi2aA58/
dP2k3iaQxhunRoM6mo4gKt2tFSDNZC2dFQRDgUIfhmTcwYSj9ZFwkM6yXCa7aq3l
H/HLKEhUB+H2hmWivhZhZ5pocSwQ9N2HHdD+YFJ3gWfZusuczuSJXQdWKwZ5T/H1
FYqliVJUHNsWB2qIEGH7sgn0Iiyalq8NbU5bFDPS7WPMOZmQ3AavjwmflYKswZtA
zEFt32wysMIHZ0FCNNw+/7Mqv7TZvipHWzc8esbAAqwLMWM5VjFLiyOZ82kf6ybb
8eHS4jHqnktCn/6+XSUHf+JD4LBp90/PhLyLvgmlNPdItjO290gzOgXZu17rr5Mo
dj6Lnx/RG6uHrTbk9RgFtQ8elTt73G8IsCntWvfpiNYzTJ1euPPROkZ86Xaqbf9K
Wv9o0uysoAUS2o/aJXNlFUYJVWYDdBZQcmoDO0U1n4ZAJa2Eo6GwyL/fa2HxFFrG
xiwi1g6t8Wkn+hvP2oS3VWP9SDv3LFQ/UlDrp/WmS3ldTqp9D/Z5hyusEspsCG9c
okoJltFDOvyglsYRTZbWRTFnwPwAYdkDiRGtg1gl2IwivLKADR0n2r5Jzl/5xJ8F
uUeGM/OaEaKk2idyBy6OYgfnpiKCBMDIZB0aO+rT3QyVCPyn5b4086YZxU/UpjNx
ZBetDW64TZ1XnbzGDvYTizpCsFI0y0jCdQVXRl9zzoRxiO+ZJItIAo4gmDKf2EFX
2wgxYP9lJ3F9pRmB9ILLKyboT+GRkduq9DBqMGhpBu4P29YGsgCEVncoDoZgkboD
Bs1rkHDsVmzbi8mn3VUH95g3rdXxDTavvGbmIv/PZ0dpj/7LhW7ZQ3izQCRvWER7
b+W8pnhUhkWw8eFSKAG0aFi58XphdylyGZIV3iF29kOhCkVjLom5Cx/t5sj+ViVN
xcYh1F7tiyCIg4Bz9ZwO1e1XegxshoH9nj4PvPBlc6fX6L9qDfleodjWfgXmw9Cp
BnVgpm98EfN/ff/cTVhkDUm1T9ge0UhD2gJi1/v5Ku0bbL63lDiaCowUm6BqM/97
C1cxuippHGCdBvUwkqpVrT4+IZPDJDz1uaGxBKw30W4BpRTmI0CJNMPruO0fUb2H
0r17xCBK1McpsOaWjTLn2oFwCpheHFonvgRpkcWqg1d3tV6fNx3Rlb4yzjGLAnoj
LaGCHe4DHtrUqCa32piH1VhwpPQ333L9zHM0YaWnQs6/XdtlIgSChKLrvV5q2zM5
oMwZZ5LY170KDmSMQPecr2Ni7S71beT8HNhd0Vz8ex2Ud/+R0TLIiEL9tAy/U2dU
InWb+ylTMshD6qNAAv0H/hAO1+Bm1kpcF5plxxaWhVYsR2RblMoHMxakEQvfN7SH
sXTE1QIMBlSraGj2TRgdzqhN9do3AwQCjlRrNgLycC4k0uMugvdbWgV1gihFzBh8
sAzHhm3cAKfIeTK9CTtjSamanHP8kEWOOO9A/AKkEjzfesiu83pn4K9ZfMIbZz2v
BirKzVcVO3aI7VT30zkFfL4K2RjagAH+ad+/KzwroaX9AidtYURbAiv2KhvdexKf
OeVWeH8pC9bE7wSxDiELWSTHyOJWxG8H0fyoflLCcIxC27A9yqsfWl2ZvlxhfxYP
pR26UpWGMixeqS8GFgs56FUuO6hXTMfqO7t6XcZDReNR/aVdYLlxN3CKWDuagREm
kn7cCAzDV2mv8IXWucIv5kaQjQQO1AUcPYogwHNk2CVWtzmiHqezyJBx2rbFmexw
l9HX3YEwBEnsgoiLtZ/6qS8/aBc7y68YadOCynzQH1z2i9aoX9mExtsgu7s9e5ZL
T7WjdqACbW/g3DVaKSSrhdw59o4tiy6ZLz8AFfGtKdEBFIblxTgixVdn4G0jVo9h
asD2cNSS2WSDWRKh4fMAd0QspIKNT3C8QTsquYtqFxjRQRJ8H/IySTcVOkGTTOF3
i/eRYaOj5SLOWmIplApcTC+UvHfNKpfrpK15suYAU+wt1otXJzwSIvfbWSUU2vq8
SKr5RP2WK0OfE0MoGcj/bfTdsBdrG2a0id/PAu7YDiw98j4/gwcsTCQ75ddC05iB
e6QtpN/1kFQEqd/Ha7BduGzaEMO6kqqZGa2bh9/50xiMGBX/yijYndnCBKWWoOVO
lDcqo6twMuWhqIs34nuN7eFZmjxcKy2wyXrepie7tA/GZIaFmDIzDUI2xqr17nAX
PKLjl/N77RaeXehTEJCYMzmyqIlGKmgYI4Msyz8QhbVn1UXonUoVAsJq4uOcIWfc
BIwCszxCRBdQwW9p0Ng2hOyD1GXquqaHmFsH+zz9CXEjoJwTh1KMVcXuApivLjRJ
+3IlqnNjx4HTLm18binRkLmtgi+1QbNvMp9mDqZz/UFfUQEIxW8Zik8SXZ6/JpJT
uOaUOJAUXpDDUaMwW1z4/qbJpFAZSsjr4XhHQEvxgcRx352/i3A4fTcwbiBR1LA8
dvzUVDaYfbu2mHysTH20bkGaan2oMiST+Z0PDocTYa0YBPmqjXLpntbmDSaSM6Ct
hFlmFDyuK2GdQYpIMm1rrLkMUKOSt+yZPeRIw6e6EIHkNiRIL10bFzTypbMGYR9Z
0prNRBsqBnJDnsxtV1FfeUQW54nMUHYo0H8zLaKZOxSYfXFr1I8eV9WAdc/epZ6R
fpCFZd5fkdyGX67uYHTXzoprcfOtrmiQxA2XxVRBD4rLyUoFwZDJbzpvWchBbhl5
CoE3Y3LRkh/LtmuXTTBlJu1FzgeoM0oWQrcfH1D/0nxSv7sMT+lMuh8aVZ2KeZYj
zvo5mLWGVHJjKMlOyVznE7mejiAu7WI55oO7cyYHXKDWfmZhIg3mzH5bF8Wx9AcK
7XWFeIhtg7cf6oZKilWd2f9pGDRTdnGEHHNSDi/kEKpdQGUHcTXiTpOiKMoQLfq5
5twLyvxL3VCoZ1jpEB19Cb66ZR4DzyqcQmj+ET58XEgOIQwAZVp+5bciRWIpBbXL
a9ii+eXJiruwcIr32s8rYuxA12H2Si44/P1M8vd8UNeafGm73i0QdcxjRZrtxl9x
Z5xyi1HB5nuMAJANhhFBCIwivQSoKHlBG1SXhfw2rkC3LmYyA8SvLj4ETroZYz/4
auDcRBOsbdnOTi7oDjRc9g2gtT2+rlGQouOQmlbANrcJJD1nphBZEDUgOwu/KKpf
LwDzbFTwWg911ABsoAOZZwrhfqGNfJvHDlv7cNm/Im2dDCJbTrPgTXjUF76IC5yR
Krk5+2qI22gTjjghe5P5hmzK8G362mC6aD0+ixT6ynlVaVDHvMoxdbJLpMmZrzRi
twN0VyFgLHPstMfhDV2jCuggVLJPzHxDvV2StW1uInPc3dO/g3rRc8XsXxWId6Fo
hCCpEJCpHwf3+PoQZMxj0OTv5WTN4DYQbKF894MfMnikGvo3CpRj3CLUYiZdSCQ6
pEKqLIMbU3i2reD2ca64EdsO3vHuculcH9I8BFTlKjZt/ptn5rQQlB4ohQ2sWZ1q
CWFWpgNoiLX3XLtcdsOJNfGMbIZafDZvy5MMYzM4eNNBmjNGeBGcO0gx4kMibXkh
p3RWvWAAPyaiQ/mUYU+ADeG4PfeYuiaJBH2bJPDvkPtpnAenu0cEzEuTdYOsUUOY
uhLejRjGoEP76pbKWfQ1d+U3QhYVI0ctikwfIm5dTRBDhBvBaZShbfGC27xZPg6A
AZ9BqqTszBGtVcRFBWIVq0gInJgEQ5DUkk6QoD5Fr4pvZGE89DQbslxa99ISLLxZ
otoS7ZpjruwM3g+PW8iE8jNgyGdC5nKahbJQMDA1a7UZPxeMQKcC52Rw9x9P0Fwt
gZcC5FSgN59ztKLQ6v2jivyowf5ItW6Lwsj6LW9EaR33mxM3E6BMSVqackAaiy9W
lwm6fM8VPzvxGM+heWfS73rjH+Mw7H3fNX3MM7CVnW8sr/TCg58Dgi2INai/U1fb
u6wV8aVTDgagNWexAXxQZ2jkkoPJ5QLtoGDO4RSjPbFExrEOklX6RPedf4GRkGgV
vOavAWKeA1sjw/aDgU0BfPiDtkriAALEOIxo3zUbVpoOTKXBS2x8S/EilX5bjpg6
1EQrXd7PQ0bx6rC/vHEU666iPBhOF3VvWW96UJOQR/O/UJ9RycBgYM96NQnN8kJb
pmghRswS3AuL6X7hVFPwkTtFp6tOT4vZBi6OhTwwHhIvCw2CsAXNUSi7whXYmwLQ
UP9TY0SKddWQZQ9pp0fqL9BAg164+uCtHIP51MPbGHFhrVLIjsXpVhllhXQ9wUe8
GuoU+msl01jg0SEgruSUI/wHRhjqse2qCliB++kPVfDGBgI0vjGfef1/E/A1N9hU
fSv5J77WFJ+RdIkrNcWm1oxnIBoOKXs+O6myXBrvPd+RitSBlZ51vnJx3V+rIFSc
gM/dCWUKcxxG5zED1eGWc3yi3+4yzR1FhnZUmRhm4nrXJxTFyz2U4TkX2KcpsYPA
/10TGMUxu30WsBSdPjMMW+L+fk6TghbpDm/DPR+Q9W1wpStdZD9d6QX5YPk0YGQq
koTymgn838g5iBOyUp3NtoUblMYZ9Q5E0SWGOYjZqPaLEuRbUuzJqacTHOYQ4IIZ
p2UA6QHc8m8Ku20atBFuC04Fbop8gd87b3GOncXnnmN7VGGneUvlklHn5ENXXJIy
uTdhzmMsCzuBxUsIAg1/+H5iHJdLL8F1lr2hixGkt/TyT4vmmiGVts/BUU/sErpD
pZZUWSo/f511+YnIIL4Su3JnDVwt1yH/oVr+Rjmnm85e5zA4FFr2Ousc2/kHjHk3
oyufauqF+lgIvSvBOoDPIl1evt+Lv1e1hJBU5utqaU1L4SQM+AtZQc/jmvJ/i8ct
qGD9u/ALiBlJph0RKbLXaZOo1HOFAZpBwUYM1yM1gj+yPW2jsc2Ko2HcK1sXFxsD
946eVoTMuC0V78KNaTRP0J4Lau3ixsFtlRAfGfFZqJnf2YyHXsFxXAd9s+3Gio5y
L6Gax4EvJtcOsBckPHU+3xru6N3fhdxvdyVTjHwIxQIvPYmyFqL1P9O6V4QMqrb3
SdxvVS6W9uHV/Kuq66dM21NZ4sJdhyLchd8x77iYCp6EZ63IG3atF5ZAw0k9U0Tn
HfBKDI2cBxtneTtTHJRZ+jB1k9DuzQIOTrPlq49Q0dtf3Zr3iU7kv/O++t7gbfcu
LZWKTMT+3c0zNL3C8I16+z7I0KyH/XCS/A8F1rnEgCnn63W+qstVjiVlk+Mu9Bui
vjUvnOZPNDGCo3em5Lfg/4vHYKm12beFNZiiIPlVDI/nPtpsxNGcVde5LxBA1oSq
raW16QhTGy+WRN1EI+AJMW/wWqUc/C9DpL038wwx3I43u4bUB2kk1mcGfR5Ka8Z1
cCDKI+uJLzAGjQt2EgiukVXL+2jW9jyuP9o8wIiZ+XhArpiLrhRutKTBTXQcxa3n
kTV/qFHYgQXblmImpxd21io0bH1zgRbKSSR45dJIfArCErLysJUbvsfS9JauY0GC
0CnXSs70idzkYGzgmjz3Qk7lo53aU5B4b4JBTL6/JvtxdvODvjrZzd8yyl/V8xiF
pfcPfuZHo2UeR1UbwotgyGGdLoCEDZm4/ILDGSXiIyVY6F2ymwI9BBzViJkfxsJM
aahFBfjsy8liMl+1y8bu9G0fN9cX/gadyo3FANQvI/z54ZVHRE6MgZOwlyISTUvB
eif7h0XOfe4/R3BQmfCiXjatF2TdF2qIPH6rkX9KlHrAkNRyFH1LluFxMOv0L7f6
qfMhWMpFkwinv6OudCV42esmHVULFvBvEEp6vcNmk+hPZFF2dbXLZvKwpsSsFseS
tcE2akyVgz9X2b6rms+5mtvIZOHxEnnLNKib3cvxoLygPXh1Etfs/w3I0pl6RwOj
tOKYe6HLXRDYqm1TNq6Rg54fTWsbgL/dXexWpjfqoj4gBhc7uQdcw3BpLYFtXapq
3IXJcRZ3iqQhxv/qoHM9wBViC7t8X95V0x4egPtts7oEGrWmB60CKJlzNuEEKYt/
gSUAzFehH5SGUE8KlVxoyZd8BdDOK6LbnN0/ijKdHsUBBzumCMWnXm6VAQsJe8/Z
3nmr1b9JcYjbswsNlu4d2fgEdYDFJLh/C4c5w/WLedNby1BVImeieev9aaR4Jrv7
hARz5a2dzJ53OQb3wnxlvNeTPsE2REXrFAwoIc6QOa89QbJvznIz8DPcCW+lmxWX
7CdESwNIUXA5us7m761xgaScKYMRtdlzcfTXXhH99wXz67S9jOVCr3QGTB4biVc5
EO+PUDumLm+WtOyy023wvCLgBzDoNs8OVDSRhTcLmow/V775E1d1XTqa7LeZT+v2
IyssL8P4/fSOTuxlgPz5Zywi15s/WhqCldi80ebNB2veUFh4702ix1X4S7Vm/Z9p
83ePpoRIEQJoSoODHLFJ69ih9MYCyxhA+LNouOUWRFU6U499VugdIhGGPnpjg+zH
7qwwAN73j+aeik5yiMbYgu36M+89YsAVbC4/Zlkd6fKJQWP6XLB5JLOuJ5MAafqo
DNycWLdTJFjm0kt4mjmXf5UqpJAtQ6hZAp0AL5oPp1C9wwAvrzG+FkHEPWZiRkeV
lPhy9wSs4VlVJ63KQlcuO7jOgaJDwb50RjaFdWqV6XWK2or+ZEujkK83iPZMPDoz
gs93fB8fSJckfe5vJ1SvI82P3V5cVfGGpLSgXNs41pfpjOG4sawH8WTb61wtpA+8
VZzqemAQAF6V2doNno8UPwaTOK8VkS2+bgLbRLYUtIEELOavSsUAZbRhAh1jvl00
buR5DvWtDH8wH6O7z0q6f+3I2S/yErNvq2TW0K0iYn/+HTMw0wDfdpMGM65EZo44
uVtW3Tn5fs5T+2EinDBKdbEsAmCreUBU5z20X53Sbu0SW5nYT4Q4TvV6PTavVOnW
V6UZgkHAalO185RHQ8QikFkbZw3NP8mnjfprGG+4+ly6cco+oLj8lf6d/40mnRRt
ksjQP16Io81aHC+Nu+UqHNFkya83Anibg0zNShnU0ufa0kQRLsY2Vz/7VzR2PO18
Rg3ycHfUcCP8f6N61dY2Q7qwN7ydrrIQwnL4sJfWa2iTCyRrdzAJrghPcrvnBwvK
8Q2iC8qRqwa33NqA0lxNcxbezu11hY0nH1s/4VrSdoBxNXPlCgn0hPLYsVNd9aP4
gh3/KkxErd9DY47YhPGHUlajI4McTLPfWMwbB4DGu/nJnxxH0aqiNs4ucx6h1lM4
iGXasdqzHFD5mJ2SkMCwyCUBMijl8noYEqOT+i10am2v8GEhrgBnPZYhoZeiejs2
1eA0IXFqn5ukHMyAB74rHD1ptnA94NjTStgLoQ30aQ5OxJm/vFmr+Si237LhXPr4
mlyKva2ItRE6mEHnhZAzOhgzEkU29ednEUs8bhol9CU6zZwAD9CQv6YX6fsTIySC
JKetfikVszvhWxRP5L9OQTyWdI/XENRsh9+S/1ecKocQqGaupoLidGuLEvRN7NPq
2Cq0/K2Y4Q/cSx2pcLE9HK6Te8Dnm/0W5YGYgY8BzdFfhOwi1FDS10oo6PyZuZvL
aWDx/U86WpaqXsvtXCBfxXzPS+3of32UNf7qVQr1kOOQExdukmo26Kurx4S7JfVU
Z6CkSROG3QBB2Gs88DhEq4LQkJGtfgu2bpuYBzL/iWCrrLPFtIKxHSq4ILMs1Cvd
DpJaVLZfnFSUdQlNbNXPwuG20HVLaY3OFclvl233HqNuPn5SLe0jlDRWPX+pw+R5
EnEERdo8a2QX5nL36ospcT27wB3KYjgnYL0CGwVBwGUskoT5hr98R92NLQutkwSl
XsW1gAq34IA2NBaBMoRhPO8P5cbQ3rOayvUZiCSEN8LydmxJsCY7FlHtZGDQtXL6
StUTYPyc8pjFMh/S9IIp3g8YMfBZuXWUzT8azi1Kl9PEx1jKUVtIDN/ifufOYAGc
RZIyUAPeZArR6fy5Rx9pRxfb1ZdbfdnfpgWtcapGbWNxbLyOlpfDIRTqHmqQp1eD
M1eUR/JkJ2em27loYOvjrBHT7oPCbJURbPwl0Fwn7DpiXXYdIMR3DxUyl85WF2d+
8i6vVKNMpFUszeQvVLwSLle5OHhgL0fMF5GtAKtRqReIJbHjIilHPRqVV1VktbyP
RNLnTSomZCKN0AMNOeCVF3djwSb88PKN4byjfDO0l5Ui6QShNE5nO/hSfR1GNGPJ
tnYWhyqdHQhJ7Bkz82bYzI8p6CrJir/IVi2yYp0TOdEEikKMAQeO2kdM4dm6wkgS
167Uf5u5aTU8h8cjXSPstdy7SrJbyKhdL9/CFjEzfUbNmFsz8RbmjiQ5a8u+Did9
0d0SAYXj8R8TNfCEPg7p2VpR+iv94HJ/ApQQx9bKLxWWdgBJtfc0Sot3X9Q72ufo
MJvXaXxHQVgdL5RexmpmuZUo5DXA4m/P5fa8aof8S4rxIPeOUSFwXCA7rUkz5Pp3
Be2BSPN4bLNvrvgkU/RTVvnujNBQks8FXtlx51wZkxvKZHOkTw2Zun0QTg+imDEe
o2vHD74SjBsxlC8AigwsJlD0i+sjl1VYl73kcu9c9XSMGWcujWCJa2cTkwBgZL+j
hqXqEmpfd6SThbow+GsyghSUBzXlERWV/75S9fEsED7U4VtkJWLdDzGNKHrDMB4H
sr/omrdq2NgS16Ol6eb1sYgrd2qk4qb61RdqiiMan9DiOOSGs0EWNniEdTYr+jdq
aPQ9Oi/4/7Js+7mmNvzDd9J1SKIg4I6LdviqOyTOwpt//uxLgiqodOW82B9l50ej
i9XcMPrDHOrZWT9MWe6a/mEbx4ThhJBaWXt2ytgVXPXjqOnnYcO5cCPAs5RBPdRo
Rmlgka55z8Myi7zMiWlsaw+lk6S9Yo5yhv8lZkNkK2OTQsqjU5LgM6eC3s+mMDhK
dJ2j8rKqX3Z5qHI3m0UiPhlYixF+Lg0pskT3EoPdcseWH/YmWgz2ATW6bsWeUUmD
xggxnmM5lUOpSapPQwg0bpFgzeAKING6XKb//GJO/3ZQLnf7376p1yY4El7CGW/s
/yMadFKOjLvZ83QDOg8dZQTI3YfqavxuBT2r6aKdMtu5z5MEp6mI0pJbyAMbPENe
jf7RYOlseE8ixvGaqCFSB86FF2qU9WqINy4gM2qn+SBCiekaT7o5oM6ZYJWU8Hy9
o0zdImvxoYzLNUDf16iQ2428lEO5tCDw7h8LyhfuGrWLgxxt+Bhnh+6TdtnT8vyt
6W445k0OsTNW1e0sWA76RFveY2XPJb00IPv8am3W4LeHnTu58WCbGkndNvW65Z87
fSkv1zw2qrBXqL1zLsJNEIVWmP9A/aVmkLsKsjQMR8A3TVCZjA5o5Wuuc00ZRv2C
EirzSTQurrj8DD8HiCEZLSk6yqgwkMBWouJJfAMUmErcGPEjVy+iFuwGk8DjXc8f
ub7K/1cNyxrRviFJf+NaD5jBwJpkZS/prEUXqlRJy0wkJMsSO0tvMu4rJCCJzNzM
orjoVerEldjwcNhB8y0GCmqY9XhENEYe3nq43QQZNmVHmQd4uaadlqWQ9EjX67fn
1x6POVtX17e/t1Rki6wvg6xG3qZ1k/URtYxb1UCqlQ9koGwKZown8s6xUP0l1lO8
p/zWhsZIYGwwoxx53Kq99WHw7dItQtkCBjjNWP9gvaWKMQOYjQR5pTylSaFZdXiw
5tS/EUmY1LfZA0++i8zSsaCZfMH3U71ivddbSU/UADzBtMv78yIyZ2kZ06BZWfD8
mpz+nDTGj5wZ0Tth4nps0+TEuW8kCUvrq/yAmJ5STqggwLK7JUqIgjEgN6mZxj0T
g0ZtWzYYHHq15muVw0ysgEf4HQAslV9Upu7/JwF8wo/nAsEvBdMNcIUdOWHv9UtU
4bNXhdKYugjcnMXw1o9sHYy+FzD120ZfHRFtybH9+f93yg/EIYrv7vxMW01Zp49e
XOdFm7dtpf5GZzlcSUJbPBbbkRoa5nE6MDxtOhXx1dvLTriPaj4WfuysE3gn2GCd
CPHeZWWt+j4+DZkA5lxsXe7NZpQe95byu9tpre0U2uCJReXeCU9WNAwmoEL39q/q
YzzSTENJPYLz+uAZJNlLl1v1QPady4atPesaqQVSXaNLkvGMTR17qiygCJJkaaXR
v0m1t/0wBQJsJ9NXF8vbiO7Sz4pQLqgwK2TI0HwPFoDgDAwPtcIO0g+tFLU6b7QM
Y3OdMgw967reJ9Kz2UZaH4FbRRLS8biOUd5oLLXB/CpAhiHYobUZbKU8pagxhZSi
0sBxH2soafiSLYC3vDsNQDDu8PUxKovm2nnwkZfIXcJvj2wWvhlpZMXdpy3Rbz9A
cUZaiy1No/8cTFB8JSYE5lkI+LwoNT83d3vfRpo7DtiiZ6wQS3cmTmuxemCArTFo
nSRm1hA7eAiBBwQbxN2wZmIkZXXSiNiMgjsP+hUXcyc9D7xXwxB2gXheFagTC16j
i8vSs+Hu2f1Huss/H945kzmKseOLWq7UytNIT9dyaPtS7YPVglifUSvyTk1x0XF5
tb60+H66qHBPxkgqK1S8keWPCKcxMd9ZqSTn3cqoxyUkSbAfRQgopTqPH6217O0z
hIF0WUXhr6Xt6pdiZRotZQGtsneNpGtZP80DqiMYbqAObuM+lJe5Sy0uVVhmGiTi
+Z5mDOuwP+RSuu/aprsCYuCDCOv98bjAa/tpKRtV9GRusp2ApkrrMW7bWWXN/yuf
iDtKOfbSL0xLb1A6cv094e8Nn2K1G2WGuzwKMGz1pNQ1Ys2fp9i2l5QLEePs4yBl
VnfaCCe5M61zbBDyi74ihXhPGVnci0yjkDyol3Rzt8yXO3ieQFNOqAsytp7pQf1q
iHPvl/UOqU1Vy91j6GvcKQWDBH9QEU9Td3lX6fEp3oEHJmzHJ9TQvpRSvXr8hoQ+
GRVn/RW5ywvhZj2c3ZoC7gU+3swfQ5FnrDEvHdmWPuO9N1jj05Cap9i1aVI7GhN8
nmnh1+F9gz2v+e2CnoL6FHebtnDbxHUdrMgVLFHKCFL3ThBPLWaHrrVBdo4fB6ll
2Nhgtraagx8M0USCEH1dZYViH0sYb1auPSlNgQpGiF+RTjsloW73vmD+CXfg6pW4
Cu8IHwX6MUZKVP+39y8uFERv9lpjwHz+b7UXJkPTXZLSwIDEKjitqYHMjQVT0ZOb
ps7Wc9vkmg+vz57HcrSye2j+YodjoyqN5LtxztiP9tdhzeuNx+3DExCJD34bIRW8
+bjoKI0+JmE+5hwjQDkBMPZpN6R/uz2n26dOK/rEN8JinZd7WJB2+OMC7vcJAiKS
V3DYwqx5B+U+sFBH4mSzn2txG9lwbw4sb/I+D1IYc/YZkc62vB6ZJoyoxoPIbmm/
YJh9OX/mPmmrO0iGvNT1KxtGP4mVR3gtpNTJkwC6oyQn9OfJHFkun5Deywjo1c8d
ecP/bKQcRGUMYCc72rwFSA/+bEatUBy0chuh8UViCC8k0Bj9vJcWySRG2ByEX5/Y
zte95j11+Navjh+knLWuhy29eZEQ6R/a8RdBPDwUm669SN9Zdw35THenk2JJq+Hv
LWwZeYyOeRPe2PqfaQuHHqE6hI1DlX7HxZVN84QYWGziOp65Li4U6AIKdqnjsipf
qke+8uG1LeiaRs6UO2WlgriXZHoWe8Z6LoHTBqCvvbSFxnyj+H3K5AEPQ8eWwXje
Nho6dhSRNpQc14Ln9Jy+7YgTdeIxK2N9j4lsbVs2Rh+xupZDxCTKCGpmxO1JVxrI
MYCbR7+FxScwU/Kx+K1JU3IMzx809V9Tcjn0Go45SBFJ+bzJwskplpQ+2xcMBT5+
XkokjzFxexMqpAEwcazIOpzCt4hnkOEQ2K30bdTUxDjIQKqncD0HxvYjvuMiTInv
J0sa8jP132vXRgnbHcYsDS05DSEpaKBhU9YKLpMcPeAzaE6wc6I2ZzG2mUsFzLtN
kfXgIa3kt0COkIwCMCJBUFqEe9tlpJq4bamarMen97gVghrC0fmmBIL/uZTsafBO
gF3AINyEZTv6u3nM5OjWZTXHRVn1jyHsOSwO7fu/zSiXIGCW+HjHxmzdNovvCw9K
f4utuqiaU3MG3HIj6zmYWjPyh4RWErNYlMRfAu+fBsxmWsC1h+GUKKh0hlPv1efl
v95f/VffpOj198vSKP8wDUG1Zx8wt7AMzYwFZ3hnEZMacL3Enq75aWq/tXzITMUM
Bh9Prj2UUBlhAwpA1ttwFf9q8QM9uUjMAyNeObdruMh+NrXuVYbQzNPemYa0TGKo
A6bUGRMmMeZWYFHVoX3Q3lZx9TEOLFPo4ORSLGNhs3Sc4OKDE0s0QgfRPH3mCsY0
SRBcoWSIc9Jv0BpXxddh7PRIh5hGxFTbqtB+OHXURXUt8A3SHGS7moXEI5absYlT
sDI2WfKsdJzMnlCkCXRvCJfgk1T/krIbbz/C+kI2WNIW7dl0RmuSTyBsnd3ZJBz8
Do5Hdn6ei6L5D3y690Bue+QKSotR2d4edpu9Y1uD0ylTlF4YT6aOarlxVq6d86qc
qMMF2oSiLtLJsyHsgRqqSB30BXeO9inB2wOG/gkWu7eUoJFdP51z/TvgMf5psJiu
ELbzqWuG3BCbl5kjjOCYmSPLkeLe7t9/qi2S6OQNOHrKItvGbl1Nul3DhYaVZ3S8
l507fHHqtz/9P0qzknvZGq4XWfRBg+QB/Cbd6hIjDhmrmH/tanpw1WnZKKCETtQC
3Raqu7mZlGWcUt6HG7rybgz2D0wFULA3KpCwEvhZVDIYC9/a3wRWvQSXX3jIfTUe
p3RRX3FgLknUlGORrrW3HBSEx4cEqvPMFoIeTPCTShYkykEKJJ8EZcLjlnTCWXbv
54wETM0AOAsdmm73lDyQq/l7qROO3RAfcFOt5VA6DFMtuM7CFSKmlM+XrKq0vVxW
ZwiKMVJOe/7K/VnHuiAfljChCU96xvJNDj6xW9fkDsg6ZMS+Rs+XDZxU1ukp/CtV
47QnnOQeFNwu7XoqmyAmrKd+S5H8efafAtpHjpkW5L7j8BzSzx4GMU9gRhjNLcu8
S8HzIQz77++hJNqemb/i6Y4XhCyo9h6q0R9hN/PA8QmgnLn++/uCqch1pqMKNYWm
v3aZTUUCyIbZD4I2RTxVutbm6ykeExf8yRASFA1gB3aSvlUs26xhZVcGpzY9qa7D
3wrevU0pswcX5leY3NEe0fXoEBZbQLB7lVhVyng4+aMTc3Lm3/hfi74J0YGHHKTr
S8cbaMX3KP/2uGRDD0AUwfE2IWvvolTUBv7yMkmiz5KbYqdEsKxeoxkuNm8ll/8C
dbJkJI/7u+J/yZLOhXt824BCr36zNq4C7Ty+p1gRg+IdwWtqVhR1bHH1o0m89D6T
ea+aIrAO8DnhrwmPIE7IKCehpkWGQL7tsCiIRIF1nkmJ0v/sR29CY+XlKGEykZ21
QAUGPh3HdyCLbjoVMjDcBLoPLdfQYtumoYTaLtosIKH5m+fuEKHz2hcpk6ZC2Scw
6zALEbc4kJHRgXdA8/DhrxdssjEivf5pdMvwjDRS73WkBroGO1sn7cdmuGk3G8Ga
9ni9xdaRexOS5aPzAwnAwykqAZvDucZ4FDwAVK7FWRkawoVrodc/UhGaLWYhUDZA
VwouXWYRgq/C7ImG1qJvIEqzkf48PDOGWFP9yBH89r5zmtn8qeeVsJ5ahnBApveb
Hk3xmGkgO24X5FnDstPXQv1IOAa+TsFyT98diJg0nczLlWZZ5/4K2ekATFO28KJG
s8s+eSNZMRb6+SmvHc7M0k+ehd/3grIaMsz9ZIPK7XU6SlS0BqvUQGix7WmzvjR9
cqJZYMVe3ctSr+NkEJVkHmTbNR2peR0L0lV0OIiIUCS8cZEmQyVruUcQM7JA/XfA
+nH5UVLBhe9byjcVA1b2AicBnjWAxKPLjhD5YEUEXvMAkTlOFwRzscz92rtfx8VK
cVPHu5kcoOE2yQ7uXAAballWZ63S9JNcdP+jhR66vMcf2r0zri1IgOd+DQrmfF8Y
hkfb5xbGWrAEu2juFPjc2OZyv4PX4MMisrHY6X3OG/jWQQiH6igBKQza1G8pvRd6
jw9NV8izearua/xqE9Sq6pGYTEMuCoJwwxhX9TFwdq/pXa9EvGl2fQvfXs7uZBkj
lUE+Ivcr0EPGvjsbNnzZmxT79Cg86RRY84457znSi90RQEKYxQ4qOF5quC6S5pFJ
dxZIXkCdkAPU/VdV1ux/BnUXxBO0sfxf0zEPk0d9S7Oz7leNZGfMvenqZUI62kI8
gIwZoA8mOWSX1FBsa8vFoHufvrjmNtvBsDKhvcgkEjpZvM5Mc11rol4qWQ3tN0Ko
ViW82QKtRPZf31MesYK68+nlTuCMYTKUHSatx3jjtKsdEZh5LZw5GorMFPu0BTlt
oPD/UB7FBzB24BQUP+EVT7lPhPm5a7GC6VhkJuzVENbpyORAq2plIVRzH2GCdzYW
g68SnrPcvplaP/6T0RSqHJLuXCqF4qw4/gXf57FW/dAVIqKewF7NYzhzI52bnUfM
YuxAX/M3Fk5Q//FDPtdu305N0Bd7lPQMrCXLlCa8ow072OSyTYyrGFN44aNkvacU
ktDwomitzsSLNei/tY/fo3oNamlEFwqMokPyYVLbgKkFRoMOTrkanhT5PDZCC5ag
HpJXfusVvys+VjhMVQZ+zI4qFiNCHp2yE8kGlh9oW605X/PIEctWd0eRSzPuGs7n
mZr4UAZv8IBGjPjKEuYT8tvJbbTsOv7HTEoktvMSGGDY7xZgfJEh5ua1+JTOLKX/
P9at9CFfQ7jaYhsctsyU/V+MlSDn1nbe5KhKxkdMsbTTj589O3bBT79LpUs+O5vW
fOUfqlc4dq0i6FQF9qqIue0g6+6DbBZyOhOSH8851bGrKitod1clTlgGepgB9x4g
JyuJki8i9t0+0rhuFardr9dmYZMerdGyubRpSDl2EhsuPQgUjy6JvvbgzXrMdPlQ
ANOKcv3F0kILpS24JTdkZJ2fFh9ANtkzxVFDCjXnmzNoQWh+KK19MyBOlvqNC4Pc
R+9k04eEye1+fM2c+vC6quFY0oQVgxWDit0M1jgiWHqvpi5mvZMh/c/ikVMZaavi
jwaDdB4dmb5nsbtKBWEUBCh7Eyjin9wRJjV9R5zpw1SCaUM2Js7KFn2zOkH71kcn
lwr4DpMkrTqbM2Q3sNrL6kOO+7jq0gtkvdIMj71XKNC7B6G8+D1AZjtPtvLk/7P4
qwHUcnBHjF2kdBwLLxSNprcabNIC5EbVqq4ePb4z3He5i7ww78TQ+hWj4dM7NC/i
RIBCozRnMFHECTbTiT4HlQM++ifJjjwHqH1AVoK81tcewx6TSpwP2GsilWjaJob+
C745LUqBAYFLDG5Y6SXNxDiuUXQqqGF/xAl7CShx8vc+LS99bpXrclF7bdzTWcAD
AxP6dDqT968rY2Y6TDJy0TPy1UJ9uy4TYoazQmhj5TcPgacBR8HX4j57I1rHZuw1
g9dcDgSVpjgfH9nKsu/wCk25uojb3rdhVLvyM2hPPolFC3Zo1mCTYY/0LcHevTk1
FUDQ/jsRxr/UZHNaeOq0SA/jvfRXSSADpiqA9Y1lrauTfOCOqGBVM/P7haIGSfuS
vxylfFHvkFDZBNbIWOP8GCcLBxqwpueZOlXbBaipIh7x4GCBE0ggQthxIYG0p2V3
YAHF/JhjEsMlsLtwqXWMMeDTz6G4DTTFbVcv9yq+/WpTvcT0QhIlmT3ml/Vs8rCs
T7HkMVOVQ/7jgBtJkxMbmdAYJIrUe1PUhWqV8f7fIBd0+mgSFUTD1WuL/kn/C6yn
lJv/Bimc/o17jSt5JamNqnBTg2rQbzEtd8jhKEjNRt/4ipo1sitbIZ5HO7HU4Zbl
m8CO5rxl3HJwHiNwL73fVdt5/dEvbS7CB0D3Ji2sTjc6BCbUj7hJqT2Nkn3NC2RJ
c/anQUW9pTWu0z+2bu199RAF/vKlSJCJuPWTmzBYueuk+l3b++DssrMnzny8XQn/
y8VJhRyYGcOLtIR5T2A0Sjc9Q+SuA9XpstBaRb9t//sw1eJKYeXZfugUIl++G4d1
Z/dbYh1emy8WLBvcBzHVAx7AGZ1f/MRsR5Zlzi2XKwBL+0sBxpDe4zIJcdtJV9WK
VwsTXuYZNo4wH5CtzG6HTHbD2AMRDDrn1UGJ2oc5kO7jBiJT+vK9mpu8WRDLnnGj
MLMMt171e8j7LRyndRBrIccFBa5jplYlbyivPATP0TMQuyY69BiRhuTaMTdC6kvC
XttK6s6iFFR7fOPFymmcLXTQmhkju7QrhiFwKvgR2Z4/f4LgzgO8qLX1avKpVgxx
OlnrkqLfb3yDBPOzC04Mm7G6BtpOrVCkuQ7ZDGcujm/NPrGu/IxyfPQ1MMwApuTv
3ycQ6D5U3ZTOnmcseT09Ce24ANvV+VbY4ZvjUynyYyESd0J5VT23EzgfNY72URzI
qEL2Sxo70gcMbBYX3tc7ZqcOaPis/Oi2gcigZzOn3lcjuxHVLfUIpC2ZPeYglq95
D6nFNvEmdWJzEWFnbrNnbOvzo4HGp6M2UaFij3dKM+vweKzxOpfG1c3cgo2EgWdi
zfQo5LhLLR4vI+DuvpqISxaxGPCLVhGKXyjYD9jFvDlClB30vrBB5s57AkEAVVFJ
6yPt63tRggxsB1JYVCBjBUNp5Em96k4Te2xyPdh31RHCFD8RDaRSC6vvyoto3ZaL
HpFDGmLFs3TZ3ivloVdPmnKfQC9wa9xhjLtywJQDcVJax+fs2zYgyNtNVcmdGPLa
+y9o+i4viHybWn4bzzimd8pdFNPzgMsQjZkGrVs+ycRaCRN+DZyhT/ccDt7w9eKJ
JYobN5qu/MOffOVzTIvgVcSwe/IdtSf3lCX6mIzB38jXo4g+A2JQsr90biiaJyn3
UJU5CUJwI31vxH995kPKOCPh+PaFbDYYweAua9cakaK5x9Q/cu5nfBc5iptK9oG7
MHMHmzhx0G2s95S8UMTXR/hxp6VeDXfYmP01SkvvxnJo4QJZA8OdH1YTu885j55m
9GKMzKOtm5//eXsAZZlGtDS8x72pG9288+pQv/4lU8Wx/sZu9Spu+DlIBg8KKVDq
F3TMh83KiC+zZh+ngy1OLzm/xEIkJ6YpgTTMGUOIXCNZuFQW9cnKXVd8MD/uIV0a
n6M+fee/LomLyNw9o6cnetOpqvSYIM/7lGrYVXAdKEvcouRPtmDiUddbG3xs9PSg
6T3MfC2rVDaIz3TuzdL5dYaHm+7iTb7vQqMBXuV30LehL8TuuZ9I6rTJDOtR2dPN
ynse0yOzloL0NNYx5qVBgMCollM6wqqunn252G0ORS4Mi/nwI1Now8HzhnlBqHj0
hlYCcjvZ1fq3dgKppuBdLBZ6R6yUaqeYsvmvyt1HGAiZxaZ+TzgsRuG2UrkBAaEh
InjSgt8WUrbEgOVyc2Gq+wJdVh2jKKAIkHUhoW+ep82JeALncf7yZUk68vK9DBck
xl16hW0Xw2cyK37HWD11jdoFcr2ItI9CKobs3efmDTxDiXFRuIcPARaWyqqMHYjf
rH4qSnMtV2t3WWQ+QLwtYVHFfdgT5PxEgrjGka86YuqIzWeiuuBekVXGRYPPras0
37Qc8KMtUDmsL1D1Jp5LaNyexuZ/iCT7G1gfed8UCLCA1GHlLkMWKLINi11hZEET
6+Mt/OcDY/1zzuzjHdJrJZTet59zT1k6m7PwJbkHH1i1nuC+q5B1OW0WN23ZcDeX
tdR5z14qa0VKFMkcyn4LoiEpjZeFZwj2VD5RpHqnMH0sZlFrxMbM76DtsbkjtdZp
ii57ndBsWxe8ieQHby6GGvgBOERFus7ApuK0jpL5X43JrQGihMK5dK413uzybbcR
BY5xRyA72d0NhKN9tf6LZ66F84QNdWqMBhZdA4le3tgMXybK7IAlJQr+LO0rNpFH
ZtKPDrFHXHxK+OEVloMjgZAWjiTjpYWl9Qzr9HIAdowGWYpGlZhpZxgva+EeLZHF
0m6nLmP8htVXBkISn3jJHJtLZxaFBYiWpily9ApaG9gGdNxsHWCa4FCJdrG3s8nL
7Plrnb+3x4+9zRxxkUd04LQyoSIPXU7Po5MHuMKHvrDI1OLgh+v3K38oG2951QVP
Z4G4TfUUUbtP35ZF+DsYc4gDMCbRQQ2urXtfINXEUq8Fi1w5GzB942O4T2K5+6PW
9hwzoLZDiR3fIGaXXVx4o7XnbR+1FKaQHNmr1o7JjV1fKVWRWI5nFWVcWHEH6H5d
IqCvvc1GGmVnqgZuCto2wH4SnqIivQAXjWOG5RuM+TsyYzIju4ozY4Ikopbh3Rzg
rtitgvFwjPOEt4vG3F+Ig6C7dhzVEuA7yw7AYHnzKU2JkkanaoxNqKJh3Q6N8x4K
yqnfQr/TTfpRfmDA5NhXfkBhNxC2mhYWlmRsfwVM9INTw2J++xDihUYE/BoOXBQK
CBH0HxuoUU0N+ws256E+p5zI8hyt4t/F1yqnLQbPc8t45cVPpzOQTq0TO9JzzcrE
s4zJjeBbuuaML0cZLZpZDnGxQqElXtGAmxt2ZJDYMOVws6IA9SGCvroj5v/nHTWD
jCz0AJdkb8aL9p2aqYUsYgOvremVNHNq0z4rPB5MnyYF/HELnr/NuUEBY25pfP3u
NSgC/ZIaxdKs0B2lwOoHhoheyf4yK9Ik/NODu7Ac5OQRTDT0zD7XOIjxcAsxdh1y
FeqHEjpaui1uqAZATj5Djre6tg4WR+JzTGbBBJglIYG1xmMszzwdV2BxJK9EWNTs
nqlZlJqW0nOXHc+mkX5wmqSXjTijnOPTUb2ifJ6xLIX4PezD6xdzAwi1Jcxox5MG
upTAd9zhGol0T+hArYwZhhu6ZQUgCb9Kskj9E1dwYt+DpILMJprz4eZNtZD3QkdR
Z0S9JrlvFqAx5Ofg+35fNsjDrsbMqFNRfZpX/+O2K5Ce8ErRlBePPWrn6h3WiMJC
OurbVdv4MW15JzK4JfWm7FMltagqLJMS6ZbgOJUdr9zTCP5af3T4A4gxX4lOe5AT
VDIK2W5XL1vRESTGKvTl1FWQcr1hMA2Li8vzfj49aqv9emubaKpJ5Iva1SL9IGUU
tpYw4nCjvmQjQf8ux6OV/sXGQvZltIX3DCXkvaAA9e85XrkoXkWK1mQwfegJhf1b
xbPOv8LyElDCjUalomo1iRQBxW6yK1Hl47brNejACrszt+qWdyPYnPrsPzjzUx33
5v5yfdfsssokZbKf7+lEXxkaulOXDeFHaGYNgQbzMksZqLWCy38DpS3TPPyda1QR
0bSPlW92Ot9Nd09X/fGfJIakPqoWv641a0l+vS3hUYobQk/Friy9CaZwepANJeX2
qmojJFVePgKqMyAZE8a7B6PZbyLpaZ6ukcozwJmn37U05IZhWmucNVqjjDpTwwPV
O5MGrGvMUQhfwbBk+kcgXsI65RTW5mZ5YYlWXcO04xpYZjp2uAnUn6RSv/AUGxPx
Ui8/9ToH2/kajy2NzVwyRY+cENJ4VcGfiVwq0bZnpN33T5lcVxyMXuKhP59xgPr9
2/gOp8QFEKlm8gjk0IiUk+cGUDcBSiFB8PR7yDm7fcoojFGmkpg3Frne/r/1YujP
F8GchTkKHyZRbA5b0bVv4lfbyVOfpG0kqwI5q/Pb1oVQvYUIwmL7CGsxcSykS+l2
f3t0HLh51Y6U57b+zjJNd1vSHqjx0cbDv79C8W61bOO3vE+Ib3/GZbs0E1fwB5Mk
zpPndynkawjVjP36RdGKz985qYSCj7B01Mtb2cQVtRxlArmz7WmjnpnNoOtqmtXL
uH26AaA5mBgrI3yv6ZkPxF02IwnKZhmyYur3uRioJjgI32FIg9qVfROTUda7bd2w
wNc/wPfNUbF2nRTa1/Qrgq/GDW16Naj9Rq0UoGXZnkHH8t3Woc3yrdtvXFauXpRX
rpXiOHcE/TYUNjlDcU89Hg6FhjIT0GyVJ8sZ5dmtpZRY2yiW5o1WzyXSNXxeZW2r
Yk7/FqsIwbHxuPFlxowI/79CYPh/nOsBgp6FyGJkjapiSDpHb5koouBtlNddDgN2
mtywS41/RqV4wRG8c1UdBkyRY+Rs0Jh5Lmr4H6xZwl/yYc2xBq8A/BmgttiMTd2o
9NBuCN8ddrkr022vVym2QTj1q/JWnXuU9YdojNPs2jpjEseIOGzEP5w8c6cMfqpl
KhtUZRWHm+s3zSOl2Mzmk251GjT91iPxmeMhha2ctV3UrUAUlox37yZbFChYV/Op
qUQZJzzlVR1ngRyEOZ9aGjPQ2uV1GGje8aQAc+crUKjbaS9mDewciFIj9iO7M3k+
LN1LtXm0S8evF6tdJVdxS2dGywYd4AHAe4/6DxQ8GjKo9gFXxbaS0UA44Gd4Zscf
Q3BvrPoGj3V//0pNglCQTpne8XXDwcxhHN1En5XeHsFks3I+wkZJQdUFnPbwhQM/
+TVQfqGpzsvPqMtez6OXA0uBytpKHldkG76e2lcOG8IxQ+UVLPe86djOmfcr9u4c
fJZGwhChzwXaZ/SqyyXOymDOhJN7gajoLoIOIxDzlvqdXuzElrfSNjQH1ZeYxl6t
0b3tiuO9i2VzqjyfRZTxjPz5J/noxsLuM4fT8MHLsahnOEIMAdvXRcNF/dLdlbvy
vR6g6X2BkgbFcq65z+K8RbW2uj2j59anDHxM/udsLd2/kQxGyQzS71mKMr/kgd7A
NN2jwPJmXGEOFVu8eTEx27hOHK4EFS+WMG6brSj8/Vmum9NL0rYqfIQL/Z3ZO3B9
xJJgO6gjCoV+v1D+S27R5dRpZ5Blyfg9ihp3k6JzYtUQ0ScDABbFtu56INFfiyIH
kaJqhipqLzGFxefAiShmGSOlKgeRjuJU/zdVsvYA1HPPiOOAbNMWdJwmpXenbV/f
pUGr6xlhW0s92bbyT6dmtsufW8DRqKw5sdVmFAmZKJ4uIsHSuk6SFfhCFFOuBiAy
d6vmfNTd32wOW/LbKS76t2mgYRlPL3dNetvppXHe0K4X6dBnYa5MNmj1hnE9eBpl
RhBTx8F2I4D/nVrbSZTY+Wb6OFADJ0qGgfbtN2u1MB40ICGjvqRHYu1i66Lc8jMC
SIMaGRGx0TqBQX2Bzo/C8Q67eBI3yLJHkWqcIELzPPS4msIkJo+7AUzVZ1fJPpJe
LHXQtxRmQ/PkfChHpXsuWUPmUHGbBMyOezwK4399drVolZ+8HYBM24oI+l5KDJ/S
jbgK+gvepx1vUk7UlKrIX3yRsnbxfG83uKoFQZtrvkBoYDdh5RjWjygV/mJCx3mp
ejhJzTE+PFak6aNBi6bAGhV6aHmxQwDcfJxjkyXHxUp3Jv+LXSG5ez1+qIhCjt7y
jLP772GsHjOWeUPYz2QjfExBzl6w9p+TPjS4rv2clMnvbgs0z19tkYKTR7wPH1S0
VhSX7hUpevxvjTNCgRjHERw2WbTOYM2bQ0Q2PSeDW88ZO7Zo8Pc0AbT8zWPmbKRH
VuAKA+dWRYPBS/dwce0XE+CliOTQ8uORbZQz9I3OR+8WVvZz+D/qs1fs9V9It8AJ
UeQkCpxqJ2dj0RTxMGOK3laQZIlIJ0jhwn/kuxEcQ231VP9934Br4etFppvDwHCj
ukvlqs27LYMu3po8i/MBV+rHagiAA/4bCxzdCg+kkWMRllcw+S0n1GBlAWPIWWwh
TEuwXmxfmOo6cNUSaxK2rk1+F78qV5a3hBLpA8HBjabHxPxsPCGTafs2uvkpedVX
JhFCv6AYTDjG2qjmOKBq2sWfz0jNZqx6Dd4tu+cqZ/1RIDYqot3p379osxbreiuD
15mmAVSbMNQSKvzcPZlxpWHmfiCvRlsObjzi66xK94nT5NdApTq25aKGOHzXhgNi
ebZehBhFCX7ZJjjauTmEQyiRCtJ5rO5UMqp5NsYMkfrSErA/YFuw8XbYKR8hL+7e
x6q/q0r3EtoEcZlHAM29qljVspwJkAyLtv9LDJA6nTTehEQwjobw1639c+QdCWuQ
A83GI4Eyc7ByrCfTlC+yVZekqrQPQNjitcJggE1UnruGwRlm2rzhnceMnUhkZaHy
UzRLap3UBT83QoIuho4Wr0LCxWyqUMoXlqF5PziXjDEz4cZ4LOCpbZQ6kqEQwLvk
U0F5EDi2dAU8w/s30Ssz03T3BGjspvZCMOD+E9/yvZGd2Q5SJo8jLw4nxf1FYOFM
sDmWBmFAMuOIihyTc8D9S97IZjMjSg8waGfHlTiFLXLpyX/MtvyZzdzIoZwhGESd
YDuMLfGWAM7hUQIiPZDgY/MWKZBMM0rOBTlqz25YClwl1dq8aN8bjYNffZmFpXDb
jAwOZUw+b4q09c7VwIslWUN3HMZeCZpB7lxnSZRufAqst554Q467KFLknCJvXgyk
BdppHUEQ5GrzA6WaAA/2PMzJljCg8/kLZkqdkzbvvbNJXhUkLuf8ITHnqT74y49e
Gx++j7nF9XE+j7YtyUTiRj+82kHlBvRdfRrh9RtTtU+ZcAHEn8yX/VrdeMaX4HP+
P7Tqnihl12zNrMYx7adL/PIqS6cFUE8kA6gHCav+6SJDsMi6jt0w0bF0pG8LkmVL
93kdMMfvh+npg2CgJpqSnDp9eVLlqdHi4zvEp8FgAabecseGbJeTB1K06yaoR+un
gFBEVmDAAFXyNYfXhHYykUnO4BlulITO/akcioEJ9xP4mKxNEB/kQgifKT+GkNt8
WGhWlbLCU5f/x0TU9Ubt+eycmukeuQyc8msPDNj9Sh8Q9O/GvwKv0nigS94ZzYSW
AdofO/MgBxZzgEJo3PF/O7pAxl2uQKZE70nbfk+XRUimFl1+MWQ2tb6yOT35v1Ew
WyQ13JOAecr7vSqiUVUCVW2j7yaY0wKhHu/6xsllI6+ax+tIcyczwu2ELLll1cl5
AGhtksimMxkxFQ9JZ+Jzvr1uoUzMSzLX0OL2DeoQ5ouolhB70Z/kaABiT2cxkb+D
hqNRpcn+2zccj/mN/xf0DkLK3PsqFzsRmuVkV+20t258PEhunGGrGalUdy87kFb1
uTU79vMvDSm46N8y4yHUolYrJhc4cqDCqyApFDksmQB/1v0Y98L3y1zaznHJ+jkJ
kKPYwGHU8X6WF8MpXp73yymrWF1eUJ6qfPYtbrA+uMmx9E/5u+2CdCOSjjULgNOv
wZ7iQD88OSWvM4TMNhwLgfYQOKH66AnTOMIxni53ZLVZys1BZt+h32fg6/toCcVr
nUKAi7rQjjn+pWF38Bgn4sTEmnncKphu53dCAsbkrxvTV5Vd1uKvtalghVK+Lelv
odVvz0YKLBrYYAVig14C4jI9ZY8lKvJevrr+fAX6ZgzCTkuQeJHKODw/Vwhe79Zv
YIbSVKRVxR+/lVH/dOTEXXDElLkng1sKfyb2mcDBnSeEjyntPg7VKrX7qEedRcwA
wYG9ruIwYYYIz3SZx1v6wZLhFA2DQmjwDbVrSMX31jHbDYWIUlhvqRinb1XvN8TJ
5Gvwz2jAQPbOH+90e3hNddBwW5wu+SCpOXDAhbv8beLLbDxo2C0p+YTMFB/+3GEF
h1NHO7aIcvDCx0Hf+wWvyzgUFEldfnUivzA5FRV6CEqPLNdPladBF5dJYHtcOBXw
zfQk82oxK91sY8z5nDu35s7oWtHDyDs72SDsHBqe2s2LKjF7lEkM0UpbJZ5kCL9f
svGIs+EoSShPgXJqbzCUKSb2PNFbCFW4mwOUJpQ4Op4l0G8SVKvZcLz8ZU3JJsVp
2x8crkoyh9eV6taQE9Rifz/XVMe3kQuc2Mrjavp6SG7e3GddY6jwvnF8qH81joum
b5qr1260fH1LXDBfhHWYBOrw3fyc9uu86gcsxWOQclpBtIQgAgt3+Wtt/BFVqkKH
DugKR/e9MIdHNsMn6NRr30Zi8ttJbDdD6hGUZJDK0IzA1FZpixFQ2g/QiSntW1eG
92Vya/dVUHXvdLZsxdfgGYCHx+5NHYkr1oIPgJNYKldOzdOZxMAKNFKO6q5qiqmR
f7ec2LWp1inIO1eEupiqduSlO28iHcKv6iq5jVSBm6tDz8NYA1QfhEl4BSCNgGOR
3eIlJtH9HDzAx2IHWx+QkUkgVnLD/wiN2ys7/zuT/rJUpWNcGvwfisix63MK2BKn
saAA6MCsAiPPEVJATieL+KKtfzWR+NDfDhtklZTcvJgK1IBhpgQ01YQtnEuNAQc0
+fz5I3lBGo1qL9siD7osCw85wuPboW/3CiXOeQHGmPijQEvqDLYPXO4UmDj4VXrT
4cXyLFHmJzHCz0bX1XD10ILbPsje+ob89o6946k/5zP5zupbzaCQxLmV3B9zYTYG
RsuOFBiL5rKQzLHYk5QEW2e5j4aRY7JlVDcHb1VzuUw+1sy0pBryLZiq8VcwEOUw
3djSsB4EsZ5hL9Joe+X3ApnFSSpRnSlpCA4I+AiAO6jrUIXRGSBZYzAaeCaLMK6n
EuJly7RlcjK8pVmh8y1eetlDENoNl3t1VNPkqZlXDIiLLvLdRpAvbHLunPr5b5QU
wfwulzNJFN1hBbQX/Vto5eSYQsVSiwy5R0jQUlBF7psmagerxBceFMaulwGIuB+x
UJOeJXwhaVPApPjS+BJz5rFPuzhMXvOr0g9J/BdP/YepPg9ceoGoIgB5WN29W94R
X9DnsH91BeJgBp819VSqini5SUygH5bFpHZayf7QJdr/Pj4hcv5qd+ACBk609ld3
FO0EwFVGntBXrxEHkYJH//NYKAauVB2DOYhErdBE+/uCu/I/Qg4ENNOpJ3Ev3N8w
8uoC6+zxl4R1ObSr3xQlwn5cA6EYLV3KwA287BdKuNf6V6j5IOTF13xHq/bHyV6M
FVmEC/4dh7pYT2VwosmedTv6U5YMrmf8VidKLP0d6N4zfXXdaGNAtE8weXPMPdbc
lS3AXGAHii2/EYUOIvjkv1R6VuUiwBF9YkTe5B3mWrPtacd9jxnZbz8DhRuZOq+h
ef6JFilkKrZbgYTC+4vlsBGIISXiQPKzwck3uB/HjpQlsUqdZZw1tZEnkyjiQLJL
Ht+055bfqlscQpBRwXmUOVpNs47mZ7hXgEHZF56N05gmKjqQZ2LBfVQFfZNIlfHU
gkiBt6/g7Efv+bPqWCiOHKEET9yRA7l8Nns2TbGXKCuuNEg6xhA3CWNiQpfCLDds
q2SP6hX9EjbxXlT04vMAnYkT3VVtG/Yqj+O3yl7ULJY82XdY0K9PESbWO5wKzdLb
qF4LbrWnWQ80V/qffVyHo1H1pYkc5UIR0pqpH72biGd4vov3KLF4IQPVzCl9976f
UdB739t671Wm1+lefaQhKIRchrXgIUgdXzIc+wZe0qVrvpvrQyNw2VMupsuCkUis
ncdC988V16+NJW+iKl6smoxbMaE+38drD57cLcMYLKyP++u+kNwMc37AdRmxaP14
4P4wq6AV3jgwTC4ziHtLi0Js0misn3M7cWYAGe1D5WuY0wMKVW5wSV72qISdEPQ4
NWNa7AQLc5hHeDJK952rRcKeZFimgYSilY+CxSgsEgjK3KKjlfsJ3uUrTSOjJeTl
u18kTjVFFw8114u3pdwmTFz/fjw69bAmbDN5WdVmc7WNYMlKAZjxQgELsSA3zS2T
Iu8vsLfPLvMnvF9hK2ALvAvrl+vTfRY4NIBbju1sFiqEzeVRFKc5wu3+ozNk018h
PhI5M8VAjkhoz0DDWDh3Tmhmh8gGX/EWMokuKabFCAgY+6pb+KkRE2U3zMCc6mVg
1fzdnBRSMwLZ7ddBrcNLF3DD5H8mAGh93gmHzTSRBN5lz8vX+CPWspAfkxmU6ZKq
bRoCdqrSi29GDqWGpmhqD5jBbPojy1rppLdxjdljmLekJT0OQDbmODBw/Sz16Nml
oomeSSqcPrAqkZPD56t+lKyEF80x03LFdFO68muYAZHQnPvfoAOvaR7UnwjAfRXB
CbzmyNtJYZ/XLQshzJWUrBIbaij6aIBH8WR1H2DFRklsRpXEd4f7HVNn75wMIFPJ
VEw7z4LHDA3hAoW63Gg0G/ddCcYX5od0nKNntXtp/RFeMdrIuQ4qhjrKkHY3kLlY
TI0mZvUbhPNqg2Aj6xS0ZEBIgc/XN5EFAf3ldGybE1bWY+mvlmo1vGSLtIo3lIdy
NpNiNDfzCOhZO6oE6YzZdHkRXiHJPECGGxAI8QJEXisAwKq6koGle4P9BapabtQy
7ucQDJgq9kafHUBZHRS+m7rvQXcZhM1y+3fX9b+hr7zN4l5Tecjc9PUeaSLG6wUS
JgyRmiBvZeS9XiXjimAyqlf23yauEdNcHa3tddxJhtXU/t3JQ5YaYVYPFux5vhnN
hz2c896x0CeBA/55gUHiapjNhdWwhOKTIpM+8625fL9V24JtG6vZRIa7ulnd39Gk
QAKYEVyehVUVo3+AYOz5Zwlaj/+ovalYHNurDXx/D0im1wAt/RYnF8KYeHOyJHLK
sh/UcBUijtcljfrITWhpo1LX7miIX284YBtRByKXrWuhDj5PJTpaMRFjmQE3vkMS
8dDrsfgCkakSGX8ZfDg/fcCinOFv7Ct/GxoEh1fcXnSkbicShwXAauiJwCb1vYc7
iz1P7ioveX8sB69ryhsvO8L0DLccQiKZRLWQfETOZHZhLVcvt2uyDMlDzV0cKRqg
oavCC+JmCTVRm85KehGMHVdLhnzCuvpcc8xmHFeyHOlREOY5hyRNGIoUfDvDFvTe
Vd9pRr3hA+ogtw7jUquUBvcqf+qHTWlqZln2PPEU6D7miD/IypTl90F805IT9PQg
FhZS3tNXauctZA/nHPJEIRV/4YIGMofKY6qU+o/6+iXMh3zDhUY8TFA6DtVFFVPP
KzSH/w5DM/p5TGT+4b5GtAj+dg5I5LuHUdf1r2ZdXojtTDUhEM4/sWh35K/D6PvL
9p8pOgh2feoYpQnCgFP9YDA6ndfVL0+WT5E3+qVTS+gcNQPRy8QLLOletk3DfZs3
7ORxoz43f+NhI5Dtm9uLB9zdN4AT42wlrM+kipej8PpdGBPhxRh57IioAbh8BmCb
h1HhkZeHrcCJdVzSNgfApB3SeC3Ksf17UuWtCFXpgc/sH83Q/PMM7GzCzRO2td2d
+zrQafF5v+FsVskveOld7ZC2t40xNoIamV5SlEitJ1/qSpEAuEXnpjdjMH6H6wxO
LUQz41Veot4X8wtu7goVXaVLQc3LtQyKEFAdVB4cBANxln28zWdaPW8mtJs6OSbO
L9mozqmOk/gvGQTcRu/tup1gfgPeVoGs27hYjl3lvNfiORBI+bpwBZ/AyVcN9ksS
oAXX1D5Ae8ZjL1AbZJbabNVLpvFP3pPxPcJWlWuSXUJ2D/+m5A/kQ+L/NLmg7G5T
fTnU+WZaR3MJBV+xnKdhJ7C7XR4QIYxvqf0pjYdbkFkOJ71e+RoVvD/INOKfVs0Z
qif1XULtCCm4izIvIQ3ftbv4guq3K5tcFs2Q5XkHzPumgBYjb9Wv8iA0i3CKfjpl
5m8fiV7i65v9d9taprrkQhbt3vcd5p95vWJ+FgFn/vj+mGlUQJQmfbWDVlLEsBT6
xYF3gHp9A/bmM8NC6bQww0Pihf4u3JtNcEH/Fq3ihjfA42ym9BHuJ04ewnPEyEk8
WkjS2QUINWXfHJAYuo22il5Ssj8+hCxBxIKBb8+urzk1ass1pQkMhnTQvi30J5Pl
vGTyRYoXUw+C4sok9HsK/GrYf901GubQfnQKZKNgFTApCc6bu0o8tI2ljupsyfzb
+x9NIFb1TjEn5w6pY54/pYR8Uk+vObD3mNtz09d++cLxkt4Adgxz63t/m2/QkhZ5
H++595vAjsT64jtvlHwQT41waRKf1Y9Sx1eAOBLTyh5dPNIq2cw7zbp9Xh3bUMAS
4IvG1M7LtNZv+10PVxU1E7peFfamfpBuONVXecyg82amrPFDk4eTEAhUxtvpOZC9
9cg60h8CHemSPGe9sqte/Do5Tdd/5qhWLaeK7I94CfpokNrMuQCnENg1GGifNm/v
yov6mOwJym/pUdNG6+e/jXRbHjAw7fEK9KNHrr62joBbZyAgZ6d7KIZKFYYLKA9A
NXgdjPWbNPH1gG+IZ2DmlRCQcgwIeJ0i8iGhppwA1YioGQTnpf4l71Y5PNT1UE/k
cwI/sGH4xUl1JEh6XHX/Wg8Oa2zME5V9SzQfWp+TqZHTsZ3eRNWGfnjuGxi440CO
SxeHrX5oOriGVsiCMe0xhY0+ZzHn0JQ856TKcy2fAn6ZRhsUg4DqMJHADl/hFLnO
+r4VL4B6Jx2oWG/XYQpiRVPqdLStZ9iVSqjyGW1Prb9uWnOS8EKQTNnbczupqmhA
ffKE9hlIu0EUpyANpAVHEK2VAGXm4ucXJaTs6AXZqQ1zBJT9hwnP6TIILd0imiLj
XGR4dhpblEwKBUXd8KuQZOFQThtCYNYn6imVnHAhbZ9st3qJadThGumu3Z0mo6XX
L1mjsucp10TzW6Hh5SITopOvOh25sXZAJzpPb4G8xlJMK+62ErSIVlPIhUkvWJsb
0Nf3+aJ8MQBP22eXrAyRkdorhwJNngbzCZ6DtxAiy4RyCHcpjTuleUF+3HCCGDl9
fl0hI9/EtD0cfyNpXbBnpTqKQqZNLGuH5v4zYtIDVWrM6CSyP+H4zV7ApC2+f7nm
xu7UvBiPB9mKP56rkEL+e6as0GJS6q72H099q18LVAjb86NWvCrlHIVw8gWq/Tfq
OeAVzIAgfBZVDv7QnUgoutBOLqZ5f7jOfeFLTDBFFgsLmvI5Rw/yGyrLwv6SgT3z
pSgTaJ+6hhfiU1K0gq9oHWqvcH7UF8+prTXi+Fmz/1cW17KbBnmUF6Yg28b/wvyt
zoIksG0FbRRWHxBX9e+e7SuqIvdjBPANlPz7vi5HOUM4poUQNwWwjUz4tAz65A/1
uD/SOp5Pp7ZcxeMIAX0a3qcNoB42EblOhK6BpvrQsKMGTB2HFl3Lig82dZ2ylVG4
2zLLNZPsTrRiImmmDlUCXuBawYrh5L7IPhhPifm6g44P6Rq4v7LHPa0tG9TPOaNG
UkDwBF57otQiiz7mva+E6V/pXFm0LnZVaZmMxx9VjkOUuX4V12QbZCOmXtVGY3db
32aIgwEsRe2ngf+KZTAbG/VSsr5rEeR32EQACqW3hvl6LakdLCpT7BaqWbUftNJj
jBbIVWmnFiiE55hehNiuBmduq6hvxO4A1me6sjr7TX/of9MjwkLzpgpYGUKThvIr
ljtpRB7oKRFTbQcQnFKlQ41mFdvs+I5xiDev8qbr95zZf+M7DHlP2AWRNYDW2CiD
/tMjk0B/8QgAK7pre0ErkReYCu5vvi4PsDkYVJ2U9fKJ5bwTuSENMW6Z1TdtcKe6
SIvlDdp7XfufRxEtidCbRFPJPv6yaIKboL2Pnp18lcy8SRTDZHF4ntYFKyny0m1P
+rE4McMq9lnPvLyjkRwM8g53GfJAyhAqL86f8cOnJa2ji6f9AYeSNM7z8/TyyWJd
Ovqt/Eyu9Hy3dzRWf7XBpEWJLQNb24/wNFE04SAv5NbtqYLYSmYG2DB4uMI2Dq+O
GEhWFtC16klA6keXLPWRkaaU9TPCSJLcVCPEBKcNc/xNtXFDl0pK2qqeWcLgS98W
1DbkaBNY92sSuOVV2RNmCDOZLYS7U3lV5PmKSgFtsOEpK9mFySplMCXgcoh7k2Zd
ro2ClJR4cb9Kxk6GrzFwDJiILoMUu4ZIpFYe7z4wuqjkU1l4ixGzghJftlBXfAqL
kETGe7whJx7s1ZSTllKLviHU6V2qA6Cxq6WweSIVuYBmW4s+6D9ee8/rRJUoXL9D
tBuAU+SHeO+mm0atjrxRDu961ybrn6mJxtJwVniMvVt3W+Q6Iyfn/RLvqlvCIGir
NkPj7e4XrENueDd5NnoU2pPH6X+2fZhEpZQ69fLxMuWHrwiprNMDuEkv0A43ZRdz
xiPVcntjlZ1icKx0dP6xO0SKJLSRoYEy7G8T7jfVHlYgHXgc+AvhM+W2rG+zy6c7
G8C4q2neGTn38xtGzbuzsZXbr2L9ZX6ie9AdKlGgOS0RA1vB2EYTA7rTvQhmLZAR
6xwjVHePn7y8Qgq7nk7DtZj5QqjPu9nBv2DqWvxtZbgBqwD2OhkPSKXVJbF3IGXM
fASjLa4EGYkHWUwAo0KlkgR6w3+rqUSDmPMY0RgEdoCGbu0Q7V9fuYDZUvHDAcJu
zb0wvmUeDnPuWFBCW77SXoABhNXs9Ai2dyF8Ka+FRyfFyzYxaH4a5GTg1SmXrdzg
tsgGlSLhwJf3GHBZBJVqeAbTSnqKnQvGN+RgEFHk+Ir75o9V2gzH6rVnESlmHtjN
njW/rfwmtjvVUvu53766VWTj9vV00EyBYN+Hi65OeMSlaf1K3nfY/GOhCadMVs6e
/oc7KHnuPEpdtW85BhQzZICGdvzrEaL79nMLIurYiG7Hy1OrTT14oIaIvR2H21hX
mw9uqDsSPC0+IJfVZYOJ86a/KQyKxGNLJhQR/Jqv6Oo6fUVbD7fido/OH0/tniPD
nuT7N8+kjSnqombl+Q+OKyWGJpYVAiHY+r+ulFcI4brcHhHqoTieAr5Vx+6C4xYQ
IKDt1S7myiAE3LH9wfCu2cGuOxLvysWuXQ6K7oy078IAxHs5gggeK6paf5E8Eqal
PkjEQgarMoTgvpZPE4JIhe6QPzFZO8UsKaXf/Bmh9d6oJOaYSHeCXPXFH1Rr6a9S
jPRRIIqTatBhkxkE+257vW8o7ZHhuapHOJpnGQwbuWHOwhbYJTnyPhz04ZItk+vm
8bodnNZKmgdKKgx9nng4ifaDcMaYPIhIjiuyMZMkm/XL2/7jzYDrwGjVgK6JbtKw
/XDloXd0n2Jf2TQlx+Kl8VCpUfZ4/n7YOgYkXdedMOTvqZ+kzUtJ4iqhmDbfqkFs
Cft3JB+kyap8+ryUhxU5VOUYKQNAj3LoXWsHcbSzDjtJrRK+jLp465uCd/NYmfFp
BHmANARjWvNtZgYXetoM5zsQEQw9jbE1x3C2j0pQil3bYynWUuq4UrN7Rnp7dSzd
fEQSBM2U1dkroo9S0c/PdnMkf1jj4cW8TvhZ4cY1LNI4unCwH8x2qO/tEP34+RMK
ArIuzQR6iKA7o8z2UR6NuIanERm/7jExsZ7cYPxXouq5mklN37CemUMrIrSriE5U
3Iw4W8rbl/5cdllxL4i3HPAUM32TtkkKkZyaB7WporR05D1IUm0Zd7yS9HOjWy9r
RZcUaQDbSzrAmoIB6cuMP1UASeoTEcLS/AE+WCBhFamoPQNnQAcj0vMJOvP0miFf
JTvprCblcA6PJF9ceCxY0x4zs+v+EVK9C5KJ5pRQsNdYXnT4/2vMecx0Z97PNJ8Y
b6YTT9N5f3nGWJ08WMoVprXerBDTGyV2ym9c/roAzVfrqyplcHraoFWwM6eZaGmn
B9j6yfLQUqNuh5aZ/EPmC3pnUK/ZV5JFehZff/TBSIMimOvgwPklSnArnTZQF5AW
kWE+TckH/REygbQ7VNaNzIgTPUzc42a0vN4IoYptOl89lr0sLoExEgPYDAvLsl1d
ApKN451I4MlgjO9ghT1Kk5mfflyqDmU4btFzKt7OYb67Y0tgOGz0NhhzfhrPDW0f
BG8dBwyClGrZl3uyrcmbZgh+qN8r2XW19Jx44vXWuG+AekUSqCpKHcHJSCnbCX8H
OIJOGXqLTh1dWdUH18f6v2EzJw+DKT/kHA2fK6IwXdWksUXJLg4QwVW+0HYVCe10
V/fz/8qUFfMVVQTKI3bnw3niL4sJVQtvs+zRf0HndvbuahEcrHsY50DktrLLC3Mw
VzTh5gaLLu44QAtSCtrvBsUmExT4X27fM9CLy2Rl/ZfXKNaVy3NKblmNTzKMOCvj
UaDxXlgOfHDD+5KUiBAUZDbNaulEeYOIL4OMPrKPavlcctrSpLHmWuEB0KhPoEJF
H+meE/Z7yO2AfL6/FDSykXsuJHxujm70GulJ9DC0WghSgBzN5NeQzPbk+z80RiQ3
HSoIETiHl5BI+/TSTZzyhlTzl1lhAaGEp66ECJ2H6gdFNC/9GscLW95zsdRdApQs
/6BOSbbwcR5lUQR0oQVdmdCE/7ooIDG2leZd6dz7KuMRmzM5dO9R0vaEklVZYrcq
pXM0+kXvmN7/HkdOnyONMntiqvEexTPfmuKnOVzviW40DuJPR/tmtuo/ktydr6nR
bmlQcghNvGY3kekxuKuUyar7gupc83nNWHgkVlJdn27hFvNw5+uemVgu4slC/yoW
XSm+Csp2cKv2zygi5+u4gdBI7jrcxrDFPtfvNUm7C9FNEe9CFzCvVrxIK5C4QEx+
MArAYra6zt7yfDEnC1iKTW3dYuJdQb0x0Rjw/GyueltaTPxy3rty5jQLhZy40cJ5
ubxjIQX+PT08LNbqA4rSAPjTM58R3bJraRq6S5WH1kkPbQ+Vzs26ccMiSjtknfv9
TuQEOcSapZbl3O6vwzxWyfZaGyI0FNv+Aor6s7E0wziK+WthrDGlP0QchdAbkpqL
SYSmO18FEgF8lasppwgd/rEAMag+McyoGRbrSRvFjY87tw5ICZr+78yoAdVduhTc
Osy/x61+WWbDGFl21Kw2z5NyrXtvVx7nYfL08XQCfunPv0ol765J7eHiSnG5qi3V
kxNtZH3AN/pQ8s+TFW7pM7DFeR6meii34PKyFqYRS36fn4jOXPOyvY+5Oia7C8iG
SHF6gu336895AUE6pF/pefRz8bp3XGFmaNFyMWoEwdBnjQG0FLX3H1/X9fmwFeAj
Y1H4kmwCkiZJ+dic5PcWS6wM1bt8EafUjI2//cM5EOV95vuP5I6lHI2C3U5CUmST
dBsFe33X+ovRsEpTl+qPOoK5vTpwzqjwDXPFg6ezdSe+rBDF3nySOZiBD9wBbhZ3
tY3eE/KMPro+m9IoaTZc9bOVrvkydi12QpZ4EHtEU81ApeTTg2Mf2rw3vEAs984f
ajVq4K5kNqk9EXOhV0eV9kWq1MZ0fi1d4LDjVfk3MayOtfM7pyANGwaf9XWgZvDe
SUExrU0WL5dWyZ29Ia87kwVxqrAk0BkOu2pII0BtK2QfrukayXlmjCswq/buAT94
sLxPLonm2Zk+GOv/z8Ao3JiNVu9TCXDTB7Yys3Ip6cMD+VkN2oUkPnXiQGRfCIx3
oQORteXut0hhRWvvrrN9we7nTt86AMi2XccpOWU4jY/mcX8SnURdhZ2lcRYTomjB
m7dBPiNmA2eZrtDxMPztswZluYXwjku1T4K+A020DWTKreRfqH5JzIsPQfVbGUoR
y6/ZKkTkxoUWwL6kCIrv1RPd8DCX1EHQMCZi8arI/TBsOK7MtqvYuK8HtgDzjH1Y
gzsB2IpcSfwB3nLd+ropS9jTOz0hbJBcWWP6bRoV/fIkouPuFbJEAEs0T9VZaAcr
PIVQl1LooFErQm+V07p7ELm5bcLBpodNhevNzqq8W7oBXM+oRvPqRaY1TQGbimlV
ssJ2nIui7Ah9X+6ARRjAorCGE1YnuXY1B8nw6wHgtwn9NciBibRPOA/5kov9+z56
16aWMIZiCzu2O5oZLk2wEaYeQz8incRHxar8956ROf/VFCfTGkA7ltxi859cRqJj
Ta+cp6+6Vihwk4oWkczZ7DqYf0hx0ZHzAgQdFwMZYlxMITUvLASdCazePq098EIG
QdpwkobBFN0WjIMLrW9hc/SKbm5W5cdSoOJl2sV27v136r1UaNdta9wAS0pT4Lr5
8SbUPlkIvGC41xxU3yhzWzUNdy3UFN/n2Usk59TlHSN+Oxbv1zU0e8zGgD10C0Va
jZxuUf7RglWxfTRuJ0s1o11S2gVCZtZo10kQ/b4rj84FYUTL6NkQnBDMfLDF+WT8
5WOUx34ro4pWPmv+/VgXsBOf7lmE9gUIWXz6eLjpUmIAv5O11cjbXTSG3Ne7a2l0
um2mUDN0q7dSFlK4aO37MEttNual4vxLXj6FqTlUItnsJGQTdwHwfxVkoKqoYIhi
rUKzMdOE+Gy/D2+NuYa9LKytyTEVsk8MO7uDmyVmmpMHPRkURkDzetRWa9tYIxaa
xYmBBS2QrxaV+PaJxKb6E3ySCtR3LNG3LRUbnn2KdJONghf8QvWm+WAVuDPh9zzr
z6V2XhfU9D7eW2tk+J58/aH4BMb0L1kE9T7XDNr27Ds6wuvbkZVkD8kDEQ0xYcqJ
CE7xpR8UG55JAALblFss3eA7x+wrII9qHY5cD1/y8BhL1Mzb8FcDT6566GALZlew
kgYuso+9Bx4n+YYt+AiOI2PFfKsPdNYWc/XjU0/ZYzuJ3GrM0qRnhv1mNHdayyUD
3hio8pwdoicfXLcgxzyA+V7CkRfF9lGu0GBknmnXAfZq60TVwfUm8mgVp+H+WLXf
UiOxcvWB1fzA58EuVrkn3meSbm2NPUTGstcojBdi+IvbVWKw3K6LDWF3BX68QLXO
1R6k0Zopg/NNdbxNi35WynDr6pCbzLtth9/8dbm6QnOUv+AOiw/LaZDy3Fw/cnRG
AkPsS0nEGLiYiKhHlXYi+Sgrha3LIxOZOiaj5K6A/gJdeKkQ5zlXjLD7BIm9N02c
cjKMZSwVuAPN3sUfUVfVOFFtFRNheGjA2oLT/h86K82/aJsgw7F07NcS1KTVWpd4
uhuS8hDcCwaC6M8hpq5dzG84XsE1oKRkFoCZRKAiTK4+xuKPoJ+fdxoafdJiXBhd
HQU21X3QmcCakDBn/V6dOMEiPL7ITlFXW7ix7Td45fmqNki0u/x1xt0VlvOmv5z+
MZNmUhH94wQwdfH8hphBYUCeRRolZoH1OMtwsqfxfRycNv2SoFyjTHfefOCQmO+p
/nzUg8MGJg49hh/rK2EKZsJ4wKeT8riaaKs5OziZcyLta1vHrIhThUEhaAtup3BA
K9Gf+MrgJDahH35t43BiMRy/98MLbkngGvL1SWWCtWULnbWwRvOQHNhUuEex4c43
Vf87tHsUk/2BerBSVtDlmwG1iDbvqmE0S+/x4JG6efow0y7iaq7ehSrnSsSb/Hks
EDK9wx+GAN/wTfFysHSDPlFwJsfqnddLrCPHSZZBoRJfXT/0bifCTgXiNtAVoxeX
195TLOo6NxuuM7UzrjRIouwLQkQ8D0dw3QFmZYMPVk1U1+OxmKrjZuciEaPgsMt5
Jzo4PxH8zCY63Fc0o1jJMcDilxFcTCiiK5y8wEaZomjIOM0TVZ8JHDFntvJ16p0q
mbyyZ6pQNKiby/1pNpxnjoNflO9+MB1uxP0ykfSM5kK2blFjnZ0sc3qZ8Tk3Dz+9
tSCHLEuUBe8pcIdg4kukbk5IU1mWEur16bVYUSk6t0IVdhNJLl6vnlvlYwz7SLsw
eTFgbTnStq982CjS0cAm9IrYDlZf4Qp1oymEm8O1kBGGpqVWcsReyYMZex7W3FzB
Jo6Rv4f2dgW16Dcr4h4LfX0Tp0+Uw6rur+prfrr9wQV+O//3vvD4Q0EkRBpfb703
42PwK8vOl/NAH/+9C87J1lXLqycoCy7J39hnoFtTIVt479tE1ae6Zgn46rGcFu5u
q+fNVnLnEFyR++GNlNeqJrK/CuJuB5cxa5xR+BlGjTndSb+vb6exzOfhPsUqhuhj
L1PnGzr/Zs5wq/fzaefN/3Uc5oD5A+XT0NBGoKlY0NOgxuZDmFUpiDdLOrz6YBuJ
ko4V3aduWZd7pWDuBlMRmuXuuo6CEBS4sAy9KZG0Nm7h7DexiP2BYfpiKLyKEzwt
Aakd/cXvud5cWfulxuz4gpGIeYn9rEg96VpHxxPUjwWNaVq1KPOVNhs8t4ArtiSj
qONFich7/Fu3ufAFEibVHUNB9GwBMwelOAVssUAiUHEastqpbAQWjNJUfoxVXZcX
UahsNa2WPrud7tZqT/KEXKpfJ7SUsWIsz4/uX9uQ8Y6QMKTV2M1vl4KX2uQ9UHpm
c8XnA0U2Pz6y/679lWo8FqM4XUVyBAzLqvqrvT59vLHioVBJDa7t3/M5MPaR1Za1
BTso52JhtM+zVOH7QBSrJgjwNdThJdNq+Wce7ScgOvAY6GRFc6fwqz8TZmcNUdtX
SmPL6DNE0m7D+DNry2FcJ+4tXZkLlMyqEc1ezrC1kknX3FFsrvgXmJE4Lyes+pCS
omsniCDDTfZ/NVEPq+56xXxrcTPfFALDOKu8u3ewLCJIqjzfri8/5Rdh20MC9wii
K9keFtnxDDkaLZ6HOk+O1cr2WL2v9zttiUZ7IAHKZI3+aXjBBBE78uZZv2pvRORY
7R6nNAPRc6PfbH8X4Z/ka/KCUZPQQEYPv95WKYPjcV5xRN5n3wNpBL+W+owXzKoJ
018LN6XrMoyrXxhXwLKb3R6kTYqJ9Ev1znZXRfOl9DexasgzGXqeUY/EYK+9a8+4
6pyyv6/rHhWK/2/YYeix+rhcL7gvnpOavsHnvEjtePtjEvOSAHI3IhP63Au9BpgQ
TyeNtEbfR0uEawp12NTEjUlQnoZf43UpE0EF7PBJgjf8uWsYFE3Bak/HbWdtWvZS
z1qAaCoMiH3A9mGS4yNpZI3IOgSqwQW9fC2SKEsNP9Z1h+wZ4rQha5DTlWcLG6Lb
Qh6wfOsL2T5YA0wQnFUc4ZjJAtiGke3D48lYqrz3QtgL8genvS+ANiOHcTaIrR09
syZL+NmH4/YQluMh6VZ7WbH6nvShiv86bb0C8Xxz1uvy+eAyQkMtXOdf/mnaYGv1
1wWrnRitKCQ7Xy2+UjGfpDBVPv6gGnKJ0OisEskx6sb4QVLOtWLMBQkG+M36O08f
pgJA8ER21XY0TQQnPY/fs7Zjbw9uq8k8f659Rqfvj6mHtrSot013v7MGMsR3oTjk
+GYPqOA+mLZ4CDkJSr8be5IW03/2LzFvRrQPw09TFEracc0lOEpCm34NIrrJrRko
O7jnIDwCdUwBbbeDK+GiTPH3+2C+RnDKVpdKLriUvpKuW3mcLR8TarPmDgv8ZVBj
HngfzH4Tj7wzuo5vtM2hT5MOPcrAa+u/Hf4JvY0DmopNppcHFUa1v3rwp1nVHTn2
LxNih76IFeM5NBsX8+Y2IAVEZBbr3Dz4Jscf5SHDLW+iIf+mljpdvLMQAu5Xc7d1
KtMB6MKLVkv+TQcqEy8ItvgpQXHz6ZkqM96FAOulxwyt8/lPUc1gBXkqnO3b6wd+
LWzLAY6/W83XPshzrBW9kovUCnDcQvxku3EHNVSh9/84nL7EnNL0amBEDvlU+Jyk
3yWnol1byXRO840BV/dD+2DLvUJp19lCkvGMOpMjEH5Kz+PUim1L9DOFcEDTsFzi
Mum0E7J8gRQZZY02/JXunlTFLf+XiQZtmNkYWpRmge2jyKdjVAt6uVIOQvJBPlm7
gtffI72SBPUtHh6M65iudWVV51cQpY8vKL7zDxnSDNXA9zPmP4fxJBZCQXnAiWe1
H+bEI3zvHphiYPTHXt5Hdxo5dQjCEsUoNaNzA9ZQ4KCj1aGxaXqBrI0wXXiIFyrB
bQwpLICVvjhrbnQFx+fAZjap4lAdAI8cSIn28Y+xW/e+TON9aEpZ0OBLgEK7cAvE
PYy1FpQW/+f6Qvq2sLwLdk37eiYb0RAO53iIiSVx680bN2rqm8ORt7l8fDzGBpJQ
vvWYFSAPqtDtwThKF4KxMgNzEChE25e6P22go4FBeRjscIVlh5V3kXueMpoOJw7D
/mJq4B03t9XjbCYM6IuH77kQkDoIFJVKH8uZtXARX5fXkB4Nq6baSmI3DG/eyh0S
5e93N2s7UGtgG5vrM0fjEC+NXHOsXlu9/BuEB3k2hdq34KO+uBYSNKNWd47mjj6g
7CO5L7JHiKOHu9EpiukaMW44GizCC5ApdEv9BOQfOqFP+TUHlXnRlrJAsR8cVhl6
UU0DyPY3WNXe7UqFTz0caEjL4BxZBsq9t540kRzX+T3rMe/otullzOifBjaOQ1ZL
58J1e0JDxZu3aYPVA3H0LVayuFURHLFfrQxNGVYDCpo0qabUV1fAQhYlaGZtYLUB
wew5WdOQfr5vqD07C6XNoDrMqE2KMn6NbXBMNv5tB0HbmcjodKRLGe2bgioJIr8C
IiHTPK1rU8xwmne9RVZGyqIoqzlZupwpp/cvyW3Xw/avyDXd8p86DplltEXZqTK4
Hxs8wvidfxmwvYthb6p7Ptu/oDAvsOmrPVQ/Vi3mcvPr7Gn/og9PpGo1ovn9ramS
QsZSNR7/ncbIEYwTzLtej0Asmb3/XfQsn3Vnsh+o0ABdmdcK9C1wonNP32i46Oky
JUT1oD0dX2sds4jjKjBtu7kj2bIVvLG4eZMPa27zd65MUV4QCuWz2x8Glit7ulOf
SPhEilr1r3p3DQQQ00zNWmEL+56qfHwXYVuM+fHlRcSlBN8R7zZILGmjFxp/8ZXS
BUeCtLi0DcIhNP7H6xLv0hwPCDiwGZ7PbPTliZov0sR4u55nW0InC+gwoKjuEpye
XaSg+69nVzy0tEle1SdXCt/7Jjy0oIRNMcvrjDOjD8Lrfl4w2LD9wrOXv9BI1M/r
W0rRvg98HmCXCl/AznLxsy9g5GwENvvYA5rnkATbVrPKBECkDAZibg9DoOtv5ooe
g+uaJjtqcUmHO0rqSMFGlGSRBvAdsZczsy1g++tTta1rxbBSeIpGJfnayhv7PuM1
twzWAJ1wrCjatGsxIKJ53kWxJm+qMFbjDU+anZt7s3z22oaZbOt/qM2aQ/04Bmg5
z2smtG8xHIb+G9e3lPSEEL4+s29Wdlet8vYa7SPwnl9xyaWdC/2Vx/4qR6yybOgK
ksRUheQJUTVfs2oVWtfipryaddBUHaHOWeUiNrkHYGOypnzlE09euzoOtPoKN+mG
BbXX06FtUsWrCSqmpn9w2UEEvpbA3znkjR2IsK9sHieeunam8l0srnjRs/kE8YEk
nX4o9tPOvnprAHRLpjHcGflFdF1jFeQL7jCqNL9T+y/rddAKfAmhqja1rMAUvRw/
2f8TK4v4VcsWSgGC/YaL1YliTUSiPaHwRhnH/L3ZgeC9slF8ePdTfHceIw4bKxIy
zNmrYCloJoZ7X/bylP0ntDyHJwTY/FSnJ+KWlJXnzikvoWagOtWfBIuYd0oJEDbr
19weHUfLhwl4chwnUmK8b1PsxoIwrvQhH9G6jSTbrH3yoaKKI6VIoTH86KFIBLvA
SoIX+OHCCoW+9YzkYG9P958S3TM0gNFAB6c9HHoYLDXLyChJivQE2iNdQfMZsmJS
Z+D6cn35eRkjtnhk9krlS4/yDFvscgbFey9SisBydqfKFOpqWFgywquXu985x99v
fdak1/xEOsX9XcuFhnKREOp01hFk/Nz9hMs/9qAMObaNQt2UNtUv1Mo/raxbAMFn
Zdk35f5aUogy2z4Ty4lBlhpZxC4WZnupnOEOSYsK1Zdjcwuy4+PXghlVtL+uzzQ4
zp8UTrzM8hgoSgbHs7OieUS8hBRg6IZhxNlEQGh07aHViZdmIpRyo5+x8vqt65dS
SvLc+04z12OBuDADjt4vfs8jZdLIrOPx3h+1NTVFQ0vOm8csnI2+8bJJw9jV7PkM
43Ar5x8vRr3w7/ACJGYA9x2EXcyTEifC/4LDkI99zPN7XXc38nQqHQunZ+OZkF8/
VqxRxqmhhRNx0UqNbzIPsxDgh6RPDRQiLduBRXYMA0FgMQe6LF5gCwgrC1s1HJDV
A6TqHRRdGV7/6C8YAd4o1O6PB6KOpNcIaOwIjChBpMKtygeHKT+DO9FetKQ/LqmQ
E/1inNZRzApNhZ2G0nsvCyVbyAqGdLqrOFIm30Ya5ZY4QCvYK1yJcrPWq8SPI6Ex
6gZfbFgaGOGfz22+Z8k3mGq02qVWT/wySWw+KBss1+mlEvVBQUGKKgrTvH2R0OLt
x/NVfaZKK8tDOjCJFonsdTEKkIEQKfV0hbKanx4jI1qd1/On5tWf/XDKlKnh+RXI
4lKElNk+9GUZ2qK3R5CvBCuoGDicxUAQ5yegrxxrGTUWHxtWVsyJJYjn5mphGSwE
KSz+wACoohLBcBHCyYlzL16VtFpcoK8MVvQMprSpsPoaHFKzJfH3bitItDzK01Rj
PFidXUv1hv50lhtzn6I4JIYVYih0AkYi3DkykrDy7wbB4qEefYu2lSHI4qsB2YUL
nYwSAd/uhQYsuDcsGvUG3ULQxvI+FhQY1elL4HsON/bjM9/TD6Aw4AOPVHSHAlQY
+N4WhMgsUwNZF03UtWXQIwA4+9ObxM1mj646SRuLzV21/RfEe085E5nUcSBqy9ln
4KNrMqDI+4YbN0dXkyhoU8TX29JKZv5/u2RWD5lcjNTfHl79BjjGUqjcsNlK7+vG
mx57Xuv/oUvBRk9tuNx9EEQbFkDmWfKKZr+2Hhq/tp0t7tkmfB9bHjmNSdtVryLo
5nk384r9cgxAcTJa8TiDF0fuIhm+633X2r/960pLGi4EHj6/cHmtKDrHTO10bTDl
tEiSjCVC35iVXh4lhOcTmZZd35EiV/yM7mOdddhchWMRi/neapOIO7YV+kdMNqWW
jXnl2f3RoVi5YCwv+IazAwLt+yaHCs0DEeRROL87G/CDeWGVUIIRRkD+xaFNQU/6
Wpzy+5FfSkpEtvH5xSTfzQz4Aa9IFUxLLJ2sG2V1GwZIu98lqhzfzzeyHEzzjcZP
YaW66BMGkIwsK3PUBOQhFqKPrSrNOpdE3oD1pNZQ7LYRnqXIBPyBL6OIBJvFicYq
wlMPn9JgwjcG2To6A9YUpaKDigfq1gZLilHEyR3mfcjts77JW203YvRVKaHcBhQd
+ESxs+FxHZccduhCIVymq9FVOci2UqzuQv4/z+vMYIPJZFu9QknMynoZLu9AGXi+
ftv+3VVzRk5BJA2DUvHXxwvW6LCfMdOCb7UKu1iDQhiHkzJ7wHd8qzVkup0rk9Zl
ZPZtWzj+xgbOr4WnJpPYpw3IVqfm5rSG/nYkDS6O9Hhs9AcfJ2eoADFuGZ5hEjoK
S6ezTzwyqL16GGYflU8DQaVelniBCj08aYnnyMY6ISrpoeIIqwsBAgUvk9jG6MvV
eub5CiyQRSrYbfoeEovPXUXYkaSNyt+wh3+ZDx5M3bAHbBA3sTNLs1kShn36zWFh
c1mViHO43ZAYHpry4l2bHOR+HPaqnymyxKg7mnEG9/X/7+jIj9SRB471BRq8aBKa
iAOHP9ma7AnYrMh8nzrQYFzSa64mbczCaWJ+NbH8T/wnzTZ3/G+0bcpuRnVpc89w
yYRq+cPc9Pi9aG872QmLpYd78vfp8g7LiG8fbvawnU2+xjyep+Uuq1hdUSnB8DWg
4INVKiS5ifglOAn50NmLaE6WLUP8xqYYH3cOu0iOlvGZ8abrp87n41Cx7Rxraf7d
H71vLj/T7bFVo9Xrf1QkJyVAjXMNmpBOAa6nPrm4C6MiJqe+y7Q7j9YYIzgpl+qd
YbtVWDZwuQFCneZfRS1IzqaP7y/nAIU00i6uI6wQwiZ7fzEtEFcwa4Y17SN8TIPX
u+s6fCB0QCqoX5gKWRD5oz3Xzo9ZOlQ2/9ZdOTCH5c4ySM7cGQ/N9+wi1FwWEs4v
lWE9mjlaqAHRqIIAzjYk4qBUKldjm2KJVKofbLbqmUpeQwworY6xH2gFvfbALjHG
ux18KFmxTYGQxdQftgeyBAubel8o5Pn4yuhdCjcYIcTUHqhRPvlT2cPw8Pp1nj1j
hcESupAO+cJFtAusXlxsusoqvO9jyF4L6juRETpfhAy9bRkSZ03dvhC2CY23VKRu
fNzoes2zjUT8BqSW/72RNI2lGmdJfYfyff9/b8SKP35VjEGdDlItnzi32piBVcBB
pa4dZ0m/Q7ztsQIo9eeAyrB8sz/XcH/RIlN1ddtlL2Ni245jkucWrrA6NdbHfbgq
Clzg22KWaTjwbNlxfOB/j9T8KFxOw+tQUEkEz4YMFzqJhIAXT15O0yc7bzWTdEI0
7cmCEQeM0uE2RYPKNciCc4YKdlqB6YNNMf7Lx5Wlj/FU1Ehi6N2sTbyhbgPLcLPX
dypRb1oHzO6EBB83Y2UhrMkhp7/8u+q3qP1AH/U8br7TgGiNUNZm9qKSCNPxvuxs
0Rdp+4Ex4gkHKTQVsb4IO3S0q8qViAcNGa9LfZq1q3iueBjQbbiN5Twv6jgp5Nir
TUNDRM/6tU0L8j0o4kAXI/0+rrV1uUkWyqvFgGBiAW96usJeZcOW9LkQ/wh8m0R0
vJUMI1+RICDa4CPq/djdd9IYA+Je6C7mJ3GxRG+ut753DC8tDSaPl5PszY3ekUCJ
ctda5QvQgkHyt4fwWO5yTwGozNS+ZRq37BneVqbhstKiVYdToQv6LjL3uLeE5jrh
q7Og6q3VeMV2pMWQjz9Dgb6DepYOfL9wuAbS8YFDKBX6JoaHn5pte9IaRfwbtAs/
QW2IPih1MbPNkGx361HlZiVJmx7vxrHqev0fwibakr3vsB8XtWMZuxDsqIN6drjJ
wyWZ4fkVhwATyiqi/2WCDm7qB1CwlH5SjxKO1on/DHfxq6UF+x0D94JQc9GQIUSY
51wajMlo0BTsET+qcPnQaAG4Obbjc9CcSzEWC3sbeh0NyPyrAx5dwxtWxqysNNos
Xf1JSQ7dgZhVQoQaV7B4swnkxXHVrMLxd3BvRxXl7q3+TAYOs/njoBr4IiEcjtNW
Ja31p3BD1exCksCz6HR/T/y7rz6il/yJ4HYzh1krUfrvDfby9wbRlx3IcEIKvwRu
qZP8Way5M4I2VqH9WaRbXIqg+U3kOpGQ7ksCWeWgbyjYW3Rt//zmie5Qg3au5CBT
I3/2qNbRmQtL6Zs7iN9LfOn30uELmVtAnFzKQZNorJ2eINUXUy4bBR0245JS9XfN
qR4UEL+R88Ij7UWDUXgcI3WxiHg+kvdVykh99/iTWulSSwlwvDrKWuk3NOhqbCJ9
nPeQHSosNlcIllocZHcE9WsCy8mHtBDgz4CRkFMQCDSQCzFUT+Ebjj9CFvEekm/x
OEByYaRPX5fcuMovwjRWZcFooRXyE9EcQZL5sJfxPJ2nxcR6xQfOFIJGvyQWdZBi
tB6Bv/MCxw/mMV1fLEmhgaSsLE096S8FDDlumHRzLPG+l6p1ewARDAJXvrLnu3Nu
aV3zVsnMl2EJZkm3u31C2X0uhhqGAJggHq0sLNGajxfIjns0PN1tI4tvEdBRyeI5
EWZmEBgbgLZ1CdDUi24XijZ/rtmZpOvM3gQxq+iO0tGfRfSSFB7CjxZxqgG9VyGy
o/CA/ihAvrtehpKkgMOB+peHB6jKhxevglJRxfDnbVAAvudftFeF7crOuuLgkTrq
gDSSPLvyg+0JgYUFo6VcBT3zFNugJxA4xMoiV2/lAG+ahbsxRwaPMLiXcn3CXOBV
6DOyZky9Uw6Smjb99N5sD2rgmEekG1SYW2zjDiPrJ0M08Ur1vaI6tIxtaHH2mG40
oMa/DA9nE0slth0U5AhT679WQ5U43SoLqt0kOiVGFH23UCI3Bu+treQpv/F/GNKi
tGHJgIHqFsQuuTveH+UFGZb5ZQOB7NXi62Mzdevpi+AlO41C02WypaMXJ/P1gjdt
T8K1mFwkEKLVZDL3C4wheQx6Q6wLnMuRC5WJX/JP6D+t+a/0rRbPw0lQP0AbzOL/
rKCv84qiG08Hs2mH5wyhug+cfgPDlb6NP6Nm0Vv+7xtt2Lz9SxWFK+S5IhSKXEfn
0YNyWcUkYu0D0KLC05mpmOhwYNKzhqaIY6peaLtMF/pqqfEZ/Xq9epFEX0aQ0Fs3
4+1z5uU+5J/CZwUaiKNOI5kJQWlUHGHEGXezTakkHkD5LN+fDiZ5w5M+5WH6BIpa
kbK9HguW7y1SX3YXyTsnpao2qIAamLUxP3dIquvRBmIeL2NHNo7sVhPljdXFShjw
mntkUGB9Zdxe3sYb7lzs7sZlfKAYqph87rnNrCDflGPGhkIdQENyYzD8suTsl/MX
7UKec+4c88y0rBFwYnGqTpA/wBrGH+47v3ZhvPc+R5JUUH3r5wqM6edihuLGjB5e
E3/x1aQObtUbOf4+JsJKDjqzvZQyUVSHNm88xeUE1vmjA98lscYmsnscLlx52IqW
fXkFZ1r9+9ky5X6rc4k1qqMNcaB8S0A+tz8Ia6vbBW6dVaGRlQVE06T2dB4Rp2h7
qODT0yYagZuCI5cMUQkIl54E46uvGDq7A7bFVd5AIeyA9mdZp/SvnzGlSDAT5Eog
jfHtYUVTumKSVZfRRK+Uc39Ioujde0/a2bA+lX/0ONq/GoITuQClgNDcl7KZzdkI
oPLZJB0YioRFsIezTLY3dWfzPBI/IYcfdsSFvpoi+hc226eUQun6JCq2R1nki1Uu
PHwFF7BrB2E/IFNv16ctEQBg+RF19WiG05SWL8GF+Jj+rIFBmcUyXgTjbgDXh6iB
W/SHjL1JPgPs/tGBstkVm8tNKbyFx4WMV0tJF4sCKnnLxA/llN0qlRdXcUy+gvAy
hTIwFz0ZCXSrV2H5NrUvVQb0IfhFyu3PHLCCxreWQTGhgrWBLC0phe2C42I3tm8P
IpCWTijkTAMpYLdantvJhh7m4dX+NyIUvHsXASIp4V49NuyeMu2D0/JJii/8Gj7y
hj/Q+pcY58KwEc331DucLzXgUhn+i9wizIgWRVaKDw/FAsPclz8hCo46/aM/Yev/
nJJsKJqs7I48fl6OEmcHGFi7yy+rxwkHD6Zwc6UeoF6LVRd7Wt42wEMyR/t4LTX1
X4AW7Z8FcUg42E/mVwfx1jU8rew8jD6r63UWdeUYo49BMQV0H4raXfXqtqOIpeK+
qjZjjtsJ1XaknePoF0iJSxfzVQVptJgM1KmUF9qg8s11V03bbQl5EbUZjHNfEQFX
wDg4h0PQKqh8aRN7lbBWhZowADL0ySyxXTIOIQ+RrL2k3XgMIr6VduVh342UBB9Y
l+HE9rkbdiN7IaAGHothZXgcjgYziuATZiTik8EjtPwcIpEC4Jsyg89yFuqxs1fu
OhE5uIIfR53cQihBpxkPikNyNRKrm/+/1k8Obdh9u5lD5aDw6iANxY+eetzTrGAM
ge/rbtriu8dhT5yo2nDxAo9z8O1657iTR6JTL76tK+BzXU+wWakYhpqJNmkxzEQE
dnvLodl/Pbc4DfVaJHDIxPzN+WJctlc6Ef0R+HPfZ9CoQjtVIWX7ANBpUecjUiiG
m8oBbibwXIromjh/fiBu0dldMcWMsUW+4ydG+93P6S6ZZV4LUjL3uacxY7risTDw
55x5yMbAWN4m4aCeQrNaRfxobHisvQ+NERNYdhhVbrlEGem6aDoDIRD9V9TUS36e
LpI+XiAc1i78WLivIGTH4ePzn+GNNi1ZlNiHqujXfgcz8iRGvMJH3+ZSNHoTzOqL
Dq9pqL43i6QkWpmHLC+0hB2YsYcJQD0Ne/N5FLEDAObmulsGfDEIIz7qnD7d1E8C
DoLrgd0BqX7+Pc58nvncaASIdtjrwbPEVzv535fO8pcjQDu9tayqbtVG7N+59gf4
jJ2NPWyatwsvt/ZxEXBJWht14by6iBONE1V1EOPtmHJov9lXKugRzaINJuuB7jKq
He7Bv3gFP412cQse4BP0Ku8H26T+F25JkJS1NJ8KO4syjEBVdhXYFgepdfMFQoI+
ZSeTOI3nn9gvOQM8D0xXykpY/2PYKhFxQLYVhNqHfCgyN//9y7HWa9mU/Ii2SvN9
B2r8fp98sPGDDlZVsYfHof0KHHnGzd2P5tpDTy7/kSq7Jp0Qk3b+nb0RGEZIpxOk
xLqCYF85MLhNdt8OdxwDhgmj8/LS6787wN1NsltPDNcrQMpiimFcuGTwJ2IJjXTG
M5fqPYv7wlIUqmhyPGbt2v0/B0lKTfcofddUCiFuevxaxe2Bk4s4Qt9aw3Rm3K0F
i/bMvJ4x2ha1P//DMhySeuCS4z0jm5mV9mmufWhONdy+YGDn6tQLotr5fMqq0Cs+
fbKxKp0pUrjvitc41GGgvl5BjkcxEOaikZspwPtbINpN9Fr6wdTczmTJEVPChkYG
SEaliZDVzucUYRWjviNfMnsQij9fxoZ+gArnMu+QkJVsFVfj45mXrZvdbzsYGuGG
tywuSbvVpBABlmdrkOipVcq48VLIkc+XB+XiWePFf+AgIqTphFWQSRi5pg4hMeyr
N/+OZMBEZKB/pu5gx4qUK+mEk68lvf1/bNpn64rkrMc46jspwcrxvCEqeEu8A8Z0
SMRm1otbIMBCyixUQAtl6Vx/Fw3XiKwNJzTRxLPf4fg9JLfcu8VmcjBstQwZmb4N
yYxPTTZ1Il0p55UE3hPERGWjgU3XN1M+At0qIJNaCqMfOOuIfkb3K+D//Gp7QOCJ
RRpMwO4OSeeFSPuZrRxDi5zCP7gclF9utxm7PP0KE7x0qWcAI2/zCSj90jB+r0dm
DNtJeMbGpuZcpsp6sCuUQEPqGrTsFJRb5kNrPJweU8Prfhkkg2btMVrbZYorVVUD
Z4M4HwJYt4Jjq7dkcS4+XrD1PWVf2DqFBlWYNXCZo7/x58MJEbEIa4T0AIn1j3G1
FwZ6sG2o+CQYcBBdFGDt6blytJG23aQa1BnX+Lhw5dUct4b2bITRIv0NhXB9fvfN
r7D/hXgx8KOWiLA7qpaVDXJsV6PUqXy7rdFVhnykf2xUvPI56AiEGLHOKWEVJc3p
7hBMVYGAcsqH10Ban4GerYVOg/UGBXv51qutqszGJYBMCD0GSiTKMLoAKOlF9Qd8
KemYZxYmslLazXRg7xXD7IVDWOd1Df7L8674cMKve6GWePeFLOrJjXp6zVtbWz8h
aLAtH7zFRhDxOtnWwETug+6vCPDUCLfFLswN7boNGXI9rNT/wIXYdHZABr+hHv3Y
YN2satMpciHGdvStqSY1rqSk7K+oKTpoGMB7p3I3GS9RXpmxlmnfMkg3LGpw5Kh+
eWzr7ohuNHWpLAlq+wPVe/nea/OQXtbBKleR0GIQFj+oAf/H6EyiLdP9kUecfIxB
mx4OcXfNiBOMAOuVksodVWWhBQrJql4L8QwCCfMrA7XXXYu2s+QmItraWgc2ABcD
j0xRx2PUNRdYP/e710Icm+KKzRVMfQ+3QdZ/mBdGwLh7lJs6Rb6VJnDuUGMbWBEn
KY4A6Qfv/m0dz4BQUo/+3qEMSWBB/TqSMAYkyaKsLyEyhm5dVFGMuKS9k+N8ATwk
6LqxktEQORAIdvR73m1VCpsYLQmVAnvaF7L/AD9M0FruDzrpVeSK1lG/gzgfWT3O
HhLLZrmiA00gfnBUl/7DYtvVmm9P3zyIOpcTmzKWN1WbVQ+OUgXB9u8nTm7syZUI
80fJJFaeqF5KDjX+dfH74rqeeR1hPHTYQkjX5oPaRGEVKse/qArOaQftNN6pkaxW
RBy/LTG8XgnaHVRGUN13tbLsYykBdv3lNdX1//2CdazE/u38QDAB+WOUizbCefOO
566tZXKqRhKZ5dN6i8xk1FUHqSYv4qDPstnSnQSQ6Nc97V+eu56M/+uwCEi2Z+Pq
Ku4utK3xN61Thwx7YX+jGWpaUTE7gNdf65HXOcGbxvi1/E0/qkoC/B7O2uIsZ7Ny
fmmuQBLkBiTf7sIFTEf8V60wdsr/W7mV5Y95GN1OGveKSspRm/OmcmK4g1KO9OMt
+udMlcmfn6o6wPvMr8iF+T1lZa43FgPuHmOq2iBgBuBItyPhSryFwRiXHatLSdRa
6gdmWKWKbOaqkosonhsUkLPNZGRLlYgLJX5mXyubc5XNXR9CXkQDVckfeRptli5G
0EuuvHG6Mbo6cMvmMDthHL6Kl6oJCe52j55RQegQP9NuSvLy58+SHd4f+tGKL9XZ
8FGhoa+ym/or4QAryzFVCSlH8+V/JmdfJ9L/FN2ieXLPFPrClOCLl5N6uNTGf9GL
PfS/M4fpIFQ5DKz+CvzH8oWUXJ8SpiioQHdoYjw6MgqE1H6XuXxO5MeET65LqJxl
B771w0GSdh6Kt6b5kNccohEUBQ0piVGeSQmy8ni+R4ySCWPEc/3SoYsTo+d6Yk+z
JCq0iPd9JHYrx2W7J+CkiTqpeWLOmP34sLQ7TbjQQyHGBZMLXpb0KDYPp40Kcp9H
u6dH5XhDKxpKp/7UIIPWAzBxeljuUyDCxodHKQTQn/w5qj/U+OLb0vPFFk7fVIln
cOYCygxynHRZ86kgJXD3fCpR8ji0VSvECOh7MUwZJ0o047/Fo5tWGIENLhGvaXiS
6JjiKBmQkTdneI+zmBgtWXZoDttfK0ti7pPKwcSS52nNVMWSb57Ai7POQ0qDE4T2
PSM4SyADIOqjNOpF0Mbu8MtoJXO8J4yLoW4NnFA+wUeT9ea8TkSfbR83J1f2ha1x
ZitW8rcp0YEcM8qXorjRpDuD/le86et4eIYQO1BJ1f2fv+MiyOh+K/Jc78et2bOR
OPVtyFd1EZynByrywCcOleTu8cUiAcM1jj9vQlLxdr30MvdzhZrmXbiacsczRr0V
ryV3Cxm52C3wDnQhzG8KiOp2jQgQe2XwDkSI2F2VMXNhDmY8HoU8XBuC2dmSbExM
Z/pajTKkClCbKqJOAo7Oa6hpADsyJh4mdQJkCz+O62Nh0lLdLK0UpLz9ErE/1qeu
qpzV473nPEt2gj9amyMAXutLP0xigBWPVehzetmOYdIIcI/FNpINJkWKUVFI1xQk
iaCVjder59Q+8/wo6NbUFKIuhB3N+Wq0f1WgC7Ks0p0iYe3L8HAOUWnC9vAItcxE
Md6sJ6aZJEXA7viXq+XbU8MOf4u+yRI0UBZgcPvod91zm2mdqt7Db47bTFjkzoyk
hYFX6t5mlJw4ncMAt+3DjTdOvPSY5HiVT9My8f/nqo6EglrAh+OhxJGO3nTKM8Q5
dZNEVHg91e/vIKre8jQ7aKRqEytbEvCbKGZsMDyChFwM1WFtYahHb2bm3h8IcmhU
FhpSmlW0zs3cM1if0vUYkBQJpQ2KhKGHjekZgnVPs7nvsHBGPWigv20RK7nDtC34
3zZjxVCZHW4R6IZOOEEJWITH9asE7l7BkeIuwWY85RcZwrtDpGGRhGPtDe0vyQHU
Ff7RGfrSFp9UM3hSo7aI3u0Td8uHUuAe8elGkaT9BMhPW2J0kbH8WWFDMOHBQOhD
Obk8yjLKDcONhBv446bHz70QRHlowiqGlVSvsT+zCkHnKOM3zXG3mwoorApnuqdu
q8iT1uzh5KYkYyRdthMyclHuyteHQ5i9KLB1EMaQScAeG1ZijYi9s6m5Yt/ZSnXD
MJbGnuHfjTa+CGCRujfPFRZJFD/K3asqlEpEazmoXiSWKwLk8/7zgJ6ScRbSCZ+z
OFe1LxzJ+LyQH3/moqwcYogViAlhmomFaefYn8Jb8GkND1Z2V//idkxEMwcVjaac
vk9EUgmd73hrmkUtePX8GwVfJBUJ5Cmt19cpoxcmaYsDtzKVe0WaipRYnOvJSZAQ
liQd++2o4KyWhvVwOp2roEvXKD1GXq2rnNRszEIw4gJptmDjXaKTEj2F2ubOPuuf
VAzJ9N45O6vLyuTRupki98wDFz4f0CGfQPfKe5Wxn6r3BMR04vfLIpl7f8RDTBWQ
2r13LW99xg7H7F5RrumNAuFwf8nRroYy8sp9Jz2P6wSzOhiyjVNeghnB/XugTIDz
dcy8x7Tm0c3DZ4Bd7bZT2lRxhnab/ShSx6MB4AeJK1SzghJG/dztNYXW7cTPABeu
WDNEjupf8JN8fISfiWMvQN3dcIwxHjjgFF8dLCkKXHhRAOrEMpQs1nw6XVCtnr5c
U0NCYlvdBmZmL4lzbmKH3ppaiglC844BQMEU7Z/DNP4IPMW0lb1VhzvoGd/+/9LN
1DGVKpT/fnBJdKlCuwuXnuJdVUWSL3lIWjRWyfPPXTxRgPZibViySeTkrLXcJzvF
6HGMPahuMSPqksb7oDHVjVTdA1HAfDxPCcyaQv7mDBBEsmufZFIDsw6hPfCuiI/f
IBP0k4MB62eKDPb6xsbMgOUHwRNiBcfhmEAVIHeUejOOBhdzm+Z85wVWV/KvUdmK
GD9+Ecv1RgcI3xERLpuMaU2ktNb093MA4XR28JRRMZOVm3qngbJO6aUbU07/pEGb
TN+hik6pk7LkM1v9k76DwbIvBP/rwd0Q7a7FswF/ZEJN1yZx/zLhr29lJe0GBYTo
hV8xI5ttjbVwus/IHUElWmyMeF1cgvGseIFxCK9ZrD7QtEmNhj4zUgZR+4UznmQx
k1drhqlS8gzjJnkMZAvy1h11DFerW35oyjJO97Kee0uyQJ2/V7Xpg/Oz2YBfuRMY
+Hle4KFmy/1TyNhIfm5NfTUBjRq2k8ZGpoI16D6aCORKJf9wxIluIEzNCuW5z3/E
dN+qNPWSuznVIPryWnsxgDtAyIs1l6L6J5cwlzKGU1KVbSUvszNmVUkTROKtIWkR
50kzxoYjtUJ5enLcgxE2skR/jqtu0WNQX3hKqtCroX8VsmLq9b7vBL9cIW3hUsv5
PxhPSru+VMyt4R9VkE1Eu9hp0L+UFBW1TSP+LH1S57RK5UZjFTHk66aig1FD5gcJ
L1nk2PZrYyNfYYsO6TY6Dr8rTNFxFe8Cg+IvkHtjio6fdnZi9zM4ZQi2QJZZzQN/
yKC/3rpJ3O7KpfAtSHl3I7O7AYi276BIKqyGkTWoED7rECPfdm3g/Zifl4xCj5g+
ZYL4T6OieSiw1GUzZM2DtjFU5cVySsru7tm18+CidOpc3Dx98YkDcIV6TmdZIh1z
HF9eC8qYG5b5vp5NrLOnZgDG3wmY/4Grre7M4tGr3WxC3MA7gBX7skkbhVm5Jv3Q
R4i9WTXq1WivqoW8AF3NIA8ZuvOLBShRVMzjEqEfezLqaG7ymADD5bhVZCdB+i5Q
jpGuw0KAyoVOIxAHt9diupD1379iKUXAp04nwBgc8PJNyO38h+bznmKBXpolo9qE
WAlQQQXmvnm/E7HSNRt/wcFzC0aJIIPNHQx42ZBXcUlVKfsF++D23dBZiy043Mhj
S0ZpqU3KPCXt+ZDKbhPrDY9pliU+JvlUQGF1pIQ9cuiG5iDJvpUq4QUylWOoueot
SQENNz+N2KwDxQRmm23jvIlS/qnNHJ9Qumz1UcMdpe0o+P/5Ck33JWCD2sQlghwJ
9WimpsgOhvD22Qnj657u5ivKGckYdaknkJX/148GtKNoZ2UOc3rosVc9Z+fW7D2o
PQsda7IHJFpHi0HH5KAxgYb1ZPwcrWXq9gsVzxT4nIRARpkCA7XMfwJVV0QItNZp
SPrccypuKMHJSIxPs/LoghYTn+NTVZKpyo56dADpZDMoCLXG59ANBNW94UTOymLq
72QbgT+Tlw5D9Fs1ie37I7/RKbVB6nzo3U+V7Jseh/BxhIP8LChHe38xLxx6CPpE
+kaU3M3CdJdGJrBSO46ubT+J+d0/7vdwHizgthB3XGvSfyGf8C7yEfPuNALurNSo
aNGM92Cc0rEFrxfLvlSsyVP/75ef7OO1p/78rYOa3Q2t9RRyx8EvCBcyqbSrhZj9
nwI1lP9Jrl0QxA78jf4hP5CKLJ7Se8rv2wyWxxj7iM9UHcDeU7yoDmpxvZoymbuw
X39z9DKHI2R3TVGlUSQgV+qrRggXyxEtED3sAeVeJCEer6JK1W4wK9/Kz+NbJuQk
36cfZaOZNz7h6evnfT7hTND9V5oWgxSUwqReHmWjAu+lIJZ+Z7Lv8elsh7zY+o6J
q2wPNjB34/+RSU/sokyTIAPnNNl68QdvLHIannH0k+kmCu6iRQXgaeLtqHiAXQxy
en6jrHwWUdG9KdtDoGjesNuuNqHqEWNp+1ZdBzJh7NCAYiF0TnpwHXNhCS+ZpU5P
YYQt34oRE7dS9b7EkUBw6WKMz5XaRJICRMITcHy/YewRwbi+Bptvgwwktx/ahOMv
lrIgQTCxrpJemIay11our6sSOitynD/DdR+ovbCoOg8Q2a44wFmyNNGlxZM97eeE
nW7KMJpb/0YRRPor4QfenkeqS/iKZKBd17t8q8c/YOa17RR9ABd1QK/JAk1L9wie
8rYRDrELHdpjpBjZbBgsahC32kqK7K45Eate1pkk9SsN4KlCgWcCQpa7hIivRExU
jS2/f99HBADpN+gBHARfd4Op4rcq7/szzZz+57zopmcddFU1meHtFDfDuqRv1334
hcmYlnxgUvljj/yq/fJuL2I5Hf6WWLSWC7ShkVCiYpIhnOSx+xl4/vhtcmxEhCct
YN3UkLp3B6T2K/9NdSaQj40T3P44IBrO7YGwAJxCSrBvHux9FNP7l+vNJMknuguV
xsJqRdH/06kTepEOkuH5jB5i0YGa+j3EooVsLmtBXI5ditZVjUD7akUmiQsdFHzW
+5plT/Dy0j8Gfnrp55/LOgWE3rag//QcqYvOj4wk2Nn/lzuhxJcjSY5zQ+qed8y7
XARAX+tqOySpiZez6CCC/WAMzDTA1csvdHCyu9qt/OenUwcqIkaNX3/wT3iOBs8N
0+zVEBMkq668u22KxIrIChREYF2V1p2LTESS23WN5UQL2jpYwCiEz7liVl3a2mFP
x1cyRP46MR2OCW+jhNtE7Pl4Ukg8d2NHnH/MZNQMmtuBu2mbFZ5qT5GSdO5kDJ0f
5PuGMz28VqSjqfrvPAB3a3jS3ANLbL9VqvbvgD9W/ABajg6aOrMvOpyav9+aAgUO
9RWtERH0q12JcXZvPWaOq7CJu6bapRwjRsGtjE2jHn8HlG+Gi18vedPpviA4Jegn
w2MvWAGXbDhYcRYipGFbbUtiMdoRCPne61xEIdFqaqDVBmfeiBJXD6lLFrTo5Z4X
Qfyc1AW70FMZaSNahIIJ4MJikxbGIC1M6GMgY2gZFj/Tq/swSOirE62HXHr00yLr
S6IBfm1Nod3MY8cHQYmnOpmhMeWhCcglELQhGxoRrZn/XqFrihpuYFqO6NCrU5dn
9dBdfcVGNNHu5uWySDfxuiOGPHRU9P3D4fKQQI3tLYX1cojCtwlwETHMwQDfxvuG
gJ7SLdVo4qngXYvibx69i8fJ3lvWB0l/aX1y1boC90jt0tn1RmGHypjkbzDb2YxJ
A/ddp+c9Bcw2jgolSkaaYG0Yj7+2DQaA8y5GGYTauXezNj9Cw+MQidAldp8CON6I
If20pW+2Wicep/yP4jfo9lYHg0bZV2m7wXjLtd83c1WG/6bN9uovHQ/4MubIy8Hk
lWYf0/9XwphxNBjwdIZPkfD8atvfO4WVlWfwMO5641ieWP7vE8hXVsOj79VuCHOJ
5cDL1Dg+IKe5iglnyfl4H82RWqJjaTPS/P4YERcTTlXWyN3qA1uHH9XW4oQdp9bF
gOQ1upb7hnhlVYypYQ4knpB3Taw/OX3UmLdiTWKe1AVJxPlhBD3IYIWvB9G8NW2i
0kwRW/GEhqzGrWO2CXVMBWP0wAdko0wpCO/1eh3DHXV4hb+8wgIMc/7O4+JM8Zob
6Le+GHKfMR9csaGTiyMT9Ss0LzQ8D5W0sKTpWkpDZvYAKo4YwpkA7dRBcXh4kn+W
lRBNfmAriRhkFQ7bjbErwE+g+eudt2SM2fRoSCC/S/onob/ewrCPbbfN+blRj159
LiGpirvZNbYclDbGdfQLaV3utFCQ8aQpLXWoWPyNntv5E08MIMIZz1Ow/Oqwuj+2
AMC+DJaAu7XF8ay0hmbozsSClyMTxNPS74r0Jhw717FWP8lraUVOKvB72WT8hHvs
mhIJfImO0UaJENMOry+TBsXSZ4FbjLu6c6ifuZ1qrS1P5dNIHfMREL+UKyr1CCf5
tbIhsi437z2DSXBKQniep7cgvakO23paIW4xlohRt3JwxHZar+TpxWKF3dl7mZKp
NixJyeQ3917XGT6Qge4YKCnptXljRJJk6aRhJj7i4gALBuji99g/XW5YkyKeyZd7
lJnTRLSHv1b0jCSaTyXweTOW8CXpuB+E27935Fr2q4UT46Aednqa4z3+DDBuDWeW
Kw33zWUn/NxmN/8lgXhCqXF1yKKAMTd3eaFGJbc27FJsyP8XHSMt7vonUj9/r/Vh
MWO/atlPQba1Po04pZ9AahUaASYLzvM1eaSLI6Tn6wAz6THALY0FzjYf8uNWLhSl
UzdYmOaJ2Box0S77rVfMDcKG1SoRDMlkWc4RvoHBM9qdjZTIM2akdA0pGbaRS+d7
77TfmYNb+b1tifL49RGQibl679KcPKY1wMoggjDd4Z+8ekRI32VTMnDokP8Hq61R
q5sv1HZcHLrKnuTWWEyE7xUzomNKeWdh3bibzFNslRqnlds2W7DjM6WQkjU9B+89
a/XWA9/lcOSt9+T2MzhREAPIFQgQvsccID29C8YyLWQ99SRqOgSzFDOGpTKDtTG3
+ab0E92FARdfB4VnBJum6jMmjuQ/ohKd3yuGV5cy/DDeyq1Vmr4wg2nWz9Ub3YWh
Z/vpMx4fQlYloMYcnYZZnC88Qzvbh9AJY/g4c7/iS8gEGNNk1KkXYShJg9+/ol/o
h/wqKPHm3gN+/iHYxXLH1FMw2fLdt/yFXOqNP4ZEe4kuY4O48nwIxt0Cm87Z0a90
tJWOlUNHqoHKnD1ef7+ZnDigrYhNaNiKFFI2rkVpo9hVtWEIsAKHFOxkKlMPMuF4
0W5jHXpVbuHFkfmxEZjMTptpSGGsbqrkJD/pNs3cAr0Ur+6yPLzdLhe7pT90LZ9M
wYHg+XrM8VR29t+nCBQnxZZ851D9G9zqLulTa74KreDThlAtLpRG2Gb42H4oqfvV
dKyf4NFVBX4txP9r0nEKGvwUXTArq2nCSvCrHT9ldhGOU3PVsjiShaAQkBcYwKMZ
XUo+S4JZVu/VORHIlfEqsOg2aTPue2Scy+1EIOHcN3m8IwkWN+yZZba5sJPcZhSu
hqtysgOCVCVu+WOFUXcnN1p3rO9KoYBEuxTQtLAUYNyBVCWP5JmyoJamJhGaxze1
5J19ShZr6b8YI1T18bo/7irsCUdSihGrmcTSFoD3MmaxOLNJZPJvWjhaxm35qgL6
LHBwcriw8OoOJ0kcKbWJs/wgOjsp0QtJvKd/G4VHYsjLJdFfZE9IfxJ1N5m3ehTY
jBhTr8gvmTvLEgFbly5wsaYC2SQ23NQLqYRyDT0tdSvzsQLTYJ0HV5lIzum3tEBs
tbL5YjwFLleCghs2KHLr5o9n7ZdeHbKXtpw8+FG3slmXdQnNoZ2YZEujKf9jNr/l
GJEoqeL5241bn4Pt9xW9BuMlFFGkr2bFUYtnCI2vTF1xhQFpi8RqKHZHCAGfzAJK
I0UbplMAYtmVD5YNkACoAEBEe+3nCfNfSN6NsRONXuRTz+tN261ulEXsEsx1t4L3
cNRGoBCQ1/oBjNsVGRdG8WGM9qWYU/wVDkMX8lHljD1k1yBm1TWPLZd2lx4gIGnX
YxpDrTlURXjojwLL1ZM2iNj417RH+ABwMVt4SrsGRIoEg5kVjo4B+F/xue35zy2K
1t8zMY1buF1HUUmwEMyHqFB2O6VMDxpDgOIl+XJMe6B/RzWCnOrUv58lQlAUpZ5h
G6rwvI0/Ls4WRJ4ucRI+3siDwJV7AjcJ3LQYCATDYpVINX2si9GZA0m9whygtldF
oWlbupleoZQUdzKF26A5R1a7Ick+15yavDkYeGu0ybpfUbPknHbes30nZ+84eJeQ
V0jmE85sZelfgLry1QtTGi/jdJZJePHg54sm1Mkd4DtPHqSaDXq+w4KeMbDF3U9L
soVc2a9IQ6jDCU13HvPUQvfGTAyUgJxzpME1j+RU4+decASC/3RT4NcRhIkGWxTE
tdHDofrk9SQPNCabEZ8HB5LUXSFpKTtrSPDRFTwliSzif19FlZquJporA98Ma19q
EOAH5aNAQr9ARU2RQO+Fj2W9+xPgoJ3pJ9Yd/41i6yGgmZvwsucgTiBIyRe4KE5Q
l4LbZdyPzqdk4RKu+ufHTKmKGKhrfnqf8OfJxyQErg2lmdWdLWa5kcJRZrnuMReh
7FJwDwDGXootqyb3DCwgk/roYso3Xlcc+bMrSFE6HGmOCv/kyW8Ut9wxR/OfkzWz
HqkWF7UIkDFiBvujaXVOCNU4C7MXs80mpIw3hAf+Olp+R0EEd8Ag9Ir5WVe9dvT+
tn21JsF8SC+H6Pz4sV6zREbgWBMTKN+7gwa5/knh1KVY36J1js+CiXjbMHB0yx2W
ohGRpbRtpeYsUWLK4M+0+b4d77iceUgQBwTDDjhAEtnCeJ6D5DsqNuuxaX1VSgPy
pr45wuUPZ2CiBbDfWtaRALXG0+nacO+XibrwJlPoO2F9Oamu8rG1gvBIUyPH2wQ0
/n5Yd7f3Lk8RgsV7IRf+cf7pGIkdCVDMestPtrLodWCzLR6jQGYdR67eCx8N4xfi
+I8rXI/kdHngRYS1uDkpFob+97/0wOmQesaj8EvdLrBg6C841XbIu5nfFr+cEmsq
u44S+oCSzM37wPRWpexYIhUWqkwY21sWXq0qaBTrnNVyc2HqHRUIrzEqA5vcVkEu
QhD6eRgvP2XCKILrNOjZfHcz/C2WoEATdyRmuvVJqD6Bh0516at95OtYs+y0zzIy
ke7WE++YXZRJRcg/Bza48UrTWcqrflSLWXL6nrdNZOCYnq4d2SOOQ24BF1dHjP0O
jKbQvCJiFMm+KDwFP6LPL1EuXRho8Eykb9qVccu/CC3klonLEj6ln89tPWcPWFuo
3X3WK31VQHgtY4qBX7jeXQm4UdRyMPqiLRL9Kge5ls8EInFnA2rYlYGifwqkfISl
5eOUaMIpCD97a2IB5lZPS1GiqV3PJItNx/qOzZU5sSWtHLDwpMqptNfl1AvBwC0Y
Qz4ZDL35irr+6ivgJpjjN7c5+tUn/kGaqaR+p10S2VqAvMwutkIu9+vI94MtnDqE
8fDXEYzjNp+EuQcFRSu68ow/xnQdvGW9OBISOT7C4Gd8t36l5k9L3aTEpmf8ciMa
6hbXyt11vAn2SKw4Rvw21R5uF63qwQ7bbwjE1GTc9OLK1Bq3P8Mp+Yr0D6iNSq6b
Z9lrG2NYjmXjQof1r2ZGyLubtsmlvVUSxsZ+ZBFLvNBnlpOcuJYLb9gM2VXsG4Ba
bZCXgJJNBhEJnhdRt9vbXZgH70c6ihzGO916heiiB9H+hQC9ilI0zwEgDXizZtYT
Vyz763cWmcWXOKHfr2yCcftWmeV488U1av4Tfm9VLlaY8RY9YZDNF8afnXsEbGR4
OQ+tOonM4d5PlKKTVAuSHb8RZX8J6fdBZKZFeDGsvLc50nfqsBdQw/cy+ZyvVxGq
zAc59o2DfQoyYaGsaUs3R+6Yr9tCAKrLoKpd91znN9IUP+CkN+4Oorrxq/vEoDt7
Njgx9aWEzLuzk00rvphc4jrcf4X/5/cOY81mVd2lYQJcdrwqil4N50jM8QsCpROt
pdeu0pHmJmC4YTXWRf58pISK32BpNXfKiD+n410jLwaDWzJzbGiN0tWCOincJZoA
tpjjqHMilWhUtxbvlko5yG/YZ3xtQ0ICdIv+I78phHQg3vikjMnzCPG/3KnNTeHK
UOcxCaLPi+3TtLs3+s2NRH9PLXckdmb7Vqcnfh+DOUdzpOzT5Ajj1D1H6hQ0xTte
iJDn4ZqLb+q0eoCT5zyWtZtZ62+AbZRSibWOPN93R8Jy7KoV2VmSoDB6afkg+dDY
VqkVZbwfy52KXMIoGE09qKrke31vkhtMAcDbuJzT9Tdek8DlpNpx3lKXQA+PddRY
g+KGCYzAs5E0XyE2ZGagVIRQfQUp0EawQsu30KjIvsMZE107PL/qHvcqn39fIoMf
qWnXqttIOexwaVNVpiqlmCCO4eSCRrUjTqbaAU50Y2l04LzIt4dWOC6R+cAe34oJ
ISogmbj8b49w3qBYNHp9rb3mrXu1yGCnAvPx8jaLjnCW8/nxmdoTW0dIiYl4NNuc
TGcqKuARxC4eamZDq6bKh3WqRAaB24nf2kpGs36qZnkb3iKISv4rfRd9GAvjFx4d
HZTocOGgPde2xpsleUYe8w0d+jifL9N1WBen6mrrsWVbpAL+RiBwj7mSnEBGuRQA
nLjkoGRjTXRGQdPg6fMdS/zgasJ2Mggo+PX5rToTdn9CouevjobTp++a4rO0tVXW
1nBCIVqtNS0r5YfERE0om3ag/D67VDsqiSa2yUfaOdUqpKQyu3QsOCr72YBSdTQe
aOUc3hMngtSajVuvErQetOhpaoxwWGb2pRvEEcGIpleR6iwgWxQ0v8fxpc1EIEaQ
LGW6scqucl1O81NZoXJGD/Epq5+YXbj+6PMa5NBlQMcQfIazeK+2BV3S371Zzxqo
sbYpqlwUTQaof0tZ8tOIql8RKy/kbW/KPTcpmCos2wUeRfKWuWA8re8G/fBqfAwy
KfD5jtLemSM6E6LSOKXr+dT3KBj3Qe1q++2d2JqS7zUAmUhrvNMlsP1NjQJLN2p5
fIvnjxp1q4oY6B1zfN8i2qXCGyX5dzHYWcfxWiTr++YCOmV4kzSzf+IOPa647pai
+nRKv9bNJho26YK06AH/456W+yR2AdYIoY+YA/drLI/q81jr06p1oN5Uc7V38zGR
9AuuW7J5c2TUS9/nYtevlvNipk54PE1mTn1urB6/4VyXOQgOrnHk3dN0ZwQuOpM+
IEQKvf8dqtOZlsip/Wch+M8VGCymCZHaGzEKGvxUgMtbgMPWn6NXzGeWOdJZazqx
SC8/qlIzLE94CplbtV/WgY035abTludDDi3yJSO6Z3qZLrK+MwMrIFlXaz8iV4MD
pQ0MlnS4uDPgjxgYwpuLN6BJhIyF7wwhCskOHdlRhdMh7YeGV+Zgo4P8GzReca9+
b/gBRB+Bm6j4+LPLSDeEbmnMfiwVHNu8PZY7iEYoz57BxTba47c9lSUbDvkq17xH
6SSWfuUxGKGMw4CYEzm4UaUdehLxxYKWQ0QbpVm3sVx/4P0k916gKZ5p8uzS8VOL
/8K0LmcLJQKPdwmXewIhyKcYkRjg+CgLyI5MGfsuicqjD6njeO+Crl4qwosdcdnk
vH5nu5EhJB8FOwmN5cLq0ByJYqZJ8I0+0uDSxexzORu7+nQeDkL5ecD4EXaRJqak
+ZciSeXbx8nMVKs1/xpT2Q2Qiuk+eioqlx7Wicy9Xpm1TIZJ+qob/xmaOr/cEMaC
aEYhvinBV5XuSh9J3oCBmM2xy08ycmHmaGZkYgfJ77LpVjTcd3iixz3MqJTuvLlp
01st/GP9+Lr/NX6F45OuKSXICToGu43pTkJ6YSplRx8U+Kpz3sGZDutpcyWEOOkE
1mht91qlHMMbWXqc4yl1zDMI8hKEF848V6NNElrXKvYmv0ckQL/IFs6ylAvTsHVb
IzLmPIn5E0uu+WuKYWVzb8AN8e9DRzDf1IOpv2xNkZk/1x0kE8KcB9yDf68AnurF
NhwGfgNisQioYH/WI+RAZgerLarb6sXBaFyppbYFA+AUMj9dCIsY7GPAp9kPUmy/
ZQvU9vVXuUfAglhjHqJTReoQHx4HGLyOvweo76IJkRzU8ifx2QBzCJtiPBS8zU5q
PsBnUXJQ5Uew68PsGVb/yY1yVA3jaJiXBGREmZur/4tgtYYZk6FIrWqIq2xBXap7
pvPuHGeZc5fi8ATT4nP6zYTvoVRnpb7j+jVwB3r80IszYY7F8P2uXc25t1TNncM9
Cl5VV4SesRwitiMzqxWTMfd8BsahLyVd5LsaPRgKt+Q6svfanRzNK2CYu+JMbeCP
lvAeCCHKgGxvPm/yq/z4yMUWhM3fv4qcEUm60VFV5/UAyLisg60dOwTS0tPS3WfU
8KHRHvWQ4+w1Llo1y023GVSQiRI/+q6Yma2eqz5LvbOOfnbX+Z08i9+fMcIQJQ+3
6GAb09A+5mkRsJx9zXvt2Etq4FNFfmeI3MCfxnd6SkcyFUSvNgYVll1b3bQgwPDC
o3s2J9cQP9xZbm28agpqglW23rnkWtN7cdsso6XGWFm6/Z728XhZ4KtYLe9J8vcQ
EcbEKEDKU/hNDHX0nhJvNje7JWHmWaaierBOoSGQnfd7YuPSd7D1zUq300MKjPRW
w3eqlmGP26RlQX9cqEXmkwuBlE1T/ilo5i/Myl7lyUDpXbCNJlHMrMlK+A/1qJki
95HZanwJs88kg7JDxKp4wr9L2rOcuBJOMuJUAco1GT+j0bkouPUS+RV30sM9Q+f6
FsVAsAGd1OeAmjUgE5rUszf6agzv5rgEea/a/qYWHO/4eDS+JvvnJ0XJHz4x5dq2
x3obSLVws0hOLswPoT8uBDdf2355Btty67P+zcIcrhE3ibSs4Ls04Al2rXNT46V9
FVCBvjrcV3R65C8b3NL1QG0Vzy1dh2mx02lN1HAqRD75sA0cZ7IH3zodfFR7lBfG
sncA28kynBbcPAU1ekGwbYOdIlCDKf3K7fYzRG/2inPZ/JOLd5bOa9GsmH67fE5D
4EUzP+rc0IX3r35j5R2/MzcBhhf5teHZgqLrLxTA6EjMCukKifCJMjdAVO3NLLVR
u14bsCqAlDhdhoEMEME6YSWds3dR02Ms3MoynDkTLKQhSZzWtcf9Dv3BIpfDWkGo
gcgguVmP4OikNt6r94LFjx3oUbDsQ7P899Szl7Y2FAioQmbkY0zd8BMmryjGLF3A
mqwOaK0kNqty3O82QBO7leGbT+W1aPueOHIDKbCMiKkLYAF13sksADSvqcBqADAK
W6JgJfclpGryWjO8w14FybUHyvlnF8uKuM8VLT+FeSy1s0Z0vAGO+pqaRwbnCVND
K6g3hSkU4gd2285P+cqgOiQkqk0G7J/f657LieYqjIwRWc+JmPvatrheWE8GY1vi
M376xnbOsSYvFUjUCDsszzbETvEuz9IMWWAcHXKhqk02ZRkEEMtMZy+LbnO4kL2T
66jnbV4diAX1pgLQzItaRWK1CqdrExVuHwfiWFYkGL1zyscrlGZSgAYP4xYBm3jg
jGbIuLeSafWFUyizJ1Octy9yAEEfQ9a0PeTtSexonXAaQ5Fg0DZprLYG0xlyU7Ns
NzXhFzwZAIlZ5L8bR9oQLy+maPiqM44OzLSJ2j9XD9is3618Wvdz+0ee8HPtDA+0
23qiIQpTqQRl4JNesofV5BHzMsbCT80H9lOnWMjxy942H7qLYuBp60W+HAhccBEF
THdALgezqGi0ZYoXZLcxKq3mDMLFWcf4w5xTn2+DO5LgNkyawSPZ1HaVPt7AkzIX
k5thPAy1ycNAF0AqddJUrhRwCLE4bcNOcKOa4M0+sYbqAXBD9sTE7i+OQ2Qd/JNu
FsCYWIIEPASs4zlft4OQYt/xqzXdHP+AE8akLtnhhdnr9KoZPe0yOGMVQpaPmqCF
jyubqeJZhrG7Zy6QzCHnNIgAwiuBUE+dX2pKi7W11D8pdRR6VRz0cjS8zv3EslRT
Cw0o3Bi8jZCYfwLB4x5TgFatEMvZx45igiytIL6iO1cDo0VUscI4XxSEfNNFBrum
BGUSIx3QjS3gqcIK++xkLb94MLazW6ihM9FBKTa4JRNDdjfkQs7CVHGbmEP3rvJq
XcrgX+O2tGh4N444K0wu3vRizUWAlcOtuDtLpxPtxMeZkNrklEn3Kjh3lcRmYoCm
tfveY1KKK3/pPMy1vbyBVS491BWkN0QodMms2WA2m4nmnPkt1oLaj3VlLriD/nrT
vIdKG0Dktxj1C2pic2KT3/P6pi+4zcHIYd7ANuTiZJ7yTLowlqgpwmcffY026Ywv
IAvDWPyxrFeOa3fohoW769xnMmbQ5/jKdK9LY8UeZe7eReAzSBbsBS/f6Vulld1V
HYW5a0SGmpzwtlnu1QKu+wwKpY+lMoGNpqZRiFDWQJVOyQ5kGv2qTWxfV2kCb5YO
OOKDEiWHKFHvav4LrxLYd2tOFxadIQhKhCONDwcOoDIShKBo3KTV/8r10TPjacPt
yTfPRVXtA62z1mmym2S2J22b7UdHr+34zX8kEf2sKDHE4luPMKJ3J4y0Go4e1BLl
E3iaBoTa+QgndAnqGgU+qF9oPlEFdyany2POVaG+54G1J4tTU6bv6qzd91L42fIa
FnSjaJuqGB39S2zFy21/DGsDO6Duib6b6bumUEe5EaT2sDYyTCjX9YdRsN+TETuY
ZQIGQEl6vpxcLyloSBx0V6UltpxstBnz3jeO+jbXEaRtFlJPjcy+Zty7wKnLg0S/
npQuzgRxvYNcmuNxhvVuuU0ZWj5HLxLHZwLxkU8m1/kCgcbddL101tYP8Ik+HPPi
0S9pR3IIgF/oGq5BEvRAq/1+4GoGIVtlluNDbtHxuzdnlzT1wb00NLevc1xD6IA4
5zbDFa/qodRuTlwRQWr6QHGRSUHE75/44LISD6UDxpsj+hcpelypDVqpIWQQ4ZeA
1ssCUaAQ2/mFb58gRjpUT9/bqC9pltdpZeuWvc6kPAWzFb2iSxfror95k8zYiq2y
SNgo6NgDIDeEVZW71jnNywZ/ClGBtf6mAyrKwg4GlkquoWVWiUvgj3YlWkfUV0NW
W35rO+22wxDlq0U2oSuAcpzx6egAWenqYXp8rxvyo7D3A9I+JUsYzf+kc3bovZD/
lvbV8zi+EEsI07+4JIXCLzP2P6Ks4m2jyvwTjFKSsH67AV+UeztG4zLLXnuk62uH
phVUiCbN3Ft7Oj6lZ/1jHoxEpclGkOVmq23y7mCTnUqbj9g3gx+gAQmvTh/DVF5w
y6My2FloSXmMEkhUMF17AFmnc2OIEdFLj6zgB6NLFFKkpoLj6yMCFt0GpRvqJ+Zl
I+VH17360s9d0u6WFoqPOQcVWtcL+ymfq0Hqqx/xKkWF86HLpAMoxax3sG8J+K/O
0FCDxYhQ+o2EJULTZ3qT2xncWR6sFYc4yCS2oj6nMph4Q/6wbhyadNDXSmUN5aR3
OTzjzS/o472qcu4TFXq6a0X4g9datqCAyO4HaldhVPnQwDIgptllFmT31YLTzS5C
/WjzMM+tcHapRfjUR2u1zK8i7zchwskwa/ialEGAZNA7mOA3DDxk6H8p8adZ9kME
D65gFhfFVKZQSgr1U4pofEl9p72zBafUJZ8VKvLsmc+3FJCxA/7DwHCdkpSr6usv
abOvcukgN1fFhgTrcOvhhHZ9/APOPk0/pd3dDCkv4A2wtWrrOfBydyp2c6r83DgG
dwKFMGc546spI3ahszYu+cMc8Ch23398PU5mAGjQ5Z0rzvAu5Qy4EegL85fzYwRz
IpgZ1AlO1MN4lK2S3DXnvkM6EOT34HqI2d76QbHVBznbREc/EaJa5J2z9y5/Ijzi
rGjIX+E68YL1ZgdHgVJx24OkoFWgKnQsWD1q6OPrBHbWHmQDHAW4h/ZHM1xIDx5Z
bDlaXwBxWpF8fZQyFGmjeN/Nt2QnhoFRrHGMpSH23ua23+5wgA4YYrQ7sMzUtIqm
SgrSD5yNjl6EHw6l9MXQsMAPxVt4exWbArLwGbpYYhjn4GuP1VtJT65D+9uYJKj0
ms0wU/+p4korxVZdjOzRuDOfIifcKuyOhLB3RREagjRHNa/mkOaLtDJzPIazL9SA
QjJ9jJqKt0omtMhySJQkBkzdOtt4WIA4noPstpCnOTSfNciS0cHKvUiWfqNSOJ7l
Tegn3RIqgNC6GyHWKQKtTp4s1DXJB4naOyHbrOmTF2j6UmbRpUOrNL7XNe/gQEbT
S5TnivSLNQTBM0Ys4/0+sBpUpk/BCxF5K3SsH0eRP/Epy/P/YCz5Ogp1tIWAAJsp
gBt2XQlgTVLRdW1cgpEEkqdgXjrzOrFp1dfL3GmAfWpUKuTfAQv5r4rPCn/Sbwwx
XMRcdb0qdIqpgGV5vCV0wWvj6RyiuFW39AOyyWGte1ggsZn7jqSr1hGt/sQniRfW
SGja8xGWmfFwOQyN843KbSAhhJC5ACX8+0FioTmbqQwDmoRcd+j+cmP6dq2Ez0G6
d/+Ven1MfOo4jKBEjsuaRHqT+tj3K/Q0NSQqy62Rx15NdtBWi/u5ISl186X/YmtJ
yuH+0kexVir+n06zBX3q2ncRwXQ6ExwnHKw682QvBAEGyDKLeCDlgRJNgz1TQXS7
3L6Smmw54ZnV2tgPXP3iW4/WAMpIvdVHoQn8LTm4Ukgc8oEbvBkyLwxhw1VKnoWo
Lbd/aA3Q+lSQNF17Bt98apKuKy95/IVuzOwjty/rsaKrRsY86YCUOS+BYQ6PrjFo
NA8FyGVVSYzwawcnFZKsIW8Y+SUxALxKePjOvvDEKNF7tyKCTzVwtK7cr3AjZIXD
o25+4YrHStgEJ/f3x49J5QGMYdQ+mfBiN8Z/7ZYGanjC08lRy1EApuFUrQEBwnuE
EfdyBG1tkTXlpekWKhHNV4X35iIWLy09u0RhkCOtZiFBLBvGottl7J7jk08ByVle
MORWwfbZ6Gos7gOhfPgBaZkR8bJoFXwO3c3k4bY9BOr35WoPNtKC7AncEYdDWxMG
AIQDMjozmri2x+PsTQ+PoISMpTzkIXYmoeXS6+xeKF2LYCcBSrVCBJMJYDMP5NBj
N4Z+5Rbvd6Pqz/Ea6HSNaKCUAGZ/0PHgK/xaU5vMHCbEX+4c7V+zTz6gP34kvNPT
k/eQaIaIDCe/TGv0om0nUeA1jL0IiGM/JvAJUcutrBSG5YdWKPP0bOc0t8KlWQQT
HK5x0/y4pX6yayaAm5aG5ncCqLRLFAlzKvEq1gwkF/auEmcm3Iwuf6krjGgr1X2i
ch6uH+I6c2+m/YCGXAwdruNY8EbiLv1Bh5ATYdo9n/s9IuGZoPcZnnVCoYqjgpx9
0BxZYO7BEJe7BVTDAvWbvwSMsE4o795h+vz3UH1OjAmintQwftvJtNUbQCVkUOFU
bsg7uQYgej+OR4mMMUHfS5WtPwHE+7bHxXSbNTUimYivAuFoaKYTUZe8+nqg6A8q
zBtE4yeQ4bMUFh0uxX4eq5nLSzQipBvJaBB5cFgVknaoE2XyEcBLv0j7LbfB1rJi
KaR2eITr6se5TG1wRR1jQgipX2vUTKIiHugRRGfpHFYn8Clg8S7lAzGKLdQWmW2H
iacc76cnGj0tAjWhZ3da4ZXjY23zczsjsYfi60bcwfdiOl03IC9555yE6f1NdTDw
Zoo5WvPPj3l35MvJnHTHTWTpLwxRpCrlVi51/eYrfu/hEng3zuD7KILhZck4tBJC
MXMIaYHtiFZjnAqe+hNSXUdxgJuvmYCc+soxFqE0Njag4hzlfmjnYH7QU4yrHJ8k
iMi9N8BBzSBlyq63MAzI4i05TTTWa71RpWWK6r6UpfJwAX1L2Y1UFaeXfC3QkMoV
Cn1y2YbcsJesxKdcdH2+ObbbX/ZC2JckbVsy9CQj+gFkPTFZdZ0/SaRVdYxdC//i
MK6PISANT+PVWGzEehhxT13Fp4qSDB2qKmLDTs9xvKA62NIfyJR8a5B2ysiSE/nO
3ZF4yKQXdQXf8nS7qjgz1QoaibtHsUmGR8Vf6+omLp4Tk2EOZkdCipw4Bt8/qAen
aZVq4TmKp6qAjYhcJ1Ac49yNw3umidYfpgV6NMI7Pp/QouRrH6YMyoUmD2MrxZws
ZJRiz3XxQXKkDTYSYBENK41gkZ9URF1rNOHVv2wBlqMXpv8oj02cChvhm0HH3RoH
+gPhnXw/wahzXate2X4kQJcI9RYF0RbjsqcGV6ZUugwtK7hNyxSv082Tlj/mGD3p
fgQIyLatr/1GwqMzSiygpNf21wohHJ7/Opu2rJT69Kt4Oqt0FKn+B3XgrUsRIAQ5
xvslLey8MRk+w6UQt57NeBHi8NmiksTlwhoDwycCBGZcVVdmcMZCulSb1n3C+qvi
UbLSrkMTsvLmE/TqNfHVEUKN2wepwBa17GJTtK5eerpE4JnEH3cgJoZrPbtAuLgY
hpLAxSZy1QxOJt81k+HYQhLmWdz3d7K1qHSxWMPNbpYDewo2HCM7PcgbJgypMYfc
ZDIoQts2+8mAjL9HaKP+ehrCmX21GmbXpAxvx+5CPcy0PYNb8vQWyOYx6NYdy+M8
PXZrrhMBiir+zVp4J5e1wBUvhjOf7kGWiFbATtWYHOnc/pbvLbw+tgY5QoxkQ8lc
Iu6qEZku5x9qQD0fUtuKM93R7Zfkt2mOt2+egAfA51KTKsDR3mUie1Tcd8Dlycqz
tZzKiYk878Gm+DRF5ar3PiQtg0lfLm7mvPmseP9BPUgmpYkWpJ9qz06iPaNi46Jf
7ZwTCvFjeTSTKpjrCRM5iwwAwu4hRNTEwi7cfcY+9QHaM/Pp1nrt5ZN32hLMVXwN
bpF9bTekUq1HixOHM4cZeXSJYtp+kO/Zam23tF/ddTntSKTv7sIkpu82Z6AkWSqc
v/Z+XVerdoJJQMxzTGXTdXl9Ehv0pLcdg9QwDYhzZtunJC2RMeah+GZuTnIvIeiQ
qIugEUTSpu2BTF7dGML84NUVdLeFejv7RXnYyXFsIPCBn4gVDCtXW2c0VyhbwY4B
edNSnvLHVSdQodi/qbuiYzO+1YSKYqfxJNl0FpGpawI6aJNSGlMzJ7Bxmc25951S
q/YTB8HZ0TlwZ/0gnvxYPGNSOphHUfdj7FCrvw4FRqkIGPjdhmqhlR4Oh/Uz7H4h
9/MdXM/KLhrb4OQJm2Dt5NgZ1FxhvILAv46cBFhaCTs3bprmb7Ce5Gi10hoFe1V+
8IVHkFHOkl8fBqkbyyfapAMCfAtUTOdanE3zOGL3FIuGCMa1wJ7kIr+GMo5/0u2r
zBM/2+SM08pVAWIH/ygdE+Tz3py60aLuDE6jLhH3HZWxyEQxPqYvAHuw6KD00E7H
Zx2FWQGisWe9PXd4xfhLwg5HY+TngSSYb+qJvudQ6metffTttV86RYYZyrwURYe8
nC3cEyA9sgLLVaRdhJBx/D5Lp+Zd7IKJSUsRJeow2s69ooWbK9qSBxQgG6V/wbv/
T+mANscDfO/1foalHdt9xfcZvv+ri6c9Dg4TCzklCKZXbLMNd/rby8ra0NgGSBAx
V6dJgsqIWdBHIcY4DpcOKW8TOzVTBXdDQZWOOlMxv6Kdvlt4YjJK026Axe77MIGw
3Fx8skblOKTMLaevZXdM3IQK6dBzRc4LGPC8Pa/jQ7CzN+Z8RvqAHCZNe6L4B15g
VP0wZx5iB26uNFfrBABJsZuAXBdBDsF1/Da51kvtYbjFvHFHloga6eTpHm5cYcmu
50a2bZosYv29WHr5niRHaCc0rM2i0hoRJq8642kp/zYQA2qht3Pj+GodsrGKZyUs
XB3QBmuUfKwMh+RUY0Fne9WR3ZA7SjQRvLKRTmFE8ZwQ/fi+rpEQYPqYZC9FpOoY
E10nf+8b2dmVd6Uqs11oRN12LkkbWz92vn/TDxqWUT7P5CycHq45IjdOCnLyljcP
ygAgsDjyye9zXJFyR0LzwJVrEcsNqHRCF/ZzJnGNVuRpvXChdjI9+aTgUwNcxcaE
IYVJE6N+bWZaApVZ/ccciwU9CaR6CgqSX+RVv8BXDclxy4C9sXxPCHiqTh7fXAOV
3ivwjpaMezeZWmBGuph6jFEcFSjtbmnrWE39slEPe4gIZc9XD1DkmjeJMhH+IPcF
Grv13LkREiSeXXdM7RHD2IRyv++KKUgyj21KE81COTID+OtumLC7NwKblh61l+Rb
5xDwbz5uaFl6HvEWeKa2mbUU8kRLWwtd0ckGDx5wBxulXzwEE8eHet2n23QT37EW
vcej2IqF8Gc7zasQVIWrvaoQ4S4yB9iZu6zq6LLO8zh4HigCRz5NybIlC+7TS8cg
Kr4Pscze/BQ2pO6ZHIsLYAMA+3q82tF+tckM13HkGAuOOstpsFvKprOIhSW8aYWo
zbpusZksUp3tOhQOEAkHfKEjLrJlulMD3PntKZFy3ZjPJ6OrGdHTnekARzSqzOMf
JRnUvOOMQsKy81CZAKJS4fckUgGklT/fyLq4KrmbNwQVl1YomSt0w5KGslTuDUGE
oh/cgMRKFnCx0LPafQP71ZwA12AU301JiL8kew4y4nZG7Y9D6e5QKd6kWWn124Dn
KlWC1P0C5uGZBW9c7QnBvy9SZaw0fMI3hIRr674pYZtwoc7QJbNbSWDQVQNeoKfO
GFhq1d4JOwABMRptohuo8H5IQSlQveJUXJti3OrVCBrqCoIbm4cg0W3VrH3X7o6w
bc9GqVOCDQIrB0BHoo5JR9pxmi1tsiZJOi+yQbjdTAVzWixyI9vlHXotPjc0YQHK
rh7/UwQeIHO1ivjDwmBJip5GyQEvWKLKsedbyzhE2yXH0B6jsOxiE1yay68F0z3X
Kz9WPZFMzd2H1aBxGh3bBkFNLcTiEymXYIyd63Zu7lLP/k3V5E0TKiQaoA81TvV/
F60VGMc67TKhy+EY/CflF7/W88e5VdztSUo2Jv0h4upu8MYzN7vyOfE28WtCsZqG
6T1pOzwYYwGamWTc3N3l9poqRcbBKlmcdp5iSSIri+SX7ZJDQaV0yiQwgb9O9IjO
Sa4E73oku5eNWvMXXpQo1uUe5MVZpwRdU7SZ9C096XVufiuvHlv/99QAXukYEdDe
OrwV6GXfZinn/pn5Wl0XCjV1eL2n3GOT0vdvrm2hrt+HzTGRD7dlxucEIwNGHAq2
hDtEtzytI+e9luS2vTEXqNwiQbcADfxOyn2IvmAowqCeEIVNesdIiX8vstJM0fh0
mZLWSiZ2WMMsDVQh4m8Dz6sraJXvdL34xOR1ou2qoi4DF2mEBVtSzfATeoI8Qx5S
1akaeFMd4zj/GyqB1WXvqopgIi1Qa5afeVP1vSwT+hPMHHHPI5ySupR096sxc4rz
ZiqAlamhIpwn6e386O8xyGfpNULom9xlbQ8qNvW2MNbQnv62tJ6vUadAs6z0IB+4
z+Q3DeOy/iXdJlimE6DZaa5x1Ad2SyKLaO7V2o9uG8zz5812YH4X0kGe0JVJLG+g
i1ydPADxoUfzgtn6gEn3hL+B9/b+Y3Xk/TpkTPgE68/uZlxjbYIX1RE/80Xh+5Cb
AlIaBmxm2Pn9MB8MgZ1bXDYrB9nGXRqzDx82fgFEj9QMRlVE3LWvxBT5p/DROcLb
/zYvC9XtHZ0VdoNudImc1vJa7y8n+X4qFJJnsBL7gWt0RydTqK5RuNBbLndzQFxu
BcNbOwBo35oIlMjUuT6kSKt2jquvlXs0iHfWNgvY5B+i819AYFEECGn8wfGeYCjo
dQ1nXJubHDlGvgXQ6sH2mtG4r2q/aMd8ZYmxg1LwVeNexZ4Vmg506nTIFGuLdPlY
7nH+O5CFv3GHeHTsbfhuSoxn7tYIRa2kBNPJCHJQebrMXM8Zdg/X+KcFUWf+SVWX
fouMyIZs29kFp5/zk+0kRBl9pREl4A74VzXvYtdA/obkHB42kW9+8bBVxRklTUIA
+xIRhvcE5Oo2SEKnWM5pjANd7l2/M23wCSMPfLnJkjkYXXQplfokC++HMldY67r/
3cuXA7/RWhWAixidrUqlS9kX6pXKyb8my/AXePN/XcPXGyCE5N7uOGMYGAgCuBRu
hgp4alqRGyHMFWy2IucJpyZ/L2Qkg3Qc8KpqtbmZYLs1LOBuPqn3nWB0SxvpZmJh
msR9lbfynmZe4E22TfusmcRMRTkrS+6uihcAypHNaKasyc9WQPJo27+YSWQujaQv
H+h049tTH/aXf21oKNK8Wp7I6b6wJ6cUV/ELGi4+5cALhjmaP6R/W0g3ymr0EfB5
TjJfNc9x8tQveiPwPnnCNNS6bQqYxl18GGe+zXb3a0tX1fmput3FwIXonNU3hDnL
XG4ZQhcmta3mI/FjFXUwO5Tl3M7PuaKjAcnvlWWHjExcDjtQ1Z/ZefgG58uVHBju
ML2W8I2fK9QFmVXlzJB/9VMw5+0pXBEjdGERWMWQdgMjri88k0Bl8I6aCcO4ZqHO
Sgwj7RsxrFwWZ9vcBgVSWX8dBiXGf0fjffLYFafBmwQBKF2+UoraWyI7fJ08K4bE
+agWRNNUTvdZJuAlONQ4oyn/qreRuTNfcfC8kqp72+tHvGChNyOcdrPa2B0dbjS1
Ouf1lfBzhqasZKH3KDyYD36dFg66gwMKOAP0cBezBhgvQMlHDrptwK3WW7u8bzZG
Qbvmk7buhLsms7OCuSVDfRo7I5kMfyOkSVGMMd3ylHnvlQckrvThO88+iGIHzQYu
OJiXtgv1A6Ha7ZQ3JGNZ1FQZLpElz4OlQgsnc8y4xvVGt0ex28GuPnMetFuSmKlY
jgH9tV4N1YQ1JwVE+8h5egMNuYAXY00MyPk5AxC+X1YXODsjxqFU8lJekxZKNQD7
glV+XHVrt9EP0XWdxfXW+Mi2tHNtw1EX0nHyAweNpGjEpTEnC0Xxytyyfu0Q79Pv
RsmOyPmw+azzXY222Yhl8Zs8bT0I2ti/mxzecKsFI8jcjDL+wPmo12PhnEbn+y4g
WL/LM1jxp8UHm73jQT6OpVo5gNxQiEQg6Yj6R04o/t2IVnSBUDI/wM/LxGqJlZPL
6C9QmqxSlvGnLdosjSq2bpjHpjnkPfcrRQ+6piBtzNDuPjeOfeKT9BudrxUHPN0J
zeYJGQl/mNhXJImn6dmDIap/Db2FvVCBN1mNONbAGDj6LBub2mxJ0ZlOkvZBae57
0Np3uwBM6Y36y9pb4C/hCfPBy//HpJ7m7exwUpbXU0a3JGxvDQnqMElrbQvBjV3z
whW8X2dFkBSxEvDOsSTJ1M8nqB1WaYp4kMilbtSDXAR8HQezqYuaL9hQ9hRKXvTM
Jtjwq54udGFom3VeCnna/QP1L2Nxw71fnEOjO9WHsXR02ADVdxQ8uOPWZQvGwrCx
BUcmOFsh4kMAzqzNoeQnVUI8aBhnDHSFbjENToW+NZ0MpHsQsiftR6Cl+xAWqtGu
Jt9jQBO77vKpnzBaWC9XASvwkCcbHUU8Sdt08wc7lvwX9j7whwMxWzvEEoGidMpa
BFdVn7/kJ6IcmmR4AO7Zm/jun1d9h6zCOg7uU0kYxckKJW0CKIfD774P4Hfx12MD
rhZhsXOcRVqtVsWKZ+WYl2WcrzGiKm0KCsrmTbdCggoWk80YzRRyqaWJZ6l5qDTr
z5/175fcRXACk2y7jGGVw4m26Tf09XwKezqugoH/DCmyCF2H1uL4mUGKZ2b1csHe
VzCDjynHix0iqZgKoYgBvotwbCPkVQp2tcCA+/lo50piZeP4Lei4noTfaPtmKgSY
25yDVlCGB8kSvSOS75UDZVJVGeGoiCOyweZNAEiKC8/8AW6WwTkZoMPLQWAYDAwW
0jy5SmUD9QCifTkiv8J4EJWzieDp/JD0qSENNvKrxcXPBZQ0YjeQxr0mkd2NRD7V
1UIVKOMcrIIj1KmxqgbOFr3jhOtjugdStfgcprzoVX4Tpd7Knhm0DNBEWfDs53kR
8DbKrQP0RwYrX8SMUdvJbgTeUgZPLm3J7Lvx+76tRkkFLRF75Y3Vobms2qhH7GxK
kbXsznZunemj80jbexYDewJsOE9cyKuKB2tFC+78dMgF5utYPnwuNziSKszjp7OF
huf2HdF9tAB0wL35NNYEcjJhgh/ULUJ/BNknW1HT2lnnPeS0z8pKPdnljBJm6Gib
k0X8Ait3gKfvgG6Nvb6dBz6fyqcWQN0pUmKaKGdShde5npARfM5Xpalk7Y+dnqZE
Kqvx+Wmc6EKvYEP59rpEkysbOLs1Kk1TfXFovTIJVjqAFktYZKJjaLGOCC5gi1Ls
e8ECxEHfA+ouh57iYQN6BQTdMBApRPT/OTmpkPVvKmKH+SO2KHNisSQIt84clgTk
DR0XMCpBgVIakss8PpBASfw3Y05zsuK0lsT2oFbV7BjOXh5+y5kIS1/gaqAF2sTj
Ukc4zMLxOVNCiCDnkTDCXZsvPqKxP8xMEA7UJreNwEpygqJ/WEc190piJCAFaqn8
l4Q/up4IQlBaPyUMD3/HGOGlK2TM1/y0+n+kdWjUpIk3R5+l9P86v0gir/mOzIVf
kuUZFfk/BHiKovmsPKPN8DpiC/co1qfdx0e8htEI7wLQeGVBKVZfjy3fqb/LK5jB
/dcvHz2oyZX4Cal3EWDE6JuHVeo6qf6eVVSZU7QjCjkJMvoV6DnMV7hHG0p5CLxJ
YTGccaR+H0MAENdc8vYSVbcD5kFuVexkNsuLSZ6e8bUbn/NzRDwMGz1ZI8OuTxR0
yuoU7vYpmIhyM4IXiabdAvYs4NOc9lDRhyNtB+ZJ5KFsES+toSHCAfXrjEY1BRU4
zry2x+0yl35bnyGEBUlGfr97+0JAXmizR+hPFm5XAmuvhsnC/Va0JUGWbDUzSMQs
fUoDZaMf5LqOly5ZFWVM/NYmDi0+GhOYWneKss8ceXJbIwsrxfZyJb7LTaMLSFe1
Hzoo9dimPUrHyH+vAXfeXF6L1ZFbWoIJPo2XtWzX0wGWRZbPF7MxEs3OT4G41Xac
KQcCkwr3kCc/+WE6JqVaMxxSQur6RFxgLVVzhBUpe6bTuVmIF0cbLtu+DZfif0lh
mwlrzcdgwLeEHswA8SQs/q+p2WsNZjILiupqlJvqslwbS8VX4NwCWgh2ftLNSwYP
myOhFsZJzKBVzkayV5xcHCQEfTkWy+cHSPsB+PhSoMR5CWepVBEOf/O0jUtSGgv4
irJtWfQsTpgYNU8YHIb3hmSabNGZ8t0s+HLgNUtWEHh3kti7rmhum8xvVXz+Tdsd
fY3BN5x8fTFTkacIx3gvTAQxX9keE9ejLRCrv7GY1rSv2e/e4gca1ho1tfeEEu5s
XNurT9Hdn496y9bE1OwHeN4QgJCzllEmEWh7mvdY+OMn4Xzgaqz8Y80ZA8Bbu4fy
SRPBMUjKPpVyDc7khDWkoGB3JCRH0NSBMZaS3pEMU9tSVuqVoML2Th2zIFT90Ez8
RWj5fQH9k6ak6i1bV9DKn4BBq5tLikY7wOzelBstiVdKvpqZoiLmBK2l6P90gduj
tPKbNY518Z3hg+Po6+3zbfdbqjqH30wpuuTXazfF1JuX0Z5cYsapy8lFnpmsQDN8
TYmAtdtBrE5zP+qL8oN2OCSzh+8y0dED2lTMjOVEKab9NpvxlWg3t7GaM0Nb4Smj
jRqSfowZ3aOfJoOtGtx/yAYjJd3B08bbxWr5gkZ7eixx8+IOmIz8zOkjjez/rim6
kU+xzLoRdfuWTtbfYz4KiyLljc9Z11hFSLxUb/dNOanJI/BVtGu7hPnUr71MylCo
W98kB2ErdZI9c248w+3ME4c+5eaYPf/PnYHLaVOj3uq50c2BFrGoEWN0KUYvHLw5
Iby9dOFnUh8GNWkWVYFaf8IOJ5K2rxH6e4Atc0gju6cdGv8dTHt2/tueFvOJBTmC
8qku+2c1nxB8SAbRRVRa6eo1pwtdus56QPA38zrClrnQopuJB4dCf+/Nmc+0YzeY
zLdzUwdYKRPrT2HxJHFT1WFABXp+rUiod6+1+1B4BktaryW3yJX9CSlsKqaKNLcm
etqf5CEzhOoDcz9NyQi3fBSMKJ5ryuYwd12TckKDTYkG/5S8EtDUjV620F7rH0/b
YaygU7rbcyY1ksJgPcp2ldSqnbd+GWRui78YqhhX9mqLa8KDh4WTPcgKrW+WJRcu
6GOCTPU2NovpQfz9Tna8mdLvRX1RdPk0xka+YBknHCajW5o9o9+9iHlJ2I6BWp71
RlM5hKNGySCO6M7pHi6DCHTaLqdailJH5q2GqOsmhtfq4UU2Do5khsezDugaRTHn
fxXjqLY2X847kHeybpUP87DvcaWMNiLjTMeXhMacR1jnDJGdSGKSmRcIge4BuJpq
uS20IkkJ+UDoHsg+isSdytLdcfRlYnKqRzqI6by82QVxZFDcFW2kKstG7eyMUFbl
FbvXYjlk9Aewz4anUWD+NAz9Tq+Z+57DpdXMgCf5ZqPn+SgiKh9DSYYY5byPpQgB
Ybi+5BK/ChU6bKrk4tiIVE1VCeUa4W23uK2AYw6mNP5LxyFkSmGCEMtEpczrrsP8
i96GGjSoDnCdthPlt4Fj0GaIPA19fYs6tfxHx1QwYHLRa0Z9JyFecIr+IlywP67F
DAEJthgWfyFMb7hQHs6Pn390S+aOX2qgyRIqEmg59+bU6f9nKJwPKKj/fH8lt5/9
ByxFt75klQKLJrSoFyVJpd2kPUOmqRdjFvV0IjEO9ngXzoYFrSiURKmmWu2UZZLI
NNsLh5ohkwl3xrIbMxtHsGnhK9jurBuoW2e2nsIUImwNBU7suvPuCUPMjD6QEp7b
tkc0bTskPFflH6prSvCirWchnm/lxKwofr56DKINJVYYcOFt9quvpcqB5pDEk3VQ
p94a+0Dq6G6rb9Pk8JxzixjIh2IRNgYXC7xzoPoWHb7OnRaD1ehhGLbz5XxQxsIm
p6Am1vD8UATgaf37u1KAgMEWqu/4vuxD85dIIF291mJpbBB8AP/oFOBtdahzUKUi
8p2/igF0p9VeK+7l2EhUI+g0sNg5ptDJjCVfrR1tzWKh1xi5hVhOKc6GfvizPYmr
8Vqs1PIgXFVamFcQRMvFv2YPPU1z9wMeCU/skcLeRngNf0wVgQZHWfZLirPixL/9
hOUrLA7DI2vwQ11vA1ipei3ENMYxzV9co6pnlaIpOTfQIbtdDa7f3+abDqoIzjlN
l4O2CNdC0VeHbSgDRTzhLpuOEltfXieNr6Yvivj8F3qwS+Lt2YGRhl64U8x6CUhR
tbBornjh/906lulpEvXRHe7c2w0EhZxJqgnKFuVmK2KmaCYjJe07Vrn/p1l6vFvR
YFlDhX9+ikcUdp34OGKYD7ocKX1Ft95xiThlLmVto+APq5Z4UkYDUGKpMG+PURmL
2452bBDadBmpuYG1sd20+BKDM33svDIviyXoqi24SkiENzeDzGAGsI1hbHEL8kxs
75xvRMVUwNrGExXLOIAT518CmN2f0h8UMKXlujo7U2tSEnGw+b5xqgjaRUNrJuGo
S1eUmH8rgjGRTIkXlkUZksyvBxiANBoHszB00HE5h4KWxnOoPtgOLnVeNJ/P9OSu
qXS2KG/xUUu9pJr+IkvNPWP8IPQVJ4Tp3Gffhzhpqc4e6cRnR4RlJIoWeugxkt4u
fkRbE05K9l1mtufrV4mLjFsWejJI+1fHHNAdiPGO1mL8cHe+wMNJATLPziTmqrjT
aydaUEulYWoc4OFDKIScRzMk6hRqGQlqAJQzyeXQ+Rgw6rbcbOWh3VUhF09Rm7w7
5XuIzGevV1XieAyBWufUFOcJ3FCZ4C5dz+FtILBTpQFZIKYsiCk6MPr9r0q/0O9k
sxhT9iftVQYll6swbTrc6zik/ixOhk7diUGbHSm7ox/2eJSk1hXQ4CF9TiPLroWG
YNv9d6VmcoQ1tyPW9Qfq6QT0QNrcJVyGQ49WyVkAqsV+acAqP3by3dncstsjHxW9
gbPBe7jnnyKLPS3QWgtHFCFHGO1aXaiQCVoruiCoLc7tOtElSGfPSJ1X2Ddq9iJX
jkSPcru7gvOQ+rS6+JvMKcYSTAdEoyhnBHEJOfa/nIImYkXctAIFHPQPkWbqCOWq
Tyx1Dq32zYDiKoLSKy5UFQeoTG9J/ulSHOydoDEDGtRutCB90A2NsBJ62UlKBRDQ
AEXyAE2GhgD2u0ptGRQdTKgd2m27WUeMXneH5kUyz7GttyymG8RY5wDFniulWYFv
oVA5renhA3fai0oJnCSP+k29MSivHtZCXwsDL/pUaVTq+ZcugG1r9zGBmmL1zBu7
ucwCwNewdWkvpcHWNeXS/ygx8Y0pyLV8ZHGwmHG81vsXzu6+jI2DOEf6KYbcxfRq
1Y72ODOhKPhdhxLT1MTnXizhcMZc2OcVVd9FfVrILoO7Ui8qmah32nDeFhw08lBr
kRDrONMajFNOUhze8zW8LqTLyE5JpJ0JgbC1CmTjUuH0Lido2h68E/cSV2SKVwZ0
uFcg3j1CvYpOplwAqyjbpub+sjSg2SA/6SFgumqKTFGodinLXHLBFQBVwsfRBoQc
2fMKxT/oYqZ/JpwdAgBl/Jg+3bd1P5YSlgmSdBBIg18s2Xjndx5d8H5yx8CGQfp8
h7YROAF8jecgvDgRmu6g1gL3SxLYDU0+DHP+NVIRBdtG61ftsvYFdXgjZiKhETou
uWJhjLmyk9au4rWo6M7hB6TjJm+EupmwDHe21jDZC8LVS0llnVrTaSnEmT95fTbF
kzdF1ZrpaX4TvzWZ8xX6YhslJ2YoFjaEUn8l+a3O0iQOEY5ABzs8dQrY9yYjcK0v
LjDzXetGOtkPJLDSO8ccDuz9ZCp0ayIsIwaNSqeipm1bxhPNYBc6z3P/bWNp7t48
fol9gW8Nm+spHG4gbaR7KaEN57x3l1fXp4F9+K9ueFbS//yn/b05UFwAsJdjFR+n
Evr6t4sYsXFZocEQpaxVpdB/1FHBYPEsu06jlmyCEYp4U7/Yp9Aw7xb/3Fet29xQ
P0bTa/u6MFJYJQRnC/99ADm+2YZcx6GfTAdE58Im7erHB+V+ePkM+1UWhGuohUAe
hzNoWKLxtnWhbid/eyAwS+T30CGq6DTT0fDmo69UuuQsPHV7W8FN+9bWF2yZBwWG
7i0Kc474hCV7a+ws1aJ4EmMf8Wq0xAF3vKhLH3mbpbImMT1LFeRayw+gt7UkuOQX
Rp5E302fESPiK256rBOIE+46YcL8vXLoPgMjDJ544Twmh+qt1N7JJb1p5O1exWOn
drpwIM27E/jxAsg6bPdForGEefz1gY4B/UXSYenwctPsSZ7dXZ2oInObhIC24Lvn
O73hSCRoo5X9ieW6krzytJAJ0NXhZohi3jxBIeAAeSHzT7NSHz3KSm7n5AHgs4cj
NpvbSF44HU/ByKyfvGospAropHlLLT92o4zHDVHC3/4L64A4ZLVFemayd5zk49oM
8eKu4+iGJ7GB+gtdZl8JagvB7higLfiidgw3LUJ9gsgGKVA/Z+dTOngoq46fPPlS
82ETBIQcuooitv1K61XTIpdcjM6bx7jdNgCZxyzI0B1EYkQIeDBBd9QLaIPpvsC3
awTOeXmyjrMbYEFdbM4MkFPExIBvLmq4zJoyxMfM6/u9i5stEVa4jKfhVkWBMNAP
Nmm6LxhbW4VHClxHoHgqJETR0WvAtEFhHJ8yh/ynmBbt/FzdGgeu+B6oKuwwGqEa
MrMI04GoBEer/CzUP9qoJ1QbfqAlWWzh3/J4BgmYDWk16GGxaKeFaUk+YJOta7+Z
VHELFIFMWL0p36Xa7rU2N67JOqPMzMXzZlAPF5x34UCy0CHLoJDLszMn4oNsncOY
TL37qBbRUrDUPkKi6Tn7WZPPvq1xnkoVFU4MptoEs821J8XsKzyB4ICddMGqvSa2
heuI1hSkm9QF2/Ytt/dElMp8jN2EoQW4obZWgJmnCNQZkRTPgE9O/qboACH+Uf+g
eGepkxChSvypVvynLnG7v+ernsYNC226SSZXTQD68/usxqDeS4zGIIaXr7eEsqVE
U2U1A+wcpsqJ2Cb+nVoIP99sMV1u6Y/7W8BjJYW2jgHv8Jiwy5gkimgku0zEoQVo
/yPZbcuxDx6gHE7Vzc8SRt8ObJWYBpcVec94+UHe9nXwQkso26qAwhs3dQGsq7y8
yIX5IPN06RZijKtcthp+mt9iPICpNf++8u110I0EeQfofPlCoetTS0bzIbz+5aDp
IhhWbzSG7tnhgDKeoexOT8qYh3EmIGy3k+U8Qbo8F9m7LYaZeYPHdQesusXQtSP/
gMeBnNdW6xeUMLintSi5AoRl0wQcC3wJa3e1hK1mDDE4dSmcNTKj3D3U3sXXDdbr
Qca5qONyoDATyiBA/0jVoC+BgKHlSshMvBHkSzTbNU5AzXQPY7nNa+wCEPVanYFY
jLNhtMnfl54+Xg6027tIgpnQi2QQ5kjKn6W4+qo8iOJ733qT19e4wlCG+zVD7ta+
SQWGb1ADWgKXmyZqYlDMIimC78cA3PjerQ9VQwyHKhhQDQWDVoguO9A3f/RaeKQt
NRcxrGbb9kJdcc8P/kWh/ntbQBU8wEofqk8E/1wrzUxEmkNRPb7S1gmmtZZDX1Vh
exAKpac5vnGKAPCaB6rRpG39ko9xIOZzagiBh+xWzWhBm8w7Yn25pknsfLxg4ke0
XqFBmqlmZzzVGHgaRci3uaaDgGHAVdsZOj+GINzNRCuNrcI/H1ay8e9uDXkhA0YL
W2kFXlpN5TdT0dNO4ykMtYUUbPNVZpe8htYqUhwEag/2loDiSKNOh0g9rXYyLsEO
0saXRgKOaaeQHcilh3lcpzjCqHGdPwevzKK0zwZxFZn02hjq8SOCvZ91dwHXT8AK
jnplZmWvT05X9e/0DdXGuLcuhfFhHyyFY9tiudl3Zb5UVahgMMTuf6JQN/QARYk1
ifgrVnVjvA+rmwtWjJA/pk2Su+N39Ew2PFDIGeeGLyUcS3a38npqhG/2jm9Mebj1
AigE3EAVGOjnupj8OLuXZhGWCXi6++3k17oquWo4WFQobu8tB+rIfUDkh3elovCb
nCuYDttwjVd4EambOr8fycw+vDz9eKNAqeAaYm89EgO8Gq8a91pN+OFl6FFYybAx
ORqhazMhxjfvhz8pyw0F6hjO1D49tgaXyFWgJmFx13I8IoJ0Qbto7cuV7sI6x8C/
p5vBPBv3Fyn9VKF2DsBg/cdWaBa1xCOqVi1mSoXSmacrN8ZzYeOxNhebzBiuO8Hn
4u0u/MrEQxXYKfrvsXKcgB0CwmIsMMzFZYgVejQkCDV7SuJY5orUH1+QmNGTMexh
7+6idDPo/n56xNDc+sTvVnJ0bJQdMgQDaOsHGaiKqhHedO+GeeYr1O6hFsS5S5gy
PSzR7e5o0dvSN9a5gMN6DEsnH1WSvFj13chO0VMbsdU+lz9gfHDJspcF7h7o6Rdy
GRkZWzQC3rOAWBZ/ForXDGGfuKb3R/1Vi7lq7AArhkK7r5sSLfrJi3/SmvX3G/Si
ZE251I8YGzONUxdTxdfqYW+uLmmBCiiAHXGV5uz5AiXOivtYiF1Ooy9a6rDwdDFl
0wGeay5EextEWaFPTOmYfHCwLdybNUnix9HmYG6ORTGOgtfcHkET3pl9TVN9QtqK
Wz1DSnfOLOC0dGtpuK/A5yRsrh+5fkMoDNGl3wpNveZc4JF0KF2WniN+ymtBt/ZU
oWqmMUYRWpnVQx+Mdy263P4ExQYxGQVRgMaTmLsk+X3yrW+2VaTOGqJOdDBecSyt
JVqNoceHChYt8vSYFrETJ6QCXdvj8bhyXKEqIkVcNKfmj7oePIr49np/0t1oqOnv
7ai85XCw8IxUZhROTuC8FuyOetgv5ZNiCVhpAU1nY6LJ3OgNRp+wHgR0rIxqZaip
m9DAxxOTl11DF8IwatiMIIPRtlLkW6yaN9yjFIm2FPD8x1ef4g7DPTgcwOqQCw6M
Bdk9QAJmwvKFqHW4Io+pFwO46/qrLYBj29qOHLjGDdA+ix4hz/EpY5lSY93ESTZJ
EYtma9yHrMeZekq54u20T9JBwuS+kS091aH8UPqQ8Sq1Uch3fBTOZHmypPJUKYmp
ivs8SjYY/JthEF3mGwOosNI1TnzBeSxr1hXWAXukm6+687VGLtO0rKIKE6PeDaOA
kAI6Ux20u9PWLxo6Ugu8bnf20guFs1SUcPTkVw3CrXz7aVNHx3xiQf2CnCtAyPi4
ACXzMcH82g8WKllAJnf7GyuCl2MOyE+CPlUUJjq3rR9qpih5ulJSFksidlLnI0wd
+qmG7W69ez60KuCvF57xjcqfyvwjjDHkn5h3lnd09HkW/thAG1YImgoDsvExvmEa
UH1ouPdFFT8d+HZFSBqJKrnBZCKJH7iUCG4pzdUD9chXBfy81PecEMyDLj+YgLCF
+0cwDUZFPhAoKtCz7TUBFfsm0qPGAdEsuJ9ujUkZ34diZNEEsawwgyUCcb6r2/Zt
lz4oFUB6vNnpOSUJf9zSxDoU4ArZLUGO2Z79kp9vVre2HIjAvsPCrpL6egxcBVIl
4Cdj7JmOUtJ1OMo/kAIZYMaG4YVv74bCWjvTKtMRyuCWqQOY1dijuobvrUfVjCsY
aF1lEy7KfgJ9DcX4ygSQP14nITDI4fwDIDt17+2k1/pjhR1cfMI+3LNaSEBorYg8
VNJYNNANg83KUIdIDqOvN7iaobTHNVwo+F4CQ19NblG3npWuADgH7/le1i/Cqcxm
+3Dns4F57NEMjBQDpWpDpllOvsLYqosdkHSim2s4/F6uri8VGtVQxv4axtO8AW46
Lw/WPIPU308EWLNdtkbjqxdqQXjhWW2xJksuhgSbwP4feJ88ftYZkQnUO8FWhNUB
eB7ZrEYdzR1Az0EhiGlkZ+uU1Cur0k3xEIBuSdBN2TOTALtr3XHgAXUBxLR2hF9C
Rcyi+b8JnPa25DorrqI3La1H+/CnCOsFOTP5IUMJN2PJ/2SqXfRZc/AHQe9lXUr3
Fi00e2vZAP7uN4+OHYTzeHGmqz15c8RpEHYHtn8r1GSSrrJt9Xm+FOrB2cXpBlEL
YUEFRBV59eg7DCkrXvunaBiK73JmtCjllrNcJ40y1DgUaJhqUHFNTKBjx/lU9neP
CTHTOkklFkbaNSHqZeWuObtbYp0VFLrPHkk4eRHyUNr7L1j51XxEv0xny69d6Ni+
pgpTKIeq8l4CTHguE0fLyC4STpZCXB49fhorRQtK8KSC4tL9freaWivaBrfiEHCE
1ViANHZ9nf3iKOM8E2fKtYKfIE1pdA4JySPV4Da/ZenHkBYXauXSVt8ryQFzfL4F
BpQ2W/5u9ifKGB02QMTT9YSmXVRUml2pRL1Wnw4fE86Y8nU523NY1G9tqs7P5Tew
JonCC8DgV6zLVlNFSd9yzAjHG9jvLDpHU4BHgo3oje/A78fz//B00Ku8WzkSTatq
djMophmo5f4Q0dW6Pqb7AQk+2L3DCemejgo/yG+dulQZ4CTFtI5IjhGyZvpMoNvD
PxVqE09Xb3DjIeGGCryc5U/6ODfZgF+bb6OfYw+pzRImth6bRx1Afuq0l80B6h+/
dl8Ot+MAMY64BQsye2BdK3x/opg52gv9xuO389MfOXEnBkngztL5F8YogZv3JvIQ
+MmmS7L6OmVv6WRx0VJB7jd3FvTWXRpfvnMG4hhL5R0FdpABgNwx6xmnod46guD8
MCAsFQv5lxqEbRSgbxd06L4tObv9PGrvW5z3hU/tVTIU/cxDb+J6vAaAj54ppaHs
NDqUS+CueVVL08OLvtTwUMnhft8I1eoCmLzke3eEZn7d8GGavACUBfFqOf8WeXdS
GAH51OVvszDfo6YyteML9r9fc32TOgKRCsl3ldAl5RCN+hHwPM0wI1fJXkrrmcgo
qSXd5eYHpbM71MwwOtcfpLYdDT9NhqMFVEIGCbTyI88KAdRrI5+bu8dFmtlCOVpl
poOeLgI2uDelHpmt58EVH8s+WLa15ufAQ4UbmQEosrACBrCK8nbhKUqW3mzDD+hd
JphhGDgrbtBqQx3TVuYKnDHWvBlnUKaXx9FotILZ7hhd/CqtNiGrRDsr8VlOZjHX
CNw3xmIZ5T9xKTHJy1J0hZl1CgjpRaf/ohHZBQ5S1tcDAs8I1PVH+izi02/Me5qH
ytJfCKqopV1858xV1j+A2QLImzeb8qOCEzLL2bSeq6fbOudaS1R/p3uDPwdBv4q5
0IUgL/HsGcJH3vhAq1BEeHGU6tMJEjVwlNJkdq/eBwvgTUuHQ4UR3CufqqdcQHW2
PStcI/yC0VPHznWOHBzgWkWWzCzNrG/eWz4LM954q5aF3EvQynaKExvYeCrtKX2v
9JbEWFmnwvU/zpvG7fVgAZLDLCT5F9yyd4sxNa8+WNa8Ec1oeUd0AYzo1tMdzEy0
4gJNX0Xz7k9SJQ+2MNyOw4goDzBOy/+/Ya6cLDVoY/DkNkXg2DML88h26XQ8utgs
d0gNRWsEKR1NY88DqmmNThoMHHpXsNJhbISngyl9f5AOgCL5UonA6djZ4EPGx3NG
SMGvI9AVK+mGokogkiw5KOmbzPf6Pk5aD4UPJ9RXQ2F3bZLh/sWSXBZXStqiJEVX
6HDTU3lRQ7x9Ak/2WKvffhspg9jERGOgTSRrGGbdlcaTwriw5xVXZOF5gAoZM303
dKN+OSYfC71G29maEdpia2QJCnvinx29iyxLUqAD8kMO12MFTP53TqTCcLl64Kje
QES768U2JxPXAq0WtH66sXttjME7OwFjersfBDwzRWNbPJEIyKSVjDYZEKtHsijK
javYViHncKFaucOs/jFn3tTBhbg9TmYtNG5h8Fczl88Dp0cGpd/HCKsUkzhM3CQk
CxZO3SznvPDmZ25BnmMfnUSQmCa1KArCABmMqIV9knifDcrTw4+l+Ow7e3Ej2lEl
HJX1SyNF/ofFtlSwTL/rHxpxhFyshKP69e0X5aY4lgY/6h4glG4RdI4JtoqV2Hjm
1nG4PM1eQEosO96AtRrQPIX5JcIkGRXeswGtpuGHF8GJ80t9u01J1WpwumaSB5Vl
loZKo0g91+QPT17uNouq6/+M5fw/vc2iQ4cbzALlhVpa7qdQXLMfis2ncr1tGi9o
vslM0YXEsKgNkKDTS2G2fYbTtF4r4k1RO+ssDHEPOie72hpUI8wgCaKyySjLeF6y
SaFG5hrBMnzBQqNawrTaqIqTt7vvUACMOAJomLf0UPvcOfmwBVGAliqzNGJo6xIr
JcnHLZf//H603sFdQ3Z1fMV39cN9njF3n90CRk3qLBWpPVppH9j357T/Mp577uO6
5RRKuv2joTTFQV2T8pEnbkJS5/H9ZU6dTbxZXCgC7memSms/UTNzkOypoFmnRMqi
mGt07uEtpaZW8nFc4N9fNlB6qaLwyJynASeRBaIPCZyjfbzKp0FukgBzG8+1jeHG
nKOCSSknUbIj1XHXq3s1K5e+EMVB6B2z6IqjLaP02lL7WK7Iobza5fSCpy+RNDJV
2HoVGkO+NT7GeD0XpX3mCZhPkCg60PWqa5Q5KJhNfbJ+yvqAYKuPY3tvArW7Zda2
/koBl4djJPhArNtSdveaG6wGq0XD7AqVzcMORnQa7hjM8kF0eoP3lR2y7qTjIjgH
qOT8xqDQTwb9X78pYzkPKWNpanxatbWc38+kEEdztyPS2qkePOi1FNwfL/wHUgT3
yQkmQz2zgsUK5lk+TvoZ4gY1JHySON3PMwpsEeWsgPB5XCQZ6TXP4391gEZBFhqI
Fp/RQMhfxc2Er+dSmr45idk+OpwR/mdCM8WfcbcVZoP/9WxvtCdky2gQQsvxLSqF
qvFoUMLBb7mXcneQOpGuUXoO+hdpYel44LcbXhuu+ZAkzgARBWQH9h3nw6o6TWRF
f9eGpMbmjXGOqAy6PjqwjQyTs4BPuo0MSai5qbYroAaz6tJ0UY8Y70pKdcK43XJw
CMVyCvPtENPWM356m7atpoFm+sWRkaoshhfV0yjyI+zueNxOVKy8lrUt8eIbeJFN
Icsp8LL3RC8gpmSvPd7/FUAx37wRjQPUY9J+CPaW36CmaYd4bfv0T34vhXYqEJ87
rWclMe/KkhSA8ne0fxdp+lOKeSXtIH3JeBUh3w+vm4eAKQABbJaSGUmrALvbLPts
hSWutphz107Xi0113UKfYri5tUL3yLbzQuN9VwT7WvYMDsMvOVeAbNpw/CoXQvpl
LXNLjUIUFkzgcHePLSwVnkCT32u7HH6IiM7QyjlmSXIQfvMfQTX0j2YQiJ8nTnOB
uXLAXAIo0WGJCwP312y1hKeWGcmQfVUTdSwjw3neR/S9Z+CYGscYGMHZAEjfPJuV
7fXwD4e2AfXLrQvC0LQLwg/tzJUBScCLrbzFlZ/YSnq7LA77V4154cBWcPoZTfEk
PpvWMzSOp9kgUOnv/geBfXnmUPWq3gMqLfpurP9jbBc222DJm1jt+pR+byb5Ams7
BXe/Po+pCIG60Y4ihXHgkgkE+AAXAvGUe0MIACdXcFZfxOYL38E6YUCC+yh74Xyr
zefH9Nx43S+XBXaMC/ScSzRPHTjk8BmjXVvJDVqNDmktMbOH+AUE+BOe2wFWo0jb
JwfvzMJiaXylEZneXhu53cr4ZBwI5aUx5MDbVg8HohXtsqhqpyT+OZjL0+UqKWaE
UKS2Aehp9rHVpqSKqBRRJbc6DQNuZ/AWddww2xWEwqM30G5JS0HbJ+xghcBwEuqt
KOaMxxHf2+0rmgb4cCdUL34b7uV/YHbtifZDK0uALARRaqGbHsVIAOHo+h0QTGvs
pQ1GINLmuUnD4sTHxAwf3W9fAiQD1KtP66pn6L62W3t2RpKYGwfsofBl3Y7TeBey
0+j5hWqXXTBtrvgwpIiIptP77vO/4HdcccaIWonEm7DRVhK+XpwEo8ueYIhVQmBK
0o9tmmR4IEH/rgSmK6KqfkRYVOV3CqyPELO9883AA/YhXTGLV8oUC/ailgmxY4T1
p20QsTTeXRC1opx6rvEUajROIMEZbRs4nWD/JHKaFyQE5KyMo8FSTydJwMgsuxPt
dvCu3fIVwwrcgs3OkY9FAZmkPl+1T+qr2lebWANAWgT/x42DScqseu7nUvTM1exI
3gqFzpAX3SqjSORfMYwgnm1AFqzdgPqBm8jVQ81t5T0uk/khcdZj5LlO/sCG+EzC
MqMNXELSQ5M2vtqvD/X5g9o2OvbKsTIKud8DYLZwn34DBolio/A1xWnsNScK0vVU
NM/E73GeUH4lsx6zHfFRpuM7lTc7k4Qt3ikmrLVdFgAvAHBi73ywMJ9xjFtRVoH4
XcIJivdYB1iwM1zRFp9mBFI8cpWPMWvx0myYGBdDU1QnqOFNVpqg9COigzU3e0Ke
JUT30pA1jfj3u768pEH2waUUUzWAqcesxM5oh/s4Qc5ZAX23j5XTXoJd7ueHo8TR
0qJkVnSlPaIulhJTpssee/xozJ6Q7w9Dhwoac+yrwVztae64SrvmyNN0SJ+HJpig
MXK1Mt2XDDDiZRfTUtCcWLziU5h0QoOhOK0W2q+8NdnneDvzmKSTxDGL83stet2J
zCNMU4OAqzrIEyy/dxetS+GBCASghH7D7+GvArf1x+MAqCY9kPFJg4QQiRmeKZI+
E485UVUtoMQdTG9x2c3Sjw+gUwajmkqmTMnyj+Y0cqk3pPU+e9wAsA3e958bTUhS
eeCIw4rkA1Ra/Lv3PPDH324cTYwaaSZ43Vq5LlZhqxN2NmRmxmoXTrcMf/3qVFfe
ZXmzjYRmT7JHnvl5/fA2ca5TeADWiSQAgEiG9MYNctahNzhmOJea/qHJf/z7bYqj
TXKM3w33AEIvkxNCCepihgkCnqSu9nBG0lrTrp1P3wxRFtic01B8pk4TUF7DlvtE
cXlt+dZK5EqPTzZACJ02ABoTHV9VFN489+NV11xAZ3qDemYcG0QfFWS2X57KP0IU
Inya75ZB/Ej3c1lm0c+ilzA/0oTsbzFjDaSHxCA26CzyVZq1yea34WtbjWE2Xmil
DAkWv/O+R3QreaaJIC+Ri9uzanJ4n7XPYQKuN5JDveroRAEuIvkW+UtTkt1tc0/u
y2hzfag4UTNUwAc4Q0H4P6VTeld50vhmy7adifA4LcDfl0exhM5Z8Is1qoZTgCfR
0g+hev5vb6OPHJQATqAIrOKBAO5flb6e78a/+x+fT0n3PuETsB0pAlBAy35zgQqN
oyJKi8N0EY6YVEgVS8Oa/fPjf6JOVMLKiRDPyu+BySZ4iRcHUf+AAjLPjPcgOSgB
dCn2Th5NIhkvgPnHWOZ8cri38XzmFhFDnFh7GVMpmDYHfFJxJCn6+fPnf82HWtDF
6jr6oEhn5xajCN7LGc3tSAMshr1ASblWsBCW93l3mvEr9uBsGoF21DAmw7V4T9Ih
D21y+duwD5x2OuorB7cVBrqrpE66lAq2QlKvtKCH2x+DCcZUUffIm0SEDYCuVCLo
dDoSl3ZTw/GWXxVwe50dHu6qt1L5idBVrIn/q78n5NreLzpmKICeneRu/pe1xHuE
1o61HTSPfPLWT0Yx6DTLZ5inKKbPC6K5ZjsF7IaEEhXjfERRS0Gko9KTV+VRBnf8
6Mx9gxOYDVJ//F6uZH5Lh2yqYy1m8bgKd7bNZCMtGsaTDk+qX9IZSnUQrGRC/l+K
kz1c9pZrPBX+L65yXWIsxC+JBs0FI7k6gjU6bkyGPY78gGqUqo2R2GaF3WTsZKjw
rqozKDRS0NYBLCPHClSFEUTuL6FdIT3xQKvq8/WRnVhKimMwhVr7g/7IGdOVpkSS
KBEVW5zhl2vi8pMjn1udORq0BscBHcROMvNiCCoElImu/8iRA+3GrbF5iivELbF/
9fRNfCAudIlGGYfCbvXc9irEJ16ZPPwYIE2YdxYAT3QnOy+ZDyfvkhCwcDD4WUVM
538zYBAxZeQ4+d3BblJkdMnRAer150JX5qequvoVwChzPkFZajre7EYSClFhwz/x
GKTnbwiOJDYTxEL5hyfQ5OjFy1cijQ6QJbVY1jJ5BXxh3vXhF2NeAzydON5H12L9
VoT0IHk1EZGtEeFjZZHMQ8nQXnrUo06GP+EhCnHdxoceaziNRbhtSiZ/CFSZyfEv
j8Az+WwwOfukUZvlo6ismCFCAl7VihubUBJd5rsbbkon+myQNrWz30ZjnL1nkE5R
afnKAPy93/vJpceEX7NStoi2pzi3Qz4dNd93MijSE16tF7xwqFw1ueeDEoc9EYmO
9CjFpQ/T5qcjdcEr2TcoGcBtu63fcrwv12eIXSih/CNf6u4BvrVuvTfoSPq+6hvg
m2F5RZdKOmcHIetv9oPy5VApiVhnv45L/IeEQxW6mWACyku6hbY6AKYn/7HVWgga
ZWPWaVSJlh5bHrF/OfWpcHSvpN7gWB89zp2d3dvzbO7YfXQI3F8SuSKQuuIuTZOP
zJ9kM+p2SeSbkthcS1bpxoc36jD3s70+H6yZSikZsSUUmDGAphd+GbJ9mDY1fSmI
eU1FlbhOCW50hVafTo1f/QD2LE8y71vYTv60l6+xh+g9EvJIyvTEZNYwpVGGAZAz
XR9spXVDoYNyVUOjhdDh6b/daXrA+H3XwTiVwQhE3wzSCD8EvIQFmd5HNNld3AN3
eVmcMp0wSqB+r5nbf03ToHajkP/jnq96g7zOErAgSxFGAsnAH/cqneaOfeVC/oiJ
hEZGIJNCD7lzrKuR+KBJie8Ia/h63Mm6uz++CuiFkNzHmQFpcqwjxTxN1cv3NeMi
hu04DMEDSQwh/f6WlT2oni0Ht/ftT5uaAz0z9lwwaX6soPd3m6Aaq11NFy9NsOKV
rzZSacCBe0WFUe0N7az3RCczUIXxCeuj6coxYmG08IGhkClVNgYO2LbeBm+8DyZA
v1hvCBBJsvlrldlwwwzuLVdKfso2bodzyRYtRq99J3vJeEQAQza3OM+cOB3tlDlX
YYCoztz2jVOahW/jPnc1vfDujsForiT3lHLGUJKPD8AQDgFWqDkL5STuU8BnhnuB
WteZRbD03xHc1WNvYqpZ3QJ5XY+ET/+vmKsE4X9Fvt6Ay0MBhk6mS9aa7A3gGY9u
536cPrT2TuGVuePwnnX6TQH+xaPCQfPWGsmE9Y3Rh5XhO6gydrzJ6TVuviyMRHvE
LaMmo+RKAjQ9FLynzVhUZAm0bb4K2ZUX0CNW65HCFzpizEmwxPDgZUhlf30v93BT
mToJhuXIAfIHUx9WwlwLr5w6IUzVLTp6qHvvqn7Y3wRLEHR9IHP5taG1YCMaQx2c
cyXBcIlcLfLwiVb+KUPcy5y2B1Yq7k8s1OTfLSS/0XtOLEttZR0T7vM4BFkxtl3K
WR7gpHpffx2u6/8gPB3sZJgtaJ2RoIOEt7YqH/1moeNbnZW5bbPsmXtcEMVJOmab
e7cfpd+qe5oSuiKE05BJ+2FGTU8ZU1GxgJq2+TD3diFdqC3ZuTItVWcnmgaSwhzk
gcEJ6xDa1AhUXWcWNotnVpfAR2YoHsQt/hD2DcpdG0ssF64Rj14y5RYxLC9gR6jW
TwauHEgw2qIyV0H95Kz97aLGef91MG8ZjB8Yu01JivzjFLT5Ek5o3cgYzlRyzaxJ
BN2IGUgg9S/zUW5L2m+5uU945cHbj4BFQci3mJ7yq6JTro9Cp7CQQr0rRQJJkLcT
lcMK6UAmlxerkphRwTG+w1dE2Q1n627DqMF3jOFjgGesv1cnZUWW2tvTiP57sNFs
kmhpRNY4J4mUelbxIdu1ntS4kbnTAoIOvxIvFLGKktQwRWPOjXXNNimOp1Bdh51C
MRzfbZ4fBhKX/pKPtiqO39VcfCkKJZ5EqEWu/mWkQrM2jGOIGA8T7IILegb+zKhg
TL4UQ6b1Si/7eEvSo8WtM2ENzXMD396Z53fi6Zfzcka/D/qaMI9aLFswSwdj+Qfk
8iRQZL+4H+nIjqgUiT8dTmx40egQoYjmlEzzM79cVGZiYxiSFSWwU8JTYlC3MRi+
mvRVbqeUvE/Do3m3mkcUXYywkMG1KYG24NCMny7QyIWgw+KdVY7ytabmAsFauIk7
aqraUKuGSeFVXYbuSRhrB+Bbd9O1bauOTBcJL9Fy65mgAF2xe0L9+zXUc/KQ+QdR
3Bm/KuZ8Z5L5Fk83UbTPEaTyElzods1Y+jISkIfL6mPAsIGs/iCI0WL6SjMyuiL3
R3jVr2HXfWIZwCQ1s5IAhdho7yvkhWA/njQQKQUuzVA6ofW5w8/K415jQ6GtfsaD
7QeDhI9UREwutTMtsyIxswdXODK/6E4Asf9lqqpVIfIFEM8KsPhSGaNb5RJhJ0d1
QqYFv2wXsMyky+QsFr4iOQeD5nu6WfT+IWc5ls9xNnY4gczF686Av71GrYihB2la
eitCdoOArZSFdc8ATOLzgW5ad28ZxUVK7CJjUVdDt0H2z5Ukub4SOkGt9rk2Dt2k
2w2jeJu023MBpWhQUDX8jEFav4+jVyZH7HRmjTIjJMKeW15jHcC/zyyyqWYdtAbV
9L7YoEVEEYGGbi+LXEPZeQYLOPXoW/9+yM9fEQ9cVEcS6mTMmL6+9x79r0JZpW9S
SFx98gjNMI1ym247feQdos1ouIyN9aQ7l2RwL2esSzY0HtF3xPH9Ar0r2268RWrl
4J+pDud/HjmxNl4XyeHD+Ghzz7Wql1aGIAZ+CtxLP8zMGdqV7UoAoOpM00c4re08
7qQ/L5G3u51H6+oKeqAkSOUJG1pW4n2+9J6HwMjBMoYUzqlX9m4D3BWGAv70YPfV
mc+L8GUgPEUia60emcFGUi+IoS4hMfPxmABWgY0za7xDBArqrHrzOaTK3+IYZ280
DKYyv+gaRwWsRDZoKT+HR3gm253/d9QHXb5JzK7RHVNgP1M3ijsoMSVwG7Dh7Vl8
apYPFf9J3o3L/AxKwuu4NyRQZYEj1WqTNBnX9egI/F88z9hokOmgRE7MtwmD5kQe
gipjJNIffpTPFEdnembH0oz66+3YHUxNYHVNZX9pRuJ0EhNQMA52r0kHCRN426N4
iUbN37zGrPxO2FNBGFwgjqPFuee2TZ/Y/i72d0pn+cqIEDKbg/Ge3YIG+BEtHi7G
dRctLPhHDLvUwAPnjmAdHP3pBHsEf8NUFpOiUJeq9CZPD1ObaI54DCPe3SwHAYEa
6LoPb3PGzvk0umnrwgsiZzygeaJy1F7o2vlpOg4Jxw2Az9vPSWLdp8cEd1/jYP3S
SQM0cNKQgap/K1ujIU8UAvtyv4EFzWL6kbsRJvrRDknKNPcW3UMd19Mfy07SNIkP
Q31zFkAOdjSf/eL5b4ZlxxLO4tevYzatZloPNSlOh0hA5G7WNvvnfIAu7E3tYN2k
IsxQ9seSnoSSXNm/fnNOt2Wcj0vfrg+UD5Gmk9vLqazq8qhLASMtI0+jXZ6733MQ
GzGHTddgwF3aza1NAaunUQdRY1WTN/Tinv/9Wk6VXbc04B3joXLMtMnw3htUko1r
8mc9O32Qs63+JfgMGlskOPVMbO+7/IcZEDnqF9Faop5WCVdjtJxQ+D7PnLz9v1cM
GFyLwk0Va8GOH78UpeHxbMVwu2Fgf5zdnrcqMKCH9XBIAdD9CfSnrlOuqXWvwVkI
N+mJhUaJHAY1+kYt/TcpmbDB0UB9a1wvtmBT0lzSV5IE7Q0xafsgGEzBgufji61t
4tU80UmvuHrbLgdlkBpY+j58Pjrzd/dlSl/VJ6FtNEG9xzXYim8McBiWG0Cq6Bqy
XxN5AR8PbRkiqDz0KqLtXxzQbbVorQ9ixrLnaivpUK1ZmOcSB0INsk37eD5RsSPy
J8iifoM2PubywLq9GQm6QXDPRoRuZjbhxbMpcjC1dLS+6Y4NBEui80iEapwIZ+kj
LGw0T2KTBYSL58nc6zoxDKI6k/UDtOFYm30ZkXT25EQsZ4ZJZ3m1Xldt6h45rjPH
hvP/0Aat8F8lPfB9bos2DKOmzSryyH64nr7dX4AAvnQoSs5XI8InSaCHH2c4+9dV
nz6+yYgLp6SnItyl5CsALA/o+RkaeauF3wGewnzm8qNJsxc5Rejl2LIpn8lHBQC8
A9oW2SFOGkNm9X1XAlNCEu96VTimyUxIZOSe0WJoDM/8FZfdDSIZZkmUbAIfiLpC
wxANax72PlSO1fUV3dF2mNaGye88SS7Pndqp6ex9fYbh/lP9Bz1EgaK9Ta9tEbpO
b3+Ggbc/7n+s35O8PDX6O2mllV1Dotu5kVQPlEDf6r0yVnjZ+IAbXkh32MRKes3Z
ijZ4tWh3NCSrIkTOfUGNP6I0nhDGcBLFjTiEXZWQZdu+hpVjCb+GrZ+YwztvjNv9
qGnpgAnapVew8YEr9j3C25SaA0Zwz6CEcXW/neDco+KWG3K8czLQgFZGRXkJ4B2g
oiuvnCgJRJmx7FXq8lCwrr9/cREHGhhU2wgRyDcYGSLXQy4QpB54bJza8Nu93aAN
lu5s3Dh/8fo/evnTMkO3DU3BwDWgFNMSdgVMIwDKlS0KmT19ICgHJbnJeapmKk71
XZQW7aJamNcFCi2LP3IMgePxeLk5ukEwKWuepQlnjjYAoeqwu7kAhrIG/9Kal9hY
HhX2mCSRzTZZ7WblMQFp333Ewz0G76gIEOvBYyHKntwE6sFC5gL7nVP+TRpPG3Hi
bD64L2LVRhliXVi0Pg3ewwQT6Hqp+tXIGJSiYmf+JOnO4v/EWAnowcsZEnu6zMuO
uy2iWPay0Ik3EKAXSQ8pAwDNTwBymrKfzXRoM0qWmHtttNXTaDsfe2BQrSmEcdOW
/tRw/0M7ACNt6SpfC1tObqvI4ameTNsvC92qwd1S1j63k+virYQZIlF4fKWK0l3k
GpAJ3GGi5Se+R0hJ1CURXHe+QJsqOK65+0fyzjJnb3OZJgvrY3shilkJR3nszhL1
g5NQ7huy3j9Dzi70NEOW8sF83fazcPPC1ehYvXh5/6QE8MJ3AiKUcFT+WgqSCoJC
wjokapQ8NnehycQb8xAhhQlRfvKYAjmX0BgcZoQVRvHOB91GGfJzVCkcQ0K5LFrt
AT5tKIX8RKWVxNnguV5DapCTh2Z9CtmlJxCM/EsryIWgBDOKLo9XFn5hyXckt5e/
koeBTuIbJbTvGuR7SihysMz6u0GaYc6WbnsriLKt9c0BvAA702slhqWe9CLyVDJa
Um8SuiBrDG9Il2dHfNQSr8liDhLEdmr58tKxt7RFre819TJh7A3ON6DiQmk8MIDw
MrBBDlWC8SqUUaMQ02jRcj4x2jvLVN3zjNh+fUnfSHxlBt3WKQcwDljbg82/2GFm
F5bMEisLrd0WUEZ593zW3GSSiBmzbg2sfm1NIMlMLxt0bbt6W4t+InI5dWtx6eOo
ol4L7iB8LOja3o8mYjaATCByDOQaLFyN2aF0UeqJBv7Ls6z/vcvAtJ5ZOmxTcmcv
4kdilUWaqVwC1drvAbo+QqLkMTPDm+CSPapwE7sIYhK4R6vV1/3zmsWk6qyimYfH
U30Mr1OUIAEXEm9kMb3S7AYUK/PQZSb/0s5Bw/vK3PHfndbo8dovPjCMBKewlrS0
ve6wQ8pc/Iu1j7Q2mADpHAOyKYYoYEsT+lQ9J+P1PYeE5gWo7js9GVPb4ryjyzg+
SSQjUhzCjBMQ/GvnUk6vrK1pesCiWbH8cPAjrrzWy4Hs89nGsT9vX/PEMwA15jah
seT2e/XmpNfCxt7ROjsRWLnEIuWmgJlB8gipqmt356XEfqO5dkvpAIJwI8uWO4cx
C6GKZ1GCxC71U1XUU3KdGYAtEmDpoglVaGKt3J6ROVq/+//ObHzC2mT9fmNeBFLx
GCynnkW30LcjgREcq+cQmNQKOdJ76hEelEnuxUdUiPLXRcLskbHotAmFYKrdGx6L
CnudNovGw1HvTnhCDsfTiLo0nVeLKAhMX+wX8gCdnsNyOD5Ws0Lk98Nu+pgu81+Q
CV0nf5O2v2ooYrBbAEY6vTxJajeGMtHtECbOUMiXmZRP2YA2AMXD5mHuo9y4Ia9s
7thmJcCUCXQqZf/rCFSEg2Q7Cl51maaLBs16dA/inQf7a8JGHpDFEoHIXKta4GM8
p1sCb31R02F43PvndDZLMGHNotfmlVTXukeuYda+i8lvTjtMXpyiX31PDVOiUyjq
NggRd/TnzQjrN67863uhyORpuMz+W6MCcxv3epNxgJnmfxFyBk/6hQoWErN8usc+
w5SaQty9893Fvc388/f4dAS88pgrxRQZqZBfRte4Mhxmtjg/N+hGybk84C6Etj2t
SKgMZssjoFdFOwKDBfdMGHXsuLU6bYkrOEvxzKR+vFdIZdvFemAG33dPlxf6X+L5
/GATBwU7d/3os8nHk0+w2yWWN9HpoaB1z+QXSuaU3KY2FGKkndpBVrzF3XGzt1bC
8VR+LB/9m1/9RgUTRzDzvP9IGeSInDY40irogwi7PV3RbdftpYl0c3bUxla7nn8e
NaHi6x7SxjZ1Ri14lDLu6tKzh+H3M/yhN2cw3yE81FvD7MAA2ur/oQYAKm8tf9TC
zLTWDMO8B73sVg9LIMzzlGoyeIH8Ze5HdsNKtwDKVQ1zGtNWewo2pK+zmaOAbe65
U6JlwcZyDOyLp03MN3k3DDJ3DGxJa0b2eSFuHumUJPz8QjDMWa392/8DuI9W1qgH
9SCCglM8demKXhb/mVYsLL9roWvmJ6J6a6Fb+l6OSSxvP/T3ik2cBN8zsQFeKmCq
NUkrkjou8LSGgOtjUPdEA8qmlKwDB3fq/Sv+9iznFTaWSchIVzKLkTSXtLrZ+nhn
q/xDNE6aM+Oh/z41ENGcqWdcNLmsl4v+Oy/sjcZn29gWJbFtW7GN3s3l06dVleQt
sb90Jat3j5UcdUTvS/McvEdI6YrcQF/TkCnf5fatLHbiIhyPU6qz7Gc0zZGRT8Bt
atpOp+2q4h2pZv75VwlyP7mNTTDyTWXO2dTXTIQPX4UinGH89teNlmXQ86nZe/LK
usn4zcwqNsfP9tHXGrNpL2QMezL30Avtzg61hJboNH/U2A6HMsSBrxm12Y6shmEG
pM9eGwPyq6D5+XAndsdhPBBUsEWxRLN+8EhKPx58MsMprsqyKyrq4mOEIafH/5+i
A+r606/rnFAHOMRFcnd9zrHNW2WivTj0p7vTlHtO1LRR4iNVqmTGXltNNVERsJ+z
/hgVtz1NVfqdmg6miSaGCwVdZ1EyKruT48qsUgV5x/nHAALSeJ5cs12FD4zu+/o1
B9tRZfpSanIapLo/nsyZL4DmCythewg8tlpnPVMfokx/q3n/JgbLLJ4holpU3vOS
g9cNU+B6Q/Wl2PWBC9/3UO/RXFrUE3voB6qVMZMA1YLctfAdfo5GQtpJYHOJBr0y
CvKoJJvQ5yl2cqSCu0S/ZN+Ulbh13jf8QZSNpQMgecqLx1LZgHX5xpvWC2QagS/w
cRMMPPPUMYIc4AdEoEDhfXpTEPCIisuq+WSX5thYC6hfKV6waQkFjYS9YfKrPX+M
hFeNlt4fT8ocHl4yk4q/CRCbnutG0O1pc57iIKQ9rXG42s4lA3d02OH4wvw/BM3p
L4mZv6g1WrPdTZxCMRIK6kWarjNYowHRKCD9jnBYDpx1aAnlrXhGNJyqzvOTOUBI
FFqGwDNEv662ALibP1e7KIWtCiPsD9REwtVFv/4/FjalKJfxKDxRm8akIQPXMNh+
uBvle+5bfXVHXx+CBRKYcoPhZ2prDnjLDefB8Haat66LS6R5QVyfSUbT/3jjJ2Rk
/9q/YdENw6+jWb1OWhPfcuWzaiGKdpj43YmnzrxabwLsmO9eAijrSzyZsKql9EfG
AWunIOBBOBc67SLkNiJA3S58SrPL1SsYXsXu4vu3kS+x+YnB7w3odtOvqOUXxO/u
kH5D/hHN5jI3YNZm+jEEROChNHqmV21Ga0UX8XXFEgs6gWYOYwb9zskyEqXtMlaw
g9BFSYjIgfYV5vHrRo4xjYTHcZsbiRmXoSzCaO5Fh3bLY3y81Bsocx962oU9VZY5
bDsvpI+Vanai4gMsNcReCKsrJOY8+a5aYG9E5ORr3imlT1VRhDfu1pbBOf2HqE+d
XB2IEtM+aBAlMPjeo87py+8ttIowFNNO6aG3/e5LFq794C3eSR/PlYCUoPde2okz
2TJk0bQRDXCgDZNOhS2kBp2ouauwnf2avNEiT+49gO55enhx70/e1N0UKrRaAxC1
btB5cMy0JohpnlBino/fRkx64LjjQN1H/MPY31O4Cw/GQ5I4emjISjqC2Gh6o5qm
mItylduqmKAwHVS7vx/+tGOZME19bgbr3DZv+vjz79puYWZmD2g6GRUxIoLo/m5Q
mwBh9lpT+AUSgn5xeNrpNWdqnUZiMujdBXh+zQY+QI+D1Ag8aVazVjlwOqE6Dbsd
e0SSLXy9+/54fgNUEow/SgJf7wsXgzRMNEdZF6o3eKPEG72YMaeXICk+smmaa2Xx
DoTcb0Fff1AVjy7gpQZS1eHnGMIYcv4MI2p0wpL9zD5qqJD9Yk25syS2j2VGHgbF
heL+ngJQ0/i593BfOzrjsPRbCnLeUNyV+vgeSmBMIi0dEIBGqYTV7KbEo9J0JiZG
wkWrsaF/9mZDNSrL0OWiEToVtXTYUepzUo1ZG8JcCcXOzMiGfiG1L0cHZ6v7m7oU
ydI9krTY1OEozbY7YIX9aoqgRXASfi4vbTchUuDlHNaaKQ9IGmwAC+UuYh1FX1XL
jr57wjUsFL5kUJGrjD4EA1ayxGNQGURSGM9e/1KOn14eHYsAop58D2hK6dlJSals
BxGkpm65bVWa/Ci+qX6x2lTdxaxnAUU37t7ofZw7NIEQvM4E6XdTdYqhAgjVtzWE
v4zsBbV+bcw8uXjpdqdtly6M8f4us8iJhlND1gY3zo0POtclHG17EoTxE+9ISML9
BW0iom8UH23gmWDcQnIBa9EV/3N1dGcQAcJGhxCTX/Fi9HIWWSLYdMhgsqDOoXPn
KskUiimqmepNl9FT+jW20Cm7vS+fiVAS+wRxomCuB8cXkc5V6nblZSnTGhIZrxTG
G6nGyIw8xUUuxSqJfRIAUDW6o3MRLofoNLXSJm9C5iEjyWLoUsmLLKKcukZO3hsB
jmeza3ZL5FWDieYig/wu2Ltxktq3kUjMSMfLyU/y6N7z2ZOqPIKQe2++7zTwbWXM
kPqT5wpOM+vXbs4geJUO+8OMKkGgxONhKmuotu8YhJLuCTGFpHOD0DifoBPKLhkN
l9ZcIG9g9cIfOTm2xXg3c99Fv110YX/vVaS5bj1PgFsOfN2UiFyv63Wxc1M8UOiZ
8N83B0Er5XOQgBgv5wUL0JPBXKZToC7lIh5cRZLqztyFujfQaYK481k/N43YEPGD
pmblh9Yi4hvSLFWWLo54gNdcnrvlEiAPKo1N/9AEqEPlNHEc+jz/5uUYjahmucqx
jNyzAdbnsa2+ogGh7T6KT98011OUzw3SaVL4+3UHUd/bwmXHbmmAzxAyI5v/poOP
QmZz8AsYps4/J5Vi0kZnKrLAmRaSmxa0rPgdBhQQ5ivIuslKmB01nF9zogJyNERW
k4gEYZmhGjFrkARikL2XesvHDJWUei/6Am6nMza2xOlrnOh70aYGI44MySR8lrHG
NJUrQv5CEPGbIJqmuX+gis8bbcgRaoH41/EwhnkY/24NU/18LOfmPoScTtCfBv7m
4jB0Q7xeK83gE7x2MqzmNQ01TXBIv9XfHwy6BvKr1+80lI46CLl8Hbe0+KiIpUbg
7ASHQJSCwBxKFPQmme+UoUPWDkr4UCBk7nvYyswQCFRyoW1eYqsDvp6c6acQ5oX6
SJvGIpyTcl3KObVO6c4SgJA5pVquSHt7phsCBo4lEVnggf0KNvcf08RRDZytPyHP
+WAbfnfQJeGbEh8cKu+WmkOhGs44FRQQko5MuCkoSy0Zrk9QhRg/ZijrnKlsJP1V
CChPsYTf7QOJOimL8DFWH2zAfNeZdzapUxjEbeR6x4HpUQoGZoFwLS5A4GpwoLIo
b8qZOln1SZRGnU+n9P0vbGS3BLRp3OaRhHffE6i5zUVoNL6OLNStBoKa46FOwnG5
fOSO/DUO4xRtFdZ9CY16LuJOkUteO8LIqolLaqPZRMu/9k1oOhWxh41WI4YkM8rh
lUirrs3LCVsuhMcERtuS3ptdL8uW8v7kXplQ3O4rF1CEbuU2xW5WRurgnl2AGsPr
lkoEvaGrkM4zuMArlq3ns9EjtM50PxPC97zfOWJZmZjrpX+t3ho7d60OjOTTkHZw
cdJ8Wn4EmguG9ig8rtSK8fcFKlHbu7Lp7v9lhXIHYLQeHBsjOeaDFBp9guEj+x21
+ZSX5eDmo1c1rweAx5mqR1nP0WIVCyo8Q7HUeVT8wQAWNZrOVo4ZzfxFdTXUeG5g
3EbSu9FSzLn3nUcYM1aFT7fe37Q5YdKfa2G0JI7Lr3CVX6yKR+liVYqYUKMH7izv
NqwrrNr2IcWBztS07GeoB3JbIFka+vcSKAiT+aEAiVKpYq/e9glMCJLlUNA1Zyik
KK1clmEhrGvwXbXeky/eAaLXlhGcBFZYeys77/WPOjb4wPyASCxZOxfxByQ+VL3G
9/D3pB6fuie2EAySqBrrqUZNdFPCX2NY4p0xuRJ9/fe47O8/JgZGJO1g5PkfobVJ
Yq5Im4glLpdhuVM2pN2o0+jn7J4HcUHs6PLVFADPJSqv6COHlMBDA5PUxIOErfyc
NJbvdVfTIUfHsdqzu/r8lAfqPggmQSZ5TGJ7DNYPvBCZaM+WHzXzqgND0pygWu5t
qMKjSH2C4yWTBVVCGln6aP9rfFNiypfziwAsmUy15OmKCoD4e7u5HG2FoghXQoLj
5RVOyhWCdq7BBG+DjzRzK7/yzWBxwpzUH8ug4zslBgpXZGHmFraJp8qV6N62Og7i
bloFnsTd+0IZVFNWNW9h3jcOOQ/bakdIUDDfxQs1Ifk4P1S/nMK+h0tFjPqUiKok
OzHtpGnFAO25XlZ9/CiONez4JTQlQYbU3J+2MHcFOw3DtHLMt8WOTlNqHc/PNM8N
0s6L0jxQddTo3uVJtj26Qz9XQl0tKmGlJlgW8Nl30rE/2VplKdyGl9gj+Hqa75A4
uXp4nkigEgIGcDwpWf65z/irWMhJxlhLK2lL5KijpvJdooprUlkbBWjg28yLynbf
zvWaTUl1ZiLzJ/HQs2gWuFV521VYOhjRjr9oqwjTv4vm3AUYQcAQSJUQtOt7cTvv
XrI0NTcS18uRDf9RNd01MJ2/4ftG9A5PhHFmFd0yfi1fI3wGWSJRo9vbkM61QdaO
nwCsnIbI4Mtdh7CcG7zK2sIpKU5RfeIRGwHOFGlXOL0m0VNkeYlyzFV4Tu7PFr/M
l2j4q1uLvb/0iL235gzCBmUMFYyQ6Uw/Xx23qrV/zLGeRpmBk+TgqAizXbtkFARW
AI0aoT3K41Ka+w1wDwEpTTl7432JmMfhzm7FRQ7eiy5hWNtL8TaYXsJ+wk3ra/VL
frdB8DXS3nUI6z1luJHMBZYJbOk3MwLiB/bZoF0UCpurJCm+sebzfEvha/UjPYhu
JV3/HmCLKxPf7pv8XmnNqbchyhSECrYZAsdwb47wDb+MGz0iZ7se5Hy5vBuSPFck
D4gy1w3KpO7qyOAtWxAk0OC2B+ljpUxF0pJblTJ0AqWf/VEE3eSwqvE8l2E+t2Gf
r2lGQCsaA1UB6pduvKchJ6ksJB5BfaOLYo5vr+Dc31Vk0uxoudvjNEauQOsxUJKZ
J8V2kK53uoAQwDteKlexNPRsTiLTBuPAsP+a782vfy9u1ICojn01yxtFPjWAWTN6
ITfvFl57SmrmZFicCqxV60oxY0ifNxh8swua+bO/X8eLbS2skbnFS7WqcKuZb5DG
VgLe7ptFjJVtzPOjdOcS82LbhetbykqadLTznOIuJ1c/I0owKcjKjYU75Jl5pJp7
Bt69JuSTUqalsyAr+WGfv7NPIXbX0fuiGuXW5iQUCyM0ObZ0ZAkZSo5JdiHmRyKK
V3PA5viN/jGrebeNUZL0gsJ5BD8wNFaSNX9gZhZz4tEbDrbKX17XPd6R/JJYcEpg
sIZOoS/3bMNkOGAt1KIEAiCTTe930imWv/loSyZmMgR36igbiEVSXGDhTJ7iskU2
oM6u+YQPOVvJ1atxTJIrHqNv8WVamB6eB0ifBj+BcUWCO6g5FlHahpuHgtukrWcf
HDWT23J97H52wXMEc965s2hkJIFzldJqahPQFqotVooQhV+X0pmZFHQf/3L+U362
KVts1Sit7U7LFldtamL3PRMCt44O1oHHW64JWIu96SYMBuCEXpC6v5L0q7/KR0Rs
vsfSQrrzNTKif9hup2HRFcBElzLlJFAnn/ibq/5bgYWBFj/6uPWTpLmS/RGJqWHC
gjGEXucHfGiJ2/+nh5c7zGLgG8ZeQ/qtWfrDeW2ksymdyKC7nAQP8/6fqw1esVRb
XdwyAVgF9VKUU1dn9SQfSAakwwmPV9qPSNe77m9dkQBBRCwgLGVkfUqS/lH5tgWs
MARtrPhxus0Ov49oKndwkzRBNVq2u9ymGOMfeBNTa+poivNspGKet3X3D0Il5cpQ
5mpYq2Ax6Tzg7EMbPHsYxs/uo6GL/jyuUfA/fcg0tfHcIw6hDXt6Y5K5MCsCojSA
tiSv/VWZRDg0RZCYXW+NO2XNrgkZpFEY7rhoo1ibw5GY6Cy9P8iNv8riOl7FsvCb
PmYftUEPgXQNpsbiPCM2erkv8amnptnOWgzmFBp8Ognu/OILQP9LqmTnR7HS4/nX
5zIwFhYfWLMrykNS7Z5Ibq5XYcOmk6QvBlJ/ZKRgxa0bmeCllJ9E6VEsyVghJRkt
MgSUxPHMxLPwYw6gUUB4ia/xQ30T+/11qY4sko31WO5aDXSpalZUsYjNH++a4lvH
oyUNYY0YQwgfXH2VxtwmUd4FCgeY3E4JJXP3G1aDbvkP6zbHJ7lhdU0Xzi9GKFKp
1k8RJQJcWgT61/h7RJkRwVpxARun73JCnzYRY+MlfbOn3H8HwibonR4sw3xCTkTW
Bxt7i+0s5Oft2WGXtouRlI7XibLySRZZw73A7klsjoZWfhc/2yfJy96wvXhaTdHX
R94KFAc9rci33Nb+/Jo0xiuBas+LqOg2U9bKSF6RjBueE+uzG+rxy034Su87pOH9
QYQc5h5NidEHQiOZLjQl63GL3jjEmUiiy4YtzgXkPWM/JhqpoOUeGC4HcRYgU+cB
1fpN1RaZwbt02MlBnRrJheEZVwQQZ+hDzLBMaZHk5Warz3SgL9EDBK1/iI+3QTBQ
1JqnSefoeldOebZp64wP1sUi7zJI+wLEKkfrdvOU9VafzhHAqt0d60aSlOxVGiYz
P7iP7TDnopvfEyyMEMsmyWxGUKoRWiswdFDCG2o07Ux8LAoGgPJkJc+4LHctdxLW
I6GDBZOmjeQ89G9lt+b7platY2fXEdjBH9ATputshf0YRpx3jvmntuyzfqUcwbm6
6K6+PkXFvBMcCPWqckb0lGSi88PiucIps5Tv13t1/Q/v+WWQzk7RNi/Lenfqv0Pr
xDzYLjGXjoB6uMiMKegTbPVzdf9LDhomY7hOwpaCsu48BQWGYozbWL/17wYPA151
i9EROA787K5me5ThrmhEzT5seXFO1RnuGjydTO+CbJ1nBpHimBU+NvZ6U7FnKW5z
5Ok/oFLPWVvU2Vc5McDi99zItdj48UvXLWssGNIS5W7p+1X7GoMB44GqfRE1Ij2u
hsl0YXjtW/ppGfVZpNES7N7HRk5KvyIfyLWlsQicOxWUynTKW3lpgpWwU+RUX2Yy
L/m1gDzKt79tmQ04t3sxUjdtGc/XZVls07Q6+A7dh+KM4sjLXo7u7erAbzv1gNM6
Dd9q/Iy+1jsoampFchUR4uf9IcvGA4mxOMCwxg5w8pVIyffNnxL9TkL0oqAqhctQ
iO51UYBKzWf8/Vtabwtn3KGt+p2YmDOZ+WlXRMG918DSf0HQ7uzfD54iPrV3+N49
EIZmnHVQg3BNQE/Iu4NRcU2BUMgGcsWZNgIX+rAH/p4N7k6pV4dXDIXzvK83cf70
eb0iFiepEqE8GaUlC8tPQ/fNzqtdxl5cid9j2JY08FiIeJCBOus3L89OZof2dqML
/5NT03WrIIDm9MONolm9x02gtiF4bDTPSXXwKPM1DNyuh+s2ilRyu6EOP6R9bg3s
dTuVuNrDv0kY2a3/06Wc+e8ccIoE5MQfLDpjzcMVvz/2RoTe/CX0Ny1+dZuvdz1L
2zBvBbgE2SVm8IsZUXO8m1808KLJIzZwoktzdDoVQyFa1pxdwGZQfLP+AToac7zm
YkHTIXRY8o5W+//zuDZOGtCm2YQyr2G7ScCBwgAuqJiVOcPODxGOhW/o1YuZjCeB
rAhdE9gfzSKWgIoZ7X9zDNEo9oA/GT0LysFmjIehSdRAdXYyNYuxNiIec7nX6lVB
LTX8YGUQ/gtykcUkopj/fUSgu3AhT0JekJJ4ou6nvIqpVC6YXkpWB4tVCeJCqHC6
GQ/F+mT0CQdRipULaH5fvtT54JxbmLd/x417a8CyocZ5zQ+bVQsoB+UClwWm6RHC
GSlqlqwv2pN43B4JRHGLLgQBgomevElIvW/Yw/fXb4eDuR5/4Mo0cuDtn4TM1FE2
nBCpkqAMxwqR7gkBBcJoUDL6W5t6gqzzuWEixlz8YbRi3FkpsaUH2isMwA/LupLn
NjlwThrpINGnxxdf2J2bE0dNrwRl0cVtywytIKPXNJZhBBlpb2goregCUqH6v9yS
3Mel5XHQ/hg1BBLrlYyeX8cmffONzBTpJOO5KtC0uiX5oLNODFjKsExDmmc5Mycm
tzixnjgV2krfNgO4cgMJ3caRN8kBehd2SjSB6B9luR8cHnznHU/smkLypKJ7wP31
JFK7nWajbLSNVRa09/qHpwhGbN/Pks4zuMocRfh3MXbpnvOSEE2kQLuw8t8s7wau
bQH+xcO06jMUy1pvzYLApr4jCPl38aXfRGR1CKwXfb/MyE3bs1Tfq8dHijfZIc/B
t1OdK/Bnrz/m3VyGnR3MBJ+dhJ79xYe21L2XnpJoLBs50X0eTX10TNlP0s2krjKy
62xmRVZkURpA1LZoMv/GEfiPgyGxc8Wi2F9YMtb6lBhCMmTwCGadBeZtNd3muWlH
UmaD08EIcODRT6zqoz9u5aQHPaM1AD/XU37pMQL/a8QIfs3ftTqopvHIZNBUpP8p
OAPqHwcR53Ba5Hq0HcRsoiqZZ3Yb9/yqYElzi9iUmDrse6ZN9CSN85OtWldzpDxA
GLIuUFggPt5YNIDerIRj/ML8WUEAb+6lFtiU1sd5sXrqtmjob0HlMuHRtfIoz6eg
/pyjFiYn0doXF4A8Tii7KydESdCRI0X+ew/BRIyktPPhQU7Gv9nLKgmDBJioXKQH
UMrRsUo74k1LRG+IuagwOuIp6dNk2kCJX+Xx43yEIqrNs/y980vjp65fiDCaSb26
JVulJemfim/v1PScBLb9B2EHED2zjh7+YOfQQRpicrEL38drtBawFPvaGvXP4rh6
pgdNLlqrkFz5+lvAfVR2xnyikss1R6/nZvWTw3Lb6FR7neezl4WjISlDwk2IYX3/
jlREOgqfb2NMgoH98LBc8KddtUOGcImPHTjq2HeZVfsYN0ugby2zLFIJySUVkhJ+
etb9HIeM3t5FPYhlqqozyzL/7eWdS8ds605Q3RYTSE6mual3TKWwI/9kieKB2GBz
nwTW0oR0mcEbS/LngLRn/q1H+vbIAjIoggXeDuGu4+8wfDiovLN+Xb4cjPC9WZj/
2hKOCP5WTGV6kCYz6Mt4LQZtrHIPowfmFV+rfHfnJWhd0+zFyB3pRsMF/8HHXIM1
JIamLr6ubFnPuNT5inzx98F9OA3UHVPTX0cG4Pbokw//EYMzMxx5jS2vb8Mgxp4/
P+PBRHsWwJ1CTb4Z0p9wJivJ1N5nPpA2jXynunSR9tvwqGS4zfigLI8TdruFiiYu
A9ZbgnT4bQxVIvkbnVSCTcyWLNzxcDMCKO4sDuauFQmpm0xctCuTEc2bAAvHYd/j
UUBrIz5rxsufuOVkrqAD/fdCxe8xzIHRU0i7nCaEa2ONJZ6Hlugo43ln2t4c2uDA
eZJ/9Gdsv6L1c5xG8i5PxOE1d9nIjPotD1sDJjPf+0VSELpuKjgN4prVE8V4o+lI
89kKybt3rBtHEtpXF+oMc0/9HViDYmGFirL+iCMUJvMOW6TGt/0R/XE9GGw3aRgA
QqkFmUlI7hDarK960sfLp38SNjTNja5dZR9D4VnS+A6PiKDF7ntrJel6HaaFitaX
02TqWHq+jkTfeDNGfwQddE2SSO3OXQGnnkT/JifVo5xn36v0qh2f2wNO4lkOlDeQ
1z7/c+oeTly+M/+dmolT5hYS4s3hjVzSi2U+MFAdxZC+aDZwJju/xgZi07X+mQEd
uLyUcupAxgG3t/anyofph2BJZphTsLNhAMUA/TH+AXj/J2yv4bMSbg35eszV7+mD
R6eKIfcRmcBa36FcEtt7GzhPOq6fv3uYoJXYFFqsgA9yoN12/ZlELm63EDuxo8B1
cAKR8KT5KSZJdhN97iNIYXzBB4j0dKcv1yCyFmcoPyWEVEG/AClXsr/vswF9xvlG
4pOBiK4h6ltzqap87nXp4Y+XhnFsJyJG0JVjdLuop8Y41GEg7viCMjxguNFjkNrV
ILtIDppOSEOGnSDZJTlI+ePMK7SIDnIxZSPLl1xAXlWyOSRN5MoAn3Bp0LajuGTe
i9QSP35id6nXaoqhjESyDhjwwjzGIKpqV/HpV+5C3MixfDEXl58ZC75Ky7n6DT8d
iXeGBDfwU6CeqhPparQ4u6mWD0jr5Xsa5rN3gVUwJMTLR0UuCdtuhrn43mq83qz/
lw9ABUhpOZ9XcRjkWXAmqzvcr0hShG16V6zc1RrBYkiUhEuIV/zO8iN1lOwjJfen
ReclRWT90ibqa47Rjv4hsFMRS1U8sSifDNNdftsAr/kPqnSKdecVCvF4Tln6v71p
qLRlNOPM3jTN5L7DK4YLEmRCC9elzSAoRfOTYSofNMv2bwvoMSNdJlwqo/suD09n
JDQRYiPLZ/y1GbEkR6iG8dj9dra9Vxr7T/+zOP23fDOaIDL8VgD4irbzkdMJWeyk
8D9CjP5sPjIxLk8HYcomZkSm1GkwvfRx4an/by4YE+8BHNCWeS4imlOKQtXETVvb
bsynbF28tXNMs9TWLY3+LBurzuunroh9H0ss0/J8W3JgNCE6GTco/XT/p0vsp7uO
gJylQGwNEJ13Um6xBMdAEufNomYR1OoC8l4wREQWoW5FQcThYDFclfRGClO96SCr
qu1x5Cbk6OA4HLBUOWqYxeYLKXZVQTeaCOotifxXQuYv4K6tSewVCuFbCueKk6Db
CbZbU7W1VtrvoGCpbaO3cpqN4uwmiPb/vllFLtUZFvn0Vzji9l1SDpOIfGZZMQEp
I0WXVB53JlP2hXgSLsZsWA3oG5GsDUbJsaW1koYzSFxx9nxLAhZ9+Ow7StPMITrh
Uarhp3yVb4ewerG3/04kqwvsVX3H7XpJBQ9zQlSzcYFiu5QLYW88NnEgZdxX0tc+
N04dtmYZG4re1bD9OhXHE2z/nvJN7AfPNMlEwzkpRHFjWoon6xveoBKbzMt7X7Ro
A7BZfInxRlYKG9QFLS3qu1jDwOIVdZJaq0bFj/oGP9VDicfyAkgcxz1RX6kaNLLG
y2qdfN6+zXK2FLKMKYyrYNZnfCilakT4oq9xuMy86kmJu9ZTlj9FgDW5vU+d32ap
vD05edITq/F28pbBwl9XEtu++Q88suXtgly02Ei+/SGlqmnBBxlaK4SA5DmJjoU3
3tOiF5EyJeVr3N30236LlnXgeOxX/vLXb3fz3lAdDNdBpASjjJyrLVfBkmbesGrR
S87qjM7AskZVBy/XCEL4GKTZOxsVf8/xeB3VibEHw/I3YdFeEhLzrCwcvtA9kB1N
5u3VWLfiRn/KU0Higk6UU9jNtgjV64dFP7L6jzBWzDw8av2WRN5SzZjDPJYkUyJs
bvSGbcw9QqyBSm88Kktb8EMK6hRVbygzF7a9JkaizPCHdHIMaNHJV+K3iCo1c7wJ
TEYIlr0N6aSZFBBPl/eW7mGGfjY9k6oV+oOcdzRKoZV4T7EtI2Z6r0pm7esRfLBs
2ujy/3Z6R3ogFbtg0tqCppInVRrpDCZxJolPrfQ1ATNwifpdS79wRQg7OLB1OYJG
b0sjmqF9KtyhUBZM0/xH6DQemC46tgddaD6N96X6vo3bcSpXl+UkdtGD46/eDkxY
SHU3vtzpYAfyr2AbjlIVwSxP3wnzRL/ztE0GHhG3SWoO8iO+iYULABgvijxHHFPx
nRv59yr6dqnsjAEkXJF2A01Hk26Lj8UUnniTUhPVuBK5kkaCdkSj/BrtyDlfLdZa
e9t4sL5nM6qm0x+JzBPXi7E37dqroM7N+6JJoHfqLyfCybLbYy2lgsvunVwj43fc
Ys4FIZB66Vg8Nbakd+amG6A0UNUUcVERq9e2s6c2YiIXFbLZLD/CU5zQQAi4vaxQ
UYyknwI4Wc20PRnAED95aYLNheaz8XcZvEKh1ZUBVupqMnyzKTkYbnwc2ynYnB5Q
3P0Ts4zu6Gz0OlL1TmrK83WsQVADXmmo6BXzX/LCrPQH89Z87Fa9ptEo44OaiUZp
Y+hCY6ugyXrqlrrOpYj6XR07ouCoC9/FftTBXEImq4ky3UVy9iCIfagTrgZu81Pd
9iW2md5VyxL4JpKtRzinr6HLUFlAiM/ApYGLTiRenq6Jz8EWwmFoV8GTf+JYMTZk
EyXJ6GKg8Ecd/yEb+WRCGNyw29lLHvG4w+/Msrt4BoKNdn4SCarAUnYwYsY0rs2G
Nk6Men/HDAODtqinpezt2EIp1aJLOuusvXuP4sgLMeR4u1anJ5og5Zuj3pr8JEsg
/LMOOtkeaqL0pvicg0Sh12Nz9G+EvEdC21718H6MvP8kIPGIoPbfg+iL+P5w2aFd
q0EZneHkUxfs9o4YLdDUvGRRV5DQCPr2g1+3BDWQnuv3/0/LRF0xxAKMW+niphbF
/MmrKT60g+260dwhO8tqwxfKngIfYna7GoattFmdzap2S2zncaHm8fDgyagOB74f
vlt5zfendZL7JVse7YZpxDCQpcIboBAMSaIV7GR0jV6x5o+BU9Irb4D3ruLnXpiI
10NLlsegaJjY7CeiOkoEj3uwemB69o3+Cx0MNhgr8VZOYygq1LfxgdsY7oDd/76/
H5PCBlqT8fCx+twA7lfHRe1hyjz/C+wrdFizEDi5I0mV0aNG+S5YCrkCVn9PISke
bphmTj5eZ1PWF/haFAhn+yojcQkzaY8jT4+eqgu2WVYTR9W/IkDgrvXTNvR92WQ3
CebQ2RX+eMPyGg7M6yF6Kn2cO89+5vBfv1qntvejqP3uCrQ+UN9J3wAEJ2WXQgiH
6GyXzvjiASzyZDTUfqM4fBGbVj/+ksN1Z0xXsvFVej/Pq0YqyFtu7W0aRfY1KqyO
WYQGoo3H02Z/ti6vqwJFAuJLzPyDRvDJfB8RWpyE/e4HKz3va8jOYahxeIdm2fvq
gY3DNeOKMkEylsQ+wc2g2vvYebn+RNQqh9lKYFrrs9GSW3H3+sAg/wCfTI0+penH
Js8ySi6ZzWp4RgCOnjxlwQwiPGi5RL42jNMhzCK6CPeCOBfXZCBvHbEkg7bQM7Kz
bJU/wwhRdA+5FDKhcVUw7WwiGH9+7+IODMzhsPtj8CteVjkng0hxSV5ViOS3OgAK
FHL8R1vHsNKoaiPZchWDhSD51j4pLzEEcQ4doDYIFbCdI33mk+O6GllGUjwK9soy
148r4KN3OjhaCAHyT8Gz2YCF6mXqkr/gz73x+ZdmjzXUaOafxTWLl1gS063tTeoh
Ctv8krJ45LYkmlgy4bONkEp2aiWsPlau3vo3TkqEJg4p5hF/vCn7INSFlGQXvcNf
NZcr+FVkIyxZ9xbcgBNjYHGBxqhr+4gbP/UJWjSTctzRdg9OodcR6IXIhqT81N6i
cRI173ArmkKYqVe6rFMPyIAiCdtFVuM0R6pe6DsVfn0IzmZ4+EEkyk0xndzAVYaI
LXeVx+LDpGteQ4jCrDpFZYIpOeFL2XoiN+WF5bxS9Oj342q7G5fZ2E49SgU4T6kC
d/fbk1zFl+hlLRaSwBQi2b6KKHJR9483WX4xVJTW86g84/l1G7gvyxA3Mq7aOgQa
Lc9fhDTpEUrSqByn/wFlOOuSbi1tf7rMGt0RxSKkPSunCzkQptcnCplRHcNrGJ6U
LkvbWWazhkkBeBiXc10h8s98SS6AJkJFhdWDAUtEsSF240+UFPHgQpuXsNye5J+K
vuGMolpqAu3Vo/CKm5QEyaLHtuNnABKzT40pxNXwk7Vc6xhJRf7NtqAXYAQNnGo8
wC/v358moiNQIhUr85ImYIqUgEup5VtKNwwxz5hnbbl0HOwr5YjvHfl38Cd2JqrC
aHsLfzfvuEdDkdPScktiekLeZMzP9+GSgswICAeJ8gv4DeJ8EaJAKM/pgTqDBi5h
okIzRhiRnIWMJwxYxymxY6ail2mkP5sHuzkcCgGEDzcWmO09RSx0b+u5HHtMfln3
Hl+0mp+sbI9mzey2qm85Niel47JZ1CGqU3NS3b85jfFaiGEHvbp98kGVcAR5DbyY
VEJQ1WJ8zM3qDgRFSx4JGnD4XeciqtADhLs3JsijfE2RCcVjg18xr01x2VIKoFF8
M1f9lRJEHO9mYctTbmrJw37GHdc9+wmOHTv3B7fuHdWkuBCKo5FAX8JWb5YYnkXx
EHIZls2s8RzCEdHWaSARTIHHTAuVlOecRMsRdFfACMetDXiIObsAWr3nBlziY24g
+SetpondZ5mwD9olh9e82v1darbX4+npwoBUqDjCEVE8zaK2RoH1kHCS/Z94p30W
COyjsaIAAfNMlCuQdmuAa/Rbl7vdSs4nrH3eMRXjqOwdUU4VZ2ZWOf6zQLsVhGL7
mkKpqmE6wZOqeNhD4Dn4oVPHa+MGldVTEsCVp3ivw9w2i+BYSWdVCF7mLmBhyglI
wJUPueVYMK9oXdBjbOfe8PzpYo0jK6htytQafO+b4/8Bnwm5XWgRRQoOA0leUqrz
Oa5sko8CSn1wdDNxFtp7e3ExUQeCSrU1/z1Mh5D6BRs1J8Vg3wP/g9YGEqI0chwQ
rpJif2T4IVUmlUkqwZCnSzPDA5a30TH65bTNuYeghcGm8dM8X47SkrNSJgjZ3VVU
3vqidebLIZlfPJB8ai9SCqs6uuT3rwGDDJRxlpbsDv/euU1me6BAapQ2PnCO8PVa
nxxWfDs0L7qdpXpMuLA6gTZ8jHNivSEjB/cpYpRpAQQJQX9trwQy7zFK2bhGdFIe
BfpqZCYfHSgLQIPvyYfbAhneauTn1uxPMolAf5GEIxmK81uJ0B9Kuj3HVxRfZoS0
X7d6vZJddOLPCo0nO4rAOKPVeYZ6utHZzuWNscltlh7jaJDt1AGtwcgOhlg5Qugq
jvI8N35CAQA9IfkS3PecyryynCjaeIdmT6BgsujaG7Pse81m4ra++l9dnwKda4iD
sUYWGLoP+eNx91BXT/7Tp/p2xW3Mf5q0aH82hCyDmryBEsDg3PByvUQGGJ/hf4gP
VqLMD90MxIFjMplRI8ZImjQiqWctsE1W2NIykfbWaY18W+pWJ2AUwWJwApQ8rRnu
sP1NZEYnBLLbpLky3LOaCds2TREHPo3pZu6wm2qvomrR5bQ036q/rYQdfjXzeVRT
5C4c2NKs+Qcp6edvNHNkxswH5X6mhkklyh9WFVeIyHLOfE3BAMxdkzQkiqZ/0RqW
/n9SaeFBsrBGqd1M9Du0vtbuFd9NXDlqsEKh/vNbVzhB7sJZRAy8uHND5wiL7YN5
ycWSLqE3OV91OP10jXK6ckmF1Am7gqWMBX6uZ9fYnYM1+2fSjpB0xTCT11g7R9mC
SDeCjkUqyz+TLT+l/2PdADgVvoatshekVr+rWw6qpZlyenPA0uQArl2lLeALGBMa
z+SP6CVW22Ct3iMTfXiAgsnJx6yJ0Vj6SXTlF0H+Vj0c6cbrJ8k8ZfbKz/ifDB8n
c+0Y0JoRRLTImgOltGeb2P5OKlZVM63gHJKt2T0kjg9QTRZxiyEnGJufKoaRF2xK
wjTWFDLClme+0Eeq4NXMWxnMqbXlGmQSPm6QyOUyDeDGm8638HULJbrEHBDztQN3
HqxANl4ql1VBn0O2ewdugTGnsp75DG8sEAlxLaDnyjGtwk1FbnVyRsOL+xQhTzQS
I91sdpy8OzN6IvRKaw3OdXjbj65ZiO7pZl2/yC0VRFUC5y6EMtEscsmoHVFfKlXv
duEx/anUjUg7m7lbABODWlfz9+zoWeZwEMPLLXEmNWm2BCu5pB7/tgDiw9nlRzBc
V9Pcn8uwVBVtL8+dHl37imRxhJTjBAFPDNYM2W5Hp9HA9k+MybVEu6rA8HAbPPuE
lFY+8aNHOTbKU+WYkQxjdtI7Wv71yK5OGxJs0kuwLK8vY8j/ods/k8vxAoZJa4lN
/ydml0kgmKf2iKdGYB/L4Lor3O+TZGblMtSO1eUlUxjtXcU4SdEF36fJcHw+W9wq
PiLkc+uW6ZJYtoUVmOX4w3GHVQedYLpRZQV53Pf4mtPtYIMZyqOM/qAc1CamDTPW
Z+O6ZIEPm5aSnPTiiH9Y6z5v9B4g2SOPOE4QJgXnKa6tJHJWnNrlUe7wn0poFB2O
HQjlA5M1gmDVYk3vt8E+ItybK06vlRC60QFmj53LsDVhgxnhxho2Pk8Q0yJ7+rR3
rJ32wT+o01aIywq97lD3j1Y1aWy9pZQ/bAYxkmT9brgI2uInuNptOHy+ug6wL0Kx
BgkzLWwI1GS71o5ReRLLL7AHWmsFPOLrqYqNLwXoZFpssas+t20bso5EEPdphYMM
6+NF17Uy3aXk+rkKTIz6xQOsnDpEN+O4Yaq7SbZUAcW5H/mVf9HYFxcs53GOivKt
08S9Gm4Hf1yYyBCBL6o2tkblGCyaxylMOGNdjd4XVsOkbnEiwJTm+AWBUeoowzcC
6gqhRZZ0+zlY5DZ3hWbW8mRMDDR72MA6XIPKE3ZSq0QFRbRz6Klt57e5+thzt6jT
ztQTogQmeGIUKfFDcGWV0wVJ3/SS/SZAoQbpGC5K7S5Kjec55Y3IGdAOEwOZncqF
5a4FRTZ+idx7ir5w5fNxuiAooTiTCkrKJ/xEfLxqM/cMhjqI7OJKwzLEnvHTk7R2
qR0vVlmKwq0VdqGfAvc9Ce7RzIdG5tE31HCJHf4NKpKePocRUUPB4JiLPUSzuKy8
FgWCTXZ4AN8tQmeVPq7txD1gWuEaXiYpF+k1Hxpa+EXgIg4X4GcPUe4cH9Ju/bnl
JCohT+7qacFWu1EKrUcabYDiLqmg5u64h31j6STsD6TPBorFgf7Ate6vPGLr82EL
++ga1SRLcOykri7C9/UFB3M7WwuW8FK3fT9TqJ34K6w535GK5X9CWnQOVTRj5MOT
quUazaHJSdIGWiKEcoMEsmG89ffOI1MUnXGRfWV2WebyO4crbBE0TSL1VEOJM/l7
AIaTtMKcENW2AOZNuSwHo8L4Su4d5b8dzVnbM5Bkw09ipImLwHJE3vNLOxHLFh5X
DeK9938lJx0InFD9WoM6Z002ocIdg/OkzTMbhg9aFbrSB2X5YNuTiDzxgdB+RTJJ
kkE4bW1gsryf8eLvCBMzXBrjrheJnBF1uvA3DRNIcmgRDa3PQjvPGUyKbBJgUTCr
XrVfPlRdQcYyLpkwjn/r22kVRmh6n+cE1nN6gO0y6EXem7VDYPYlBIc1avJ/MnU1
azMhJUgGAWAkdY3+W4ouNflgETJn25Gv5+vO5rMecjW466Um+E0aFEteWALTSIKJ
1WMtHIMOknU6ViHOmyHi8RjXyQIxsvjJFxXF/xAVpwYUEVtGyKLMwydDGBI1gw3k
PqnIq2D3L59teUTfGDuS4Z54pwRAtYciYImkX5V5M4VFjnyO4Qkb1Hnf54n32+3E
gP6ivR3eSLAeyvkpOGmGI8s1ZoiHRWSriW0t+qejBz35Jd2k1DPHSU9DodaXKQgY
Qh52gWia07zNHBiKd6NM+p9sEJZa7BjNX+vkWnQ2W1gB/7CHfaqjZkx1PkiwnGCq
q0Jm3plF1W6uc/k7jbuf9UlFEftk3TesGwcnqp65JSmge+MDx4pdd/l1s95kRZv8
U4LNhlXUPaRUb5zFPcqvqww1/TED2EmjPmE1/H3V99zsX2xDjbOjqyoH94pAz8NE
D6enPmg+pXp/wcbEr0h8aCKMQjbDtYavxVbB8cI5SAyXmlwdb24acFgz0rB1vJwK
eZvU/qCUVnp4y/7FguYxOxfl15GlJ+Ghmf1QKb0r68kVNAfLfo7iyf86nGojF3/c
4j6zNN9qODj/jwgWgiQhcn7qkGZcziQQA1LZnug5bwdZacja3Vp5d3/VKfOKUncA
qG40R/Dk112AxkwkPLqtzqAq1qMHH6Cpu51ibi4QAsfUtiGU3iOe3SShMwpn+h5P
JFMq3PB3w2CZ2MJXf3aUUex9YWiesjo+nIThnS+Xj8lhsQcK4hKLnq8EDySCMySH
/ZtDDpEor9UxulBCK4dTkvS4/e63OSEs4So0LP6eI02NTk9b/mmLW/3u0YR1/kd0
zSIrfaMdOBdxOxSoJZDa6kUN9QUq6w1lC0eo/HYlZRaXbU64ttlOb996ndPb/Mhu
2OBDSdW9EsezECjLrXlffzaVIa2mdwrLwsPJ53FphTd1x4ftR78P+VWJDePodBWv
hKy5i3UxelxVkbqAVSpJxTesFQ2Vv8LfY5bXN84ElROl4InuBh6z/BzlUH6SRDJR
wh60ISCpB2NfWfNcnwSlrdk0fKbq39OwPGkth/+kiTe5IZokRE2I2ugv9WruFVTh
gd7ZJHO9PP7LxjfasBdY4UUvA3th07K6GpaMOKKf6l8PoHnmwZzqaSBcDVDqyZLm
jPGNAY9dM4Nk9KL9V2wtp4cKBFMclxSsivZKWP15gpWhwC62GEL/xyzR5mwbmCPi
6g2YvkUAbEtQcAkbJ1YCPcqyfm6GE7YT27JGgDlDTZhUnIrTaDZMkUBJ0IGqcf0I
GSmkmwUHkXcXfZsTxe9eoH+nG1d7DPyvBZxiDbA0FIR/95P1YnNiX1lqYlyWwzBc
mOnAvshHYU4y18hfsWTXy5/nsgjZDA7KGoTKEC7GLldz5uQfpgoVEi9yYkWFDQBy
bUw4mlZs/WOXC9lWKkulLeOibt2McHueRNjHgAbYve6hwvOtN6l+vdtDtiQZSOKt
6XzgCioPk3+wwYcqhE45m7w0Rhajl+jBMXW4EFn59bTKeSg4m2Nc693APBHFhi0X
DSjlKEbDd722vACTu83M5jTxQbQ3Z0vwoIzXS9rMxd8cO0Sh5O+fObhw0lmgAyrW
PhmU43YCELC+83aiSvxYBVM85qjiRjd9J7pf7Y2uARc/whpJsVFDx+V6o+HHkYQh
M1l1CmNyk6x5JayP7Xm4LgJG+hPTx7meBfG6m02igknZHavCkmC8vA7pQ7iaS4yx
7NU7SYBz/VKLMK+2xNOLz3cIzko7Rt7GFUKylVg5+AyDHNCFETDBxA7zwJKg8m6s
nDLc0Gj8np3bjCryhuiHfsTCM6Cc/dnm+RLXIt70zvCKI/jnPuxWsxF4uyoJZvXC
Zs5KvipLLZONGCJICjC4ncAU7noKCGyQHDellIn3peQDeEJLwY5dXVbFhjbwaCm8
OipVOlKTRsdUCoJXnkv9IgPs8lC3jmPII2559FHG0MWvI+RFTMZvgHa5seyLsajE
z60znWDNjzXXwKnpD7uI4WmhYgiSM9sxxm+u3BsA+wWAmHYOjhS5GY/okKc1nsUu
dcC380yAe6JZ58oWtJUkSgASPho8VDqkjpxt2Fet0mBGgiZNt+ES025cVIft+EQq
Z7Dmj9hiv4kqLDU5NjbrIFpP4CbpGttpbKfxk+hrJX1EcnzGJnGuylf+Xn1pvIB+
/b9LU4XXvVCFtvgRaXJeDnpwUymXsDVNsOv+Vvf2eDCFpQ2OKUFLXNTpXSm9VO/s
gjsxifldIfRuZNcS0ND21uSTH/YInI4aLJb0Cz4kFQeCs1SEybV2QD8zyuY45fRv
RiZtGlwKwpl+QfRNj+33gchbzDz/JfVAm054KS7NUoOIOe0dBRAreIYKL9i9lwOy
XmsqKuAzZ4eEfdcyJODJEZ9D77QeMa2i39UPyBdMxhxWMtjY1WATns3LErPukn/X
iDlrOHipi/Bt0yaURe3004nvLLGaJ9C5xN7GV7gG5naQ3ZsKzRGIEaVh9XmuAUBq
wzpaSn3nhwTaY+GBV8P7OQl9DevZX9aX5bTGli5Pp3FJAgzMIMKBIL/W/wEo28YE
HxE4RJcmDhd1JCXiSP5VydwEEP++OAIiTAQmQvupa9hUwjJpXOgu2voQcK4LcpxS
3ZM9bbChbzgkNDFL0XEOVQ0VKkiBo1SDgHpQOACxH+G5yb0wULvu8tl6zYn4oZDw
tlfSxx6SkByIPKj0whtn+MvyueVm52pPAWbrBgE6LHnQwAilCfKgLaozM18jyieD
ZmFMYDf5RhOAnabZlVfZS4cA8BPjYiMwhV7OEHQKhLVBdKmrnjehGLEeCHSrBiD+
CrfCQkWRhh4y2ywCHdos4s4KZdPbbSqeMb4LSs29/V4wPjIS2h7zTCNRkk5Nz5HK
6O2UVXPEz54XWqpR/hRr0XyUoNr1jHUpz+CLFA2GxBRsACxC2h+unRibeLsqM5zp
43kObgDDHKqPr7f0DZ0u8n7u9xZ4vEKt+HxNFxM2p0n1uC+IRDXqfs0mlSOtKEKn
qni+5qAPEX+Zfy0wH6GLAbqTpUCs8vMOR0+YZ/U3gIS2sz9Thw1erzhCrOAVYMjd
IFN0AAtOI9LPuBfmnUxovd/RtAAaXCefLrH7Rg92+o508as29dhIl09eib/x2hVT
Kmzpg1l12VpTwW6pNPsxjxiEqDd5pmuEYDfBGkF99E09BzoHxVoAjQcGLFTUm9wS
hhuU8IepbA6HGURoNvQfAS6kw3N16nWPCu4/5lgxG/mIUDsPSIfb9D2eRHhtcpLj
TMB+X810uiuwLoL9xSmJLiUkGyHlePWfQu1jfVwu+jZJjzXSrbobrLVg3z8J/yoh
mYGFFyzjakJDyakYAWRUJELnqX1Cj3w1zInK5T7ZgSCd6NfweQk68YtFSK6bjJCw
RaEUE5Czji/ds7rRjQMsMqLuo1Jkx5vVJcDZ5IqqpeXEDCt5eRMnoFkHv3KH+WGy
Yz/PnE1onT9IUJjbPrgSLeNF4HMYCMvwG8yxwy9yUn6YlzfycxOvBvqo/VsomJbD
vReGLyWRd6hKN37esSTJfrcag2rlVCsxAtk2UsPZrfCQg2PBkQMFul1TSczhcbt1
BwwCAwXE495wpMiAzAgxEyw01qcFCxY8Y5pt3/HVrbvrlpVgEY2xWGlyP2sND64v
4DEenncC8X6rJe2Pp4Y/WrmI5s2IBvB5r57lEXBW/B8WOCypJtIYLeFRp08arA4m
WTkZCOptMXz2FkT96R5Sc9xbzpqsZxzJ86jzQM4inSG3d3plgI52wBkVBgt6EdPR
1cc+RRaRw5hIxfiKAbH2h0aU95MSTBUgNltrmq5MylyoVoXpASxPRsU7rL785znQ
vBqhFXoOjU0KkYaw3PngIUiSInUzS90T01JlQVoN5D4Q4GB7n12RoPzWdtpbWXf3
RDh3eMCgLiBG9QenUIn3JWbPyk2kiUnTD5Jf1KRbu5rXo3OmCGMpvW8ZF4dEWdlW
LKNmx2VU92uAZ7DPBXzLDznys52BKE9qnFdZUt0O6m19rsSCl807nLLEZ/pzhtmp
7GMqq9uYrJ3Y/8rPZv+K7qpeaMoPZQ1oO5D+5MqS1C/WkNLfkzAmZDO5+U+LgRPs
BKFRt+9mIxqsFZi83RvVERJ6/fh9OlAWWPEScBkAUwRvrSngjFBIVQs9nES+IV4n
V9KkqyZXZntz2ow70BJ061La9zZ4/gfQuiTr73A7bkr4JG7WLYke2jVmEENKWM7O
csT2XRXHOnleru5REnZ0AH14yc8Ov3n/FRrDiiPxGO6Xwp+oX59LZkVZHaT19qbS
jhycJcKDBlgqjkxR1jVcb7gdwbCeW/05/AKpS9WOxMdJQJS8Ea2iu0irOXSAWqWM
goEeRla67EYmfcpTzrqQs5W13oZ3Hg71LT4eF9PDKJrer0byWFOr+tPXSllSMMxr
juJ07J0sRIta68nUQn4Ls8ng19kW7l/uGeDfgWf3j2vT5nPuWAv4SZizubKJY6VL
9Ci+XUBwJlyz5r1nPcR2U8/SmOe171lQsgaz7N8qk84DBTVo4e0UpMJERp9OzP3X
L1tXL9VXgZlsHrJEJR3RNltC5+IjZNrCGWPM4TSLCyNDMTthlrHWcHCSbSVPrHYk
WiSVO4gNRTKjfq+CJ2uEKhBHjTyqVlDrGLNBhARGHZFOlo2Izx0nJ7hzfRxjV1XF
ittKT8hGUYeSDYdXq79ew5YxopgLw5+6tlPxAVoELyJfzJwFmcOtFgBEZlpA91sY
YINv2ouBjIe84j/9+AtgvhNbbgA/Gee/2ax+GLQr0oqQqXF/cxMbfNBi/FhASG/8
/09U2AK/rtNy9FXLfKlJCqYi2a7VANn/EdZsTpYinpK7TBpQgTfH/Xq5MvfS7lBK
bIBKu1yd8R2H5woBp6nK8sBclChbwoQ4MPCf+nQUS69fxcPUI3yuInn38qVLawv+
iQlz0IlnftaL44n55Gzf8Om95wVg0U+/GpL5B9akHAGMEzY68tuImXxYQDdxg8X4
NcXpuyyPCXx0mlccH/pjB/b/QfBpCbFN6kIkKkGvUzj0kOsTOg+olcZW5pQn7Vk3
QccqLizIF7QMwO8te4COTCCAdUI31eCRIAZs2X5qr0NW+5Ujip1qZZKQQnz1LPFz
SVAF9qB+zVM4CgGk+aGcsFBenrsA7wtCQ06rfb2PYij+Q7oEXGQEdScWX+caMYeq
qilJ9wUMzejCMLrJu9TLAaBVP/ImUsbeaMPsl8N6O6Id1uYcMIYSyHORonyJ4MON
AZBoFqoZgiP0SXTSWk3OI1l9FMNpiVQMjfgVHOGQgNLe5TTuQg86sbcR8mjGmP8w
x2B+YSuEM2k0nYRjdjNeOfh/s7qb2ITVJNJyz/H9YVkSZKxV2D26nYDHjUzjRpWw
ibH17fhtbiJfGP/uowTriiJsGMcJgl3QjbuKEN9FGaH7vpTHP0b1xTqZi7C2Zteq
dj21J3cqe5CknhLlrXGe1bmyuTG910/t9H87ubY8T7TT3+nkJDQyfwYvcOVdldsu
R56mEQkKxvXdghc0y8WbVen8vkuPRiM5GJp7UPsr3l1J11r26Haib6aaH9aUFKV+
1raxCTYCqe+CsKXbvJtPNI5R5vpi2OxfP5Uxr0gkApuqhOl3qzOaqPqO5SR4Yrdr
FZQhGfgC1GHJ1a2IMQgrtxXbx+wr26f5Tltvfn++eM2FJY5YC/JeDip+CcrOgV/3
DMpfmhYQzSQ66nT+ZKv5oCapRnEpS8TGh2RqV3vaNfImlHTCmNXhZMwhtTlOzjvI
6ynb0g6WVG/xXucY842lM9LzoYtyUuqHdl1u8bOl1oh7HEkD+iRkYk2WWCjyQ9u3
IV0Hklmh48cquDHyCo3DeFVQBSBpS0txC1Re7D0wGgdMBQW94zDpm3Syp1uhLK8A
sZ2WiB6gQ/zfh6Eop7uKlsIN/r9bdFrjkdTErbd/4vULwfdVZRVSVrBsjSob1bbq
9D1rlG9WVG/L/XTpbEuDzLmOS9o3cAAJhpf92XwecER3XfNqDT3zA+nVV+51GyCZ
GCuWhv1PF2nLgYOMidaMBEPgAAmgJ+uBkD7GaBNHir7CiZA+mjKd6zFKf533Ipd1
fSCAnG4H5/BhSzma34ttjNHfDPrIfYdcTedZT7FFNyoUNvRMHAcEHY9ZoLX1UFJS
Q4Fs9jIsycLCCU0nyCDbNSCjdb1npWZk0lQzYDLNhp8z1EIZtJNS8dhAS+VYS3FN
a/A2fbyJpJTspelDazWxcGN1GG6ttmeneQ2O3wjOWq1XMHIsEwBtvJ/JVXCnOPIF
2773nWdc5Rc3CqRBXh2SdfAkL6vykbsA3Jco7NwFyPm4/TNC54GJnBYY3B+scO3/
+E9r0TI+b7f+qWG6GnU9Y6Oh1SA1zCMbsDpAikxGyS5HfI/dSqaT3sGfRnK/si6L
UnKSS2YJ91950KqtI/VQt6wGAmQzI2R7YG1nWbsqWmZ5G8iyG9nzDZOlGxPRMhSa
U4PVxJ4Z3RRYjHrgqb8eZ6bUwGUPtuAajpsDA2RWK7Cqm84Wh0GsGGVSKR+DAhWt
1aJA8Qkz54/Kf9UvQvFc5OMYlP4ujd2rCx8Kj4OfpkhteGwtAMRviPdjPH1YZI0y
l1EUToCICDO5CYn98ex7lBXwM0eykxP9xnTBfatJai4kwS9cP2YC7P55ScdWWCyU
6KFaauLzqut/BQ+Y2qvFcTIFC/3bFwvM8yiHqNUErFcwexD3W6TzHrY0y4K/zYkL
GZWHvjTsRfVVqcS2MMqFkM6fbpPkQETLGyhy58t+6xVr8Uw4PBxGPeALPdtn0bNC
GfBozfSTsQ0Msrc+s+qe9jtdUWRGMAb9UtKGc9JWF1cs1tXSD8LBXll5cjH4fcX/
E2PbTorF0hAasjiGENbz1ZxCYKdj7b6eTEXpsxgaufQOpM85ZvwdVr8AV/NEpgk9
DdB/1vazvVZndbo8p+0exe1ttmzL8lgOx66pHA421rN4M5Qo+2LZEu1/ygMhvlsC
xYDws77TfimYqQ0CCNVoqGaVrybKaVyTv65ytXM3ND95qUrOICbCyZFGvsVlhAZl
QTeMJLPZ02Mg1/lyUqmSfKYWFmHeUYGYicItGXi4pu6A184wxDxZ+WK/iKKUzpuS
Xy0HGLJxTRPTqBbPBfWLXASEG6JZjihTOWSPCOt7jgvlvBMVde+e2BES2240gETV
X6aq0AhnNqs4DxQPKBfvYFpNUAhk6NkJGucXUxSR8Qsf/RckUdQ5CmCOCsaFC/nx
gzHaV2MtX1fOoRd0bfV9ltQx6wyQ9uMkQU+PJw7HOgJezLdjJW0EI50P19KJygUC
XW/j6+EGIBWkz18Z+9aFkEearo5YXjRxi77mK42YsPrI5MpUx9OpVzBGbqGUCvGi
8oXEuxcv1uSifDHnfU7QLWSuOtCpu+x4TpqqcMbRWvybhcIpPpGyKiGFdubTlGNO
o15muYAQMPUoH9jL8fg9xKaXX88E+rL+xWJqBQh24YK6DFJAighf+ZF4TPyYet79
JGXY9hAI1tMzHFiuCLBomTq5o8MYWx0X7poRjgauhsljomjDwJkBArprTgznHilv
OE0Jbk7JoCJbuvcBmyULjkvUMOdBblcKvW2nmtt7A5jgNBpGb+DiQCODy3JNbhT+
Qjyb2ZFdEI2zCLKYT1qz19c3KZs8ZiDJ3CUEE/u2CmeMjQvQu1fpUgWueFkp99/7
gNJ6QL4KNHnNqoIr5ldDDTzOT98miErLUau9VHDaPeKvS13/0vNn3/MP3zidc7UQ
wSWCcMWslRuA1/nOnI4h/u3cKNVejvgQRfrrsb9ZzgEdTkboatAo65biOgAksAAN
A3bSlp/GKBjnwecBc4VBQDcZqv+/cw16YQZOWJr3WrZgWfuO0HQA+0gDdxYcytFh
j4SLZjE6OHbuEFTA7IaqTT22c7x/UglRaDe84tGcnt4znndlnMfJR1gfLGSimfXR
y89ASB8rgmThx+sC4DGxSw+N3b5tRk3Q6JfyNwPIthNO0CxHgqd5G8mIcQG2wswl
n9/82ms6wkdlZDFPSct3LIXlxJNuOqlPMUv8vyuxPFBdyLc+3iF7GUaAk1sm4c3I
AimCDj4ei5jM36+2IhhZcyNtxN9q0+yFDxDHUqxZvwOYINRr/m2VoAtrCvzHjrgE
9120QEtexW1fb1nqxSXhoqku/2PI0ahO4vLWm2QbCcRQh0Qjwp5/OVcDXLy5LOw6
6Fqgu69loNex7VT6H6raHT7gjlyzKOsIRpEFtV39l81yEICmemL3cDW7qB8PXq6+
LqWXsgfznau/MWvtpCzXKz6aMHKliOHNJaCQeG1D0O20X/P2aowOAd3y3H61SmZG
uOViXyA99XKCdldWz7sUFJAi4FQU4JGIH6mUX7DpNiMaM+AAXM81LogWmFKkrQAP
CzS1Cq9Sw9lo+bV9stF486H6rtrrazQTffaSi+f5sa8aCB0QU9B6dDFrc+tbnO/i
sRQy9w/pqy1W3PKMYwxe4qWcRQkgtOnB/XysJfakrtSbave0H9VoudHQj2WSM9jA
RHlbc4VlMUyjidHXvlooD5alX4Z4x1SGc2vstLX3Hwdev7mirkmoV5CgO5AogWWf
166Hwf+80Ac+HApNmllJeuRwZsp5ac9i6sz1FTKiN5n0+YpT8NpNC5WCcXzarg1W
eFIBi0pyH37ACyFbg5g+5IsGeqU3BbNTMHHPMsu6ZqKJNq0gkUdYKhEQL/w3ldI4
yKOUv03zcZLyVBUj/w642f+FTiQbUyPBZ3aCkLlfiYlPIK+SAPNgh6DKFu2CW1oW
bractyrc9ClXInZGHWXm76cz3V8+J2n5YvKyNj1YV1+tVqhYXpyx8MtuaIJ+tfLM
UkRYSyIb+Zp8w2t8M3rnl2+7aZcD4sN6rjMl9sWRNKRv/usLowIrKAF4jI6I7ZmK
9ssVA4zxxsXrQiPit4iHuB7g98RmoLjGZudpdb4VF+PGa1doUZqt02oPJJiQBDuf
75jNDb5FuYi4odK3F3tv1sB/Od8L2dQPHAac4KntQr3tiqB9/ikPod8aLT8L5l0A
tT7wER1XdgOkTanqGmaCkYb+zqXMrbAyD/tHFH7XvPGjj0XE/j9sYG9s1A44Zaea
RJH4qOvgdVo+p4G2go3ZZBV7nXoVZalpok+9ayqZIhGuGS/wPX/jqEMWChioNMjD
asuD7UMlEwNlzPneVq3a+s4cBpz1FFMQElK+wpNpCVpnpyRwSNM5q8+VjfowPyH1
uE1BQAhloWH3SDlfO2tHUcRiO3wbUuaOQuYJz5/NUzMFfy0yXluIoR57waIbpPGe
Cl7umap+vB0BLXg5zxzQdOzlphGPYwZNSlmGVsHsJiDyqYG92EhaH0dIewNY0dJ9
NKYUJPcXgYrZYrkV3Dza+N/zHY74TH/z5DynULYVopX9ICclAViL7kAVOWXfhz8e
d/CDIJK1+IYnSFVI5DV5N1AWrI+RuULAP0BSCIS6d0VGuAbLSCN7L+k9JQEoqRmI
YNYFPyyP/uOfe2cFLWeJ3i666DPV6HGVLf/knEuda9JBpJhNbNloHJAnwcz1HWaw
PIGlKT+oTS7C3B5i0k9DKB9d1lR8elJzjmP7WtN9R9vT7Vb8YIjH/NffGaeetwMQ
9trnBEtQr7ugnQWSDeMVh89+Z4zQVc1fa6ARtOotcH9Yyf1bfZ2HaP220RbNoxsf
Zh5SzZ4hEOUuo4gjcL5wb8uRGOmLI9IOY7MOj1C6Edna9yD9MwNtR08hMDG/rASF
b2NgCgs4tuRn6bCmsJCeJKDcVI9wnQHWDNeTVkKitHYcTjyWeh4yjNoE9nIsmRUj
sHkgeka3ch0KiVqL0WF2lOb56fs5er13WOrgesdDCaFY6Mo9dWDxJPKi1GVy3xOa
valjiwWhxjCm+HBBj/HPLY+zjDZQ6AOVF6ru6HPZf1PHSES4cWAtrtv25b1FU02V
PqV3raaq8dhvmNOW79NB3wLrwE8KSq3EWsnQ6S7FyFIKxLep9tsO0CRTvBirGbKn
jNWWHGBWt1UISQJAokkqNQlnO/TpxJwlqnNYVJMC7nowB7114U9uJ72zxympcez5
eh6PHgIIlvcDndg/DglrE4LKgUK7xfNtGKTNR448UdYuSvJXZBjULFsn88+Lg67p
cjaNbQsRKJJriRGurweDAtCOggmdyS5ctY5lcrduZl5QG88f5zn9hnckpFedRpit
OLDNfwre7w6gX+monWsjiyxw8PRxhAmk5jfRRYArbCTUNqqrA6oo32fi3Yhq1sKz
YfSGDWQcoMlxoR7jWdrH//+fnbDGiGHqLRlbDKYMAkEz1pezWVi1gFV4hbpZi+aJ
fPOt2XpdTA4YnXjnApJ9G6/S/HJ2qVBZck8Z3/LtMMjuT0c3L6FfxGjuA7p5eneb
DkkwbVaSNT4P/mDnDoL890EPI9AXrDRAvljz2Va53sZ7ocM6nuh8G9KZ4AnPqNIi
ja4zYkaw4gvoLOcckt6DUmMIhuyS1JDY3KsaN5NaS1W2MZOX5RAH07/DnnsmDG/z
T3qOsknms8404XoSCpj3o30FaLZJhybIdTF0bhHbTB9LVUCYQDPyMYNeDqjslU48
Np+vbm5HUI2tlQvF56D9G2/2uQ7Xcn4vomUazgqOgf4uAs1VucwEWrZS2MefKfwn
l9TKhl3eXXgzGgCUtAqyjI472fYDL8QR73eoUUjJ3ch1Lt8W35m/J79AY9rL6ScN
pig1oMrp/E0D5Nctw+7uOCecU8syEl4BdXqDg2qAEq528HFHbGfulFkYhLffD0e8
NoiZ7N3a4v56bN4oG8Lip2ClqvvctSLbJRSR6uoconhhp130LvlIFkcISSVw2Ds2
WU34H4Xg4qt091QBIO2Yvymjl9T7QtjQ2VjCERyT2srd9uZp/klAmw0lEKtyftQ8
+xc2fLNjIc3o6dGoFOr0jwRk43BhXfHaeqxlyQwE7NeFajKtUNBKBjUTEc1TYVZl
8WLOr7pPTjGFiwdAqIXRJpl1q7038Ezq+Btmb8Sb6aO+IO6YSmF3XrG6eUstNoBi
0b2FNIt5pxMjUGEmHbXRlHehXmmLkOATAp7qkT0FvUsaQijs5oBrYgVxNhtolxQe
KlpJ+Y0kjENJXn26i0sTMGh0EaqM+g3xNg7I9kCJwiJYKQpDm7vWyI6rCIX9XCq/
fPA+x5Qqb+JxrRWv5Kr3rcSAZg0E7/mhmK6Gdi+p/2Ugra+EE45GjBTodnTKciuW
K24BrdiII8DNUhjH+/1O3sw91tuX5oVIQNLkTFA9CHcmhsFZJaIwP2/0iyNTcyKP
tbVbZ5xsflM+7r+PikzyF1qOHsUWD9OeGw8v+r3kbSQOHPHuFjMojZUng4sGhJHx
+BGQ+6cmcI45V/MDLnkeNGVxtO4mvQZVRdjuo+PTK4vVBU/5PI4NIDeIU+0rZ30n
G8bqlw5gEw6T8oLO7imXy/cv4QI1c+m8TOT/ytBH17Jv7/RD1d5QGEkxFk/upLNh
opVyUkJO68HZMlqKD2z1M1MvIPpDkrlyaULb+++NcFSOBnApSN81sIzXGfhrChGh
WstJXAnFUPBoU7lnlu2SZj9gm12R1E6vVunEv5H5UaL2dlZsEAAz3NjuShJ+A63B
48cD12apEw3Pe0HoOUljddBJ5wdS9tvDPPRwIAcKnFxg3gy3gtIIg+OmOeWVhT0p
/QPvWpoM6gmf8zJHUzH4dNQeibBCk3sKcj1929JeRhS3mdIyl3sGrXetFlveVAEe
U1ePmaKH8LliO/KXHRP3D7vpEH28Hr8RoGvaicKGD+YlQwNdHMJPaFjxR0RMGPdW
SO9mF4C90WwNBrJgyBXdF37UybRKXewrWQmgFPeURXNU+aFQ4ziDRiJiJ7OcwBUf
kwRUGhKLuWJoFfK9lAQXglQ9+Fqibstml/o0sFBJk97z9Z6gLZ3y7UQW6SSzp/vA
ZYf3Lv+GIYowA4bZHsc5bsUyMQVOwYRbnnL270p/aegHEKjLCCtKhMQdv2R2KJXB
GZ+lKplzbKenoaEaIjw0pPyA9u6J72kEqId3yeiYoG5f1RL/xgC4VLSl6BBMFWXB
FaiB+ARyghzSSsIuepibqC1ZQXidaMB/kBOSb1E0e3sezSrLuYtnAnTWAdW9a1Xf
WJG7ZX3IHRSag3wzzsV2FGl8eRtn02MX7V2VQlBpURpRy14eO6XE7XEB/20zZZ4g
JvyVXWHiOyOCP3Rj13N14LHcczeon9+8HNb0rme2e6DaLZ7uwuZwznOnFdJ0IIJt
P6k11V3kk6WI7qyIt+Gl+7dYbcW2QfSdw+ErV84RBGPEp0U1iqwOJjxisGMXg6go
XMdrcuocCQNcHNP/XIIZma+vuTe5NVTGfIJVq/Bf/PUWI5BctqvdfJPCURvzTVYG
ArLk9XfmHAoa9eZAQXdlPnJ22oTRVD58nuasdz6cIg2xsafnpINEFk15gSM6r0TG
Y8jUp50BYasLwot9Ai7OozXfDr8xsXY8e6Y0Fi+uDIBt2F+3+fhft8MHgZyT0Ofr
EOe0tAc/zavVzUl3HZzJLvM7lGfTK93We5J/fpg57uVAl/K4gWnQi2DCummRvovn
yFf3A5B/oKaC724SOWgL85LX0eiyztxzNlGxSgz7mxnSiJBWi/9yeU0vi9sEUM6k
BjvnmZOYJKUvmOTSRhxO6vEyAhqxBTD2a/9eMegHHMdbMHs3Vqw9iCesZElZskfM
gK5Rz5lrUzH9fCPxN+qCWw35Qou/IfBUB5sUpJZQDVtfPV2DYYb/+4mWu9XcC/Kk
BD6O0eYrhbI+3Mo5RQiz+Vj9lZJPkgMT1bVYbxqYi0R9wVEyYT9cxGl0VUWrUptR
ZkqMLDT2z/dvuh7I9x6BK/cBt/CzDlgEkwFw3NhQSNtrW75qfWIRrDW8mTbtrTNH
fPIywRQVO0IJu4VoTVC5b4kklaK+TiPAZPEcmY9v/E/K92ePCvxsiaWXLUdxjry1
dPTwNKhtfcyUPrfEl+ssF3Wu2/exTCF2HpuALIpKe0+KldMjR3sBwnWDlJvwkIr5
a/qOSe2teqYQ/NN5wV1KP7sNNq4ApxLiE0SW3HB/eKUNPrdDNjDeBU7vquL+d3HH
61eMy/jJfeDkpoqmik8c2XMfbIbZGxLz6GipKWcOGqexvXEIt9mnuZ91beEVOXQx
+flEy50edS0xvQZi7TAn+vPoybxl0A6KJ3CV4AG8xRIQtf4JXRDlM0KTbQ1ycgzp
TPauKChryN4BNmqrilbbvFlMeTIBq1iBBDpPfLPYjhjk855nN2JttuzZ+aQQ7Lei
vwuG6A5jF7yjLJxgGI5fpJh9Pth+olQXgfGs74oxh9TsWuCdZDpVknImqkcIuSx7
VYO7VLvWswka7QOCmhUG+B30CXVabH1/EHqU4KchdaI45hj4tGi4uqBmbys4snxb
t5opxtxRM3b8wwDaXrmpUZj8pE2uCdFJHujnMGuPdylIc6rlv5lYu4YEoL8arSHx
Ro2GIYo5QW4zEfX3JCT1hszCUuUqQ5374CHI8Lvc5R3m5Q5mpLSQ706gm0OhRpO7
zJxQWsR6mMV3jgfrc+6gs7gj8JX6M2iIrsvZwbfLaZzsxEFCGsbU6pkv1/I4t+TP
CxJ6hnLevm7ukeqbaCwZozgj6OCk9MKBopfELblalsTd0dJvab1+Nj8cS0vwPJhY
gr6MB0rcyQ8K9pOOpJXZpkfON3JQWURlyKXbuiHxAZfyeywBgJm9W9IlCkeYzlIF
7NozrWaKqO9JHfleSWDO9dAV4ticW75M1RPJIYeQJ+EBVDoS6SGFzh77BNJ6pVYo
PQB0Ye8jzPdRQfnBbQrjGL62H+qzgIpIZ9mSLQ3Re/GBbENR6gQK/zHlC7VQ5UKl
NfyhBqBsB0EG0qeqKrDP+qlAGzgqO3A6BjIOCHenUc3NNkMtxdc0WiLytjcMhiWu
gIdWY1GRM303XatbarP6dGLp92AcnONupZ3qmErroJ0IYWmbxI8fCeoBzZC82gwy
QnQndBQngpWP0UlNuyEgXUH9i4F0fbw5cHHtj3JxqtZgqbS4UmLJ7+Pn7bnSgHiu
L0co4QFsOYuHjHsX7Ec9xyhkhuPb4+CxtauwnYFjAPdDPyQtDTSFAL3TbyYqzL2J
yCkWr4Cht3S5G9fampoRvme2h27P4t0FtqbI9syKOckXrBeiQ1TaYS53UW4WPFGc
BUSNpRNxiApSfijmQ9G3qr6B108tYXN6D160RwGyxfzMqHTkwZ/rI7bK76T32N7G
8EcUsjIOv1QqIpLhHlcgZw02MGuuMx5LK9xhZwxgjqBWjGWOApGgIdAYebu4Etz6
uBlyIGHfAWGiJhy7H7GLgIHr8n1qpdzMxqzAvMXiEh48gPV8z2K8mhqy6+/r/5ur
MVMTLh/RGzJeG6gkTyT3+m21lxfca1LoVhXTF52/kldWTvLKay7chaTY51U9/ITx
yQF/K00MGOGOg9geZeYX5vxpxRSU9DvfprLTru+6l86s0pJFsb/qNn+tswab4Ii3
m6O7suJGQiT+jIGHMHDs1EXpQnpPLZ7UBWW885frUBcN7IshzcqvmgeoCbq4/IhZ
1C+Cj6zvYH+6vkbuaj2HBoOk8HYQrnzf2DV+Gp4le+nNFn93+BIDSG/CQ3J5bbK0
Qm55AOAQs3Q3uW5p+bASxWLMJk/NExW94OO7Vdus3mFnmh8Q6nIdYFiG79qzTTuG
HM5eWSYrPom/KBfkWBDYN6NdNe+SqZTyEVV2l8JWC9PZeOzvkr2vX/GhgGYEy+nh
a7qLMUasotu9DMLxKFWD3mdfygbKq/IiTFNDwI6OeP7us6KeUlraasDU/nn3OAZ6
LrNCRA5jAMzRDl492ekzIfCch2fdA2Z7BELQio863m+Vl445+TdMM1KOOW3Yx4B9
wgZnwALPeyQsOG5ZfChEh/vu6GTBjj4BafYVSLmcod7fPi8ZGJDFmli5yf0QEJsw
/HzLmK+eSUyzP0tNhAohB354hK9PK+Dc75Pq4uP6juH542zFT/sBvxGOo5i5X8Fy
ndyQRFErTLqjesPbUoTzRV8nGpTTIe1KSJrcl6PH5ix2xRB1zPzLyg85CFuNsSlL
s8oe/Uz7YrFJ8QC3tTYsTy7xLZsi4dNohlfB4QnsO61U7H6T+aQNot4Uos00CDFy
301d3zV7VNCQM+JmJljMWLaV99qORnUdIk2L5wppa1aGtpBoVY1AzLLXmWDNPdgB
3j/yRtQyq1Fbc2SvpcieQ9ogjSdEbZ7nQe2/QmfA2pMYiI90oOSdK3ZItoo2nLlw
NptK0ujfa37FpEdQl7kHW0aoS8liibt2BEsRbDTHIzOKpyfbmMXrAvujhvyefmMN
0gijRVvyD0doBX4uxy8zYKXBNLL+N246ZTOzW6JXfqRx8Fok2dSRTRHs7ji+lwKd
cdqCrGDOWEzpuWkJddDKelXB1pwzjHid9xD/9RMhLG9r3HN6L/v1RpB9+VnKPvJM
sUcgu36XmNMSHaRPLX5j+uOU5d1A0TjIRch4630kHSHG9IAp59hfttJoi8yCaq0L
fVTZ+M4wCJ9/GImGbkWdPbs0g7WTlYcp29ca4F+dSLoKHXnlv0nbEXz63oNb+otu
Ped2Lki5ZLzPMijckWPp9w+T+6J3YRIGJgbLkjYq8b+vj67hPFgOdtm9G2smxN0U
Uhwm+ocilNiaWexThPStvEj834G4wPJsqGEvRWHs5/STEaWRerXo0quobVkdEbFr
sM0+EwhRvdMmQ+wtau1VuLtMQF6qYWeQC+ZJvhMoG1bzBDveAvjn55YcpBv/m5eB
JeO3K1fkf8YAvQ3NQ7phkmKYxyIHbUxJZQJIew6ykk/sP2Rd8Q+xzYfcTw0J5LEs
D27TVuUYGQi762k1nFSVZ+5X9BSw5+NETCA1Aqt6ur5Qx4+tHpnct9gsT2ZizfLz
fV3V+KHL7P9+lu65588rSxLg0vz8UWnbyPf09HhCxKw6rZbIFXermLOY8prTYZXC
cu3JvqbkIj0bEazRaX+Gh+lRhOjoM6nvcFtMZ4CS4FGpu7ZSC9zvjKrVC5p3KhOj
1TrmGx+2vwjlUgaZ+CEy/D1PRBLRxKa6NaMJOLGBqcdXSWIZckw7Eud63xAcWB+t
RO6kNw916lp2vxhpMVQOskkgFtpmEbYs6+zscDZQzIW5FmEs7nLJ94DcZ7pdZvHI
1eqYpYNpT4yMJIOs7wUw7vVaExVugS28F9WV2ZI7FWKRZlijBC/usSs02oGZWWOm
/nKC70FGSxMhFxktdzErmabJo3OcFBOJB8mcEqplljMkKap3lvDUSMCW6t/jvSs+
TAd+VynC0AzESMVDno3r6H6QgBjyQtDsCFCGBZp5hCyD6OmDeGGNy87y18Nr8K5u
aCoHejWyWG0CItiMAv8Z2GT8J3s9cgMQuxIBlSU6nY2rOWhV4P5Zy4X1C5AtiVkp
IivQ0Zfp/XI8ZTOD7XC+pnbR2+Tk/cFyFZRmgIxTnBZKI6lmTzVtPIxK4a5mnP7p
0SOCFSFJB56HZvQ36zQWgxzrF6Y3U2eWOjv6YeCWKqeZSe3ICnpiaW6GLAGblCY5
+sn48GhVjutMNLFRG6J3bpm35V3gP0A9Zb0rSckfYl51Q9AH/zq+17RpZn3X3C+y
Zdvc2bmoHISMC8Gxt5anEECdz5yCXlUu5IU7/HJjg6dxlVERvONdHjAEzv6IVBn4
yK9yVeHcWvTsVCT5X6MqMKj3WWq0tWuLG2XvfcaL22igdNUb6szscQ16vEm6/MW6
UufJ7uLI5itmIbSmfxKzLLMVgOLIdowvbfXQuOXrEJYmpmMNkW54ydlE9g3aNZKZ
Bxy0OR3F6D5ginZPUpt4H1eGGCYkl4Tmab19WyelOfgb2hP7LR+Dg59EVqVAYZM5
eZ3gpTaKmFjmjlAgfiExmiI1s0IFYVsyBTEtGW9VUTZT5ag5Yk1nc0nIn81X82KL
PQ0FsHTsvV/jkCHNUfwelSPK4f1WEJ0D81HLD0EjB+x2FunZRUZVRYT+HL54tM0H
OMQ7OS43lEpl1XF/Oks+1o6r9+Pk6Ympg25AlPMJCgWXfxUH7ZmGHUUPvUfgl7Ih
YXfxAZaeg0woEqyNDLeL9IVjjLKtsowlzBnJ7qrpU3GNNZSFho97hGqW6Mm1mqwO
Agi59d6d/UwSaoyzARqnrKca15PnlPEKZziVc4Ni0PRmafIKmTid51lVHT7p0LUD
GK7BDptnPQDqxdyLkNE1NM5cCRCezTwH0N2UssTHke9QrWqh8AI4pXJCwn7vSUeZ
UJMGhVkmkXr9NAybFra1r6zmVE8/i5Z7z9L84GDVBsNKYhvPz8lgLRx4vSHiBphj
RhiVBBc0jftH3CTWMaHY4skLO40eBp6r3N7fyw+KAGuqEvfzsAIQRJizHxR67kCV
wyyJD1hJnQ3YeQEVkVPkPStQ7HQyP6C2apk7YBgoJg4g8/chbEuTFzu3ZqHnK6rH
GWoOOJdBi+AH03jLpwQxB4ZDy3mVo0Iwo8rQO9tZ6/Tv5z70AcjU54AXw5NCZEqM
2x7ES5AIj0ToErkbUsUHDg7jlNrt8+83FzdRdQkVCt4RqnM+SJyOGxns29aFDWIU
9pWTz+3SRg+Ghspl8FZ69UCVVZrF8XKqvlUd484aydhKODbST2NBzR3RCitOZgML
zjhj2Q5yELKcflBcHPZGAvPc0OF2vUD8amTElDVIGTOxtVZ5kAkEuY55iLz+rHTb
LyeCTNjHaZmuF2sRnWzg6+/Ivm8/6oX1x/5rn36F02bEd5jLQvHlCsS081Ula7C9
Ln/D28MC/Rn4VZJtmEUc8cs/nnIR6M1MWMVmyzwod+pIw7gRYUsBvXsUunt+2QCt
Gj/3Qo/BXwBY/k+JLnzzsm2xaqaeeDEBzyTwzqLZ6EM897vnAl6/14R37H5iLIx7
nMy/2Qejb4v0DPj1ZwG0L1vphT+9sjpl/RSKA4ldOTUJvMsA/nwKTKQMgmi/s81t
2hg3ykdmnDD/KqIN8fS9U/88a3lquriPuEPnGW19aiwn43JZ8dL+p5x6WY/LNbtR
IHO7QYUzJ8KQ5n8gVV9KFsm/KHbk5JyZaLaXT/MDc79YssQDwJp4Y70DuKG/4CYP
qZ0sjnnbL0JeoZ3kfwNxwVeCoLLJXePRW2/ZTIkOiuPGJQBa6Izl7tuVyd29RtMV
wuf5e5xgfm78q7oVYxf/xX7WExAejFe546NtaHV2W5SHVC+oTbXQjOu50oDAXsBq
odqZkjKOumQM6uqzNmo/TXoG4lJH5ZaCacj7Xjyx2uzz3u3TB1sp0g9Q3DqVIwdj
4CwP+exff+Kk31XU73frtPJO6BiDawh8WDIpjw6BrnVmEhcjXtnktsCHSDj1JpJx
s+EIDrXMtojkw8uf7PV7KT6GC24Gk/EufBZ/UvHs1jh0Jt+qtb8WshvOIAPEhY+J
XkLDfpUQUTVKJ56ZuMrDu/VN+Ukv79K4fCf8mTlTtym1TleW5NXC+GIT3Oimqp8V
R253yGVo9sv6RzITQjZRMYSKqepdmBbX/g7guJI3/oFURmoVQd3i+delNSoR5DOV
WBuhvG/Xmyj1VSJNLwIlmX4+g9GWivSSUdvsw3s6mHrMdMAsKXIbmtrvB2ljF5N1
VTxeKYTs99RC8l5wC/bW43b4iHl4uwEqoD52nLV0E3Jl5R2fSqut6D/LZ1MdzpjS
3JlGypyG57Vyj+T/OrG/oK3T/VIvV4deX2NAEyhjy1Nfy3u2QKeq/bVX08gUbzOl
fWl9MSRjjG9H9kYOXyYg+mOw7bEppanhlQgCzPsiZByk3QBasRIsxYYwwa+qSFfM
0sb7Dzkibv0H23mmdw9vzkc86RxZ4gGxIuNNFmoDiSZF3vK9Q+LuKFQuoZY50VnC
d8ggoFIHmNM2PQcmS6y3K2IDPZo+sMRkhUhE5wEr3svkaTFIDy0kekD8Lffb8BdA
EQJDZJsefRuutT+m1fb516rCM21UbwYtM62KOfn1MUJqgYLTB21C+s5Mawje33Zl
a7xHcptXw6f4LdRW9Rhyv3W5k/tWdkdL74fj5UiGkLVi2PXGIa4FPgtJ/gsdRxu0
l5VkscXTha8AJl6jC+5T/+13TsfAg/nPalXGWB648gvqYVYZt+NvX/8mINqgaoNL
zVcjlwUQH4uthw27uC7iUPtDY3KEPO6cl5k63zc4Nc5hGzOXMVnrEIdQaYE96a35
y258+TcK2XNKdenvfoBPbMW8NbJo/g+bm49OsrFca5BZadqYivK4JF+rgvquxr1t
lyARpFItH5dFV2kQ79svOideDNbQMxOnNhe49c3uN7Cq3PQsEQKb5fqoppcXFqpJ
eRGjedr5+E+KKF04UMQCPknZGENxeWirs9usRcEdUBYHypad36gJS9dVVg93squo
5lcqGgdRMZJfmj2vOqwEWsBkJh2mbJdVdolVMoI25Q0WogObytBUnQyvBTzJeUEa
xrn182q1bDW4a8WPQo6Ba61AVp6PfgIQgzu257rKaff/OMJM0ZyZrFloA1Tu00Cp
5uAwnJNiAKRr0Prx+vGohUlkYQhqntacYxEzQlntNyMoT8FPU0roCRAx1LVTo0/f
JetqIVOn5kDRgoDdJ091W1MG3KTJA84c9Txf896h2He620nPKUyfPkX+w7XNSMlj
Zc0t/+XxQuWgAdmaIsiASQSKDaeqKdpqxfbxc4/CeEkI5I94+sE49ll/1+tMJvoz
KdyGkWi9kbLTBhdiuUAkmb9HktdWUoy9socepjSksFXWK4po0lQanBUgqNhUpr4s
9maTl97adrrZsctnJAHNA9qZ2JiIiMs+O9TBum4Qj+wDdGKMfZSAkLaSBc564nyQ
67PP3IrrQSiuzrfZueFdc6pZFkCvSfalB81OM0XcrpdgveWC+AvxSpmXN8d846m1
9U3WVIr/KKowJvecrZCF1q+6cuHnF6AB+EvM2wMpDETLqxOGXJ5i/5I8BEqUg0NG
4gzkPdsk0VPhH52o9hw/fz2wqEN8FGTH+j4BrAkOYfTStht9mNb+DRM7bziqH7WI
1OAmhHPNjiVfh1TkhCzYX28FYYODyAUHk1m0KP2DVVoIrLmav9SeoAjx8LRQCWLn
b2KkbVJovbOAeyPQ1PO8ZVaa0472qyLdA++cubudnugTTHJMUwa+dsnOZLkaPG96
1nvmMDUr4ClpTiH/o3XlVCCpT8doZEQZ6Gl4ptugAfTRuid1ycVoHSBZeJXyuxvs
xnI9ylNIyMk6qxmGu1jdElufXUy7EE2nW2AzeewrHa5yfEgJGBtm6BW984lWQUFv
yU+NWQi76wXMVXb6IsLnpGudiA+NIy25sRMUpk/e6ONl2aEp4wKVz3WtNu4I03m2
gjEJrTzEZOtNY+uX4Wu76kCgLPbLCN/ZnJaXKXbAPzxTmVbF2dxW3MMrkwMrq6xU
2S+p/GjgdWgdNln7AjXI3K45Gf7sF5tNI/Zmtgrxs9vYBHzOjvLxHfUWX66j3ZfK
EdldQOK3TJCLprMmfKO34TJ9YmxIqnJBqFdTA7GbCftrqg9kWfaUv5ouEEuvu+iP
GBOhL/I55sYC4O3Iq4YMWTIsFXfkJ0xfuOLMnsnebtV36qKP0t7qpKNRtRWeHiW5
BkCqIWMl6Jafdt7LTLJykWF0ubpL2oM4Cn27KkJyFaA8Jpe4iKi3qLVGcgKiQFaM
S4+DezJ5uCmSCq7p8LiS4i8e/WnR1xS7i8dKRN6B3nCo4zxU1cr5Vnj2/XdYPgVB
qX+qOSg3wv8UcuJ3qJ12eaAqr0ylb50D3nSGD1kWQ7TMnfaU45L/qzHovVw8tnbP
mb8g2fLtD1FySJDhLbqYlIc220KkLPoLbbTAxubIMBZ7MdgYSa/UxTsBpfKLkB10
ZlXnpXSLkW1GZnp6/29eHhMiwJhysSunWlLM4eCbbYT9X94txfHzmFZSPTU7HZNW
77WPEIwq9W45NOvByyYYmyj2ztPIeh719WFqRsSceXLKV8bizjOiBRlVX7DYp1ij
dko/0K3CvoXT/c1ZX6cVSY/Zo/6AD2l0JYC1pg+n/HLVr1hYcuJtEpNnUq+hMnD2
9YSMSPPyROnrNL0Hw+eZNY8HVTi+/QTyrx4o9H3RCxOWdJxsFjea33/bYUtyasRO
cf6wCKZMJd1eN5MUq2bu08bZ+r+o4VsCLHB7hlb9JsknEiWBSk72PuLl78V+EzLn
WIlF8J68Q83tEsgoAc7W9T+qaLF6ySg5LOQBYUOnO0rCbq1SZQPXTXJ1AAXAWjaA
uXGpzpGvKVx2zZlcYCX/Evkdlqz9r/jyRT9dK+sHrM4RQjvdF9QDlrFxUqqXlobw
mCdHYIlu0OyS5YTd+3uhgAM79vjmln9Mqs0Z2emw0TIOJWN8IbSLl/YOausVAcVW
mVOQC0rSdXHsLyY6kM2zBjX0v4aaY+UJYScDT9hY/s9FOTZ05cogVTHgrTxBRtgu
ExDPNYhPA1JaxN8ytoTsW6j38tH+H8W78LFFQrB4xW2q1gWzUWnAv2OQeVQ7zmAW
XVv757C+Q7/we8p8X5djvxNu6H64fEQqsNTNecg0lEqMLEKbHY/w7GemK7F7GS8g
TdbnvJPn9IPlJ5P11z+5IGvif5T3oo37aBWaP9uxTTeUMGlLTQJPvd9o3c2ZZAEl
UW82Ux78uJh3pMglcSfDK9n2n+LbC1yXIJjr+xiOz1elglH1s2hNAaDXk19Tvaqt
uTKMOuPZpSbkoqjpQ2j5smJqDBPhmM0J8oN+aPwx/I2iyLYMs7YgCRubG9OeUxgW
rOyROqNLnuqaJHLvhI6YlZqIN8ZiL+0Q5V7hVJE+bFXfxgxaOXJvw2JQq/MEPDYx
iEYmVaaGtTI6gJG3Qp6QBaXxL+9WRGAygHrRMLxs/breJRKReP4v4J7AYvfRcs/g
VJBRnrCVkJDsZJLppmU1pk3iTA2Q1a7ybwG5kj1xK5twnv0Ciy/iAIJczKg5rKC3
MS71/lQ9EVFFb7Q0yOIcBV4eTPdNiQ2Eg7E8DPVqJxYdT4jDSP6M0nuWYeNJVNRY
D9MUBuv6gYKFMQgv2K4mlSbRTl57StwUxU4kHlMF0Du5JiEVRm3ZLaBwmUHeAdfk
sdTX+xZPMkQ5FAAxEsdGs+oTyrK0g5bsdtaaIhQTQ1G98+CztFNKhkPr3rbJo+gE
eqs/igbWG6mmcW6qqmlXQ6LGNx+AAos/TkGORyWlYT47ZRtYze+YcMGN04TO3cjd
0rDcJfU4STn01L1omLde2C5PGx5JuVoH5gOR6+ZeKF1vk6BYCBtUyXQi/yM+HTaA
DgAtczUYCW7yYYIVk+pgPhQLepEOJ2JloRfSqESvGOjP5eWZuLBcIfy3ebaWreD8
6217hAaJ3EAIZKFj0Pi4J89P+sx1UhI537XIzSpVY8d8e4ssgxqoLHy90YRQb7US
3t4Clf9/aIgeenKNDJHd176ArqFgy7KU/m7Q04qAaSv7H4VhmTKykqiEtn+Gny0G
mwVk+FZnFW9vQHlV/a4UyJ8nAy0XPcoRDUkQfQW6wGGwYUG4MxrRSiTu39BLn21I
SMQ1x5fd8maWgA+X+wkcSATo2AifVeGQ4M4L+DY13nY7zsoQxvegC9dGXJOBH2hp
B6wFXk/kZkWAzByF8/aloWfWwc3dwsRhffAcDHbl/VvzvakX9KxD8qhS/VtIeUq5
uiTbXSwYMjQPky28hvGog5dyPjp2fLm6FJ9rzMOjjyGFYzMWftq1ltY5XC4GkcVo
AIFd64AMOU9+MD6DWLxYI3simOTdgwrobXZIE45inVqFENZPhGtWY6FlynQt4j1v
/XGFK4d3ibu74WzHajl3kEXw4rbODprWwTsf2cQjL2Hp08MJYl2b09kQQFpvNkKn
cQpVv+0QDzlv2S2wQnXD/0ym46JOYXceL/KaiJJBWjczc5aEjKS225g1871d1Y8E
jWNnvsAVM1EYJhCXEfhF/rTGHK2o6ZwZZ0kbnqxFWmFzcZiw06948rCbXDILBBTk
sjVvWtK7LgTFW7RxIk3dJS76oz5mdJqkJpmH72VxkdrF9jjPoPTn3g4lkciE6/NA
TqTyv7of2OZRFpskqi/oECXyt0hlRIcJ3Z2Hd1lQqiLV0J59cEZok3eYOaWqzFzi
nL8Du9CiKLjlwfIKUmvYzz0rhj4OCifd9ArK47XIYHn1MjA+b4mHvLVAaqyZUYj/
3r9xddsMI5Okv3zlTgrB+qAsd/F5MdxYiCEN1hkOeYmpx23+zC62+YY1CfjH4WCM
Ot7xsDPjF52MslgZSNyxUnGgeVpuMEWxUCVpTxMKdlpe8jhb2dzj2/BPRddths/4
XGUm15KkfpJV9j8DjiG0/T6pcYh4Yy3uOmHigKe4yjC5MZCzObMNTkwoWQltb2js
xLt8fq8o3tMQS2O/oLTQD2hiE6jMuSTx8fo42ndieFD19/D2C7qSTFSt3s6EzBFy
AejTASfJJRuZ9TNcIdE6h1DWk5c1PtolNdI9WQmqMEzjjm3cN1It4rAg4Dh73RP+
d45RrRXNqE7E9xVuZYjCGYSDvyawoGRDyuj1v4DX/uWCTvpiXCFlrS+fkHYB360Z
CwX5TSRLlGKtr9nd3Qanspm5B0Q0sXQEB7ddthRI5TB61OagRvwWKq3Fv5s8UbcC
Mu6TGUw8mdWHV6WzNgwo+jbBhrp4ciLrjI5pFpvNcauRtKuEeUCbtyG81L+V29vG
xUVJhakYfJ8uc63f+ohS251RdRE4IEm/YbCJsukdh99G3flNXyaj2nIgTGl/cino
ztTWgr4UPlfNawmIGjkXB2AFMkLh02OUklUUZcw4cEu0+XaHnIdmdzWc4KirMlKB
dmLuJ14hx7Vd6E+1cddT8UOBrMC063sCimqwyOczTDBMdNj+DbNgYs0LFjmrqYDk
9h3sY3spf0XLfXYnaXzYq0vBOTLhqoj+8OXeV5bkL0mdUuroD4VK2sf2iisJ9zoE
0QGql6hVxbsJo/8eqAOddqLVbZnHmPkYN/7EIYft2AFHL6MxDNIiEi1aqyCxmq50
vJDTDhmM0nyw8HHHebUH+rDvX6kPbFRZUR6X+mECwsmDxEjj6k0TxpGqAyjGc3a2
T5L4HXYMod7ebQorCpBLCeh2IKbYL5kq9KW9xvVx07NjTtRksAnHCK7gDcGmcyLB
zuaeWM8iw314syeKs1sRrfx9l9041O0cR1NP4C8h+92JJV35hAPRpr3v2bGnKs/9
WXWSwGPAX/leVIp4WBiQTPqyyBhGIrGkKjErk4vfZF4U46fguxu07huYMhaeXlrm
RiK775anFqJYQRPX0hdU8Pl4EcewsTgeP1NQuW+dj2uPAqGsrFQ4IwD4QIJPy/KB
NNo256UYh3rg2MKXPMibyKZ3r4L7Mwj6kaaZQA3GRhTRmNXQHN1II04cPYCcW1Pd
fz+x2LkOO9fPjJIkoFb3ernJ1hclIFR+FbyKsTSHtN4G2LA2+AV/h8yJRT0rcXpV
z4fcB+fAbJ5dT5ztxr/NCNXpikXZYYllFoHXHibjBSHNqLVuTpzIzdhOPL7CW47k
yGr23TZYsFdT1lY+vQyunP+ykDpD9ZxrD6aV4u/Lres8q3n5Jl8mYK4BIDoxMTzD
UVFKL7gfR2ewuO9yr3TLTYj7t5jMps4P7JQUQrD2v0a2WakWyQGu2X39p3dVNjQ8
hz/UD19pnAaRpHRJjZ86HydEV0yEtv2R7cGEWLxUpINE0bT1OYPwuT1QE1w2yim1
u1o+tWu0jULqiOnuIV/7chdXpSVeJdl8UhowNFR3lAxAyUaqnY7FUw3L3qXxh0ZB
bQzIAp7cIa66R48qJSuypsDC0JbjOmBBaL4y2138FFvwltDthLCXLp/A1ttxdVaO
HHXakC6ObkiLFwm1L5Vuo7ImgJTOp/U8/U8DC9Jfy5NNC+e448dTU2Dx8Ova4ps7
zwlXBp6j9iIhkNBgpY7QeBeD01vEsEdlYVNphMc+0McoLaTo1HOYU82FtuL+n+BI
GbyGZ/7xUn+78gnkRBSCm8rUqkgjrNOQ5OGV4BWuf9pxFocB+74RVqfUpz54Euvj
I46PypqfCCxPM1xBgqqfzRnUW/8Gobnosm0QSDzolUwKUtR6WLSk23Ejv8Wac8Xm
cr3dysViqyRTaqqaBcO0vBqBDrWx1JYzdaSocJDO0CEHf/ZOk16rfIvJd4RJA+vF
q8FvdSIMrXbJPROMaPZaB/Go7izsXfdJ9ozqMEmdkxHto46+30o9adfa8sOA3Bvk
2Dd/XRzwINoRacfhjnk7BMSR5otQaop8Os1527VOmH0bhaorH7YSwKOjSYoalS2/
PwrVXow+wbZCiGmQ/nItN92xQ8cd4DGJP6W0Un/VRhltXZufYemHMhZkLqSCF2fp
uDpQIZd0nB0jWo1q+w7kSR9v20NecSF6yqITXQpsKk3NNUacAwzeuMB4WE2Z7oqV
R/eeQv2n+uhgVxP77Bza1nu86qegM0zruNftXsXojuIN5MseaqfQG9jkZx/doxxK
wJ8znYBDXdhHozILB65P7zg9Q4tUppXNd0dT3LCZN/Rf8JucukhNCrYE/IALeKBC
yphb+xpAhI4SorQ6JDWHyEXnmwj7v1oC+RXB8MicheNuvGOWC5Tfb4GXrm2QOQcT
wHBX6z2vWFUOoYabdeqUhpm8rDZO9Hmw/CzIBOYzDuoTZtuWCQon5ZVbkjL2hMa3
f0Xsh3aLw5+qW3MFs1Hr9/fH5UHGwrXCNCs1CKlfwFZOaoPHGRyg/03wyNLgLsLR
01VYEHmkrBM5udNmsgmrrKJ3N8XohVGJmFF2m8OLlBGxs/HOb6erY2XjGWLg6Ay6
yEsboIQHoLZpJ6DGJISZ7qKPyLr6QEcMOX6DxzqePnJQbmb97BCb/3dT0YJgZR3y
/ZGH6CKG2bZ4RYek4jr75o74zaC9Kwxs/80/z72jLp64zKepskCSsfzUWABVWgJi
GeVQRasUqtEg5rM8rCpaw3rQW1UnynqEYFcG2vF2ESNBZ01Ikq4w1FQH/g/tT6Nc
m1LZ90tYHKzgtUwaXLNf8gG17eJnM6UYPWuBysCPyo+nWbDo65NOQOBZhSPAhawj
gg9GLQxXjKbdwLmZQdsgBcek7zuh3hUW8a7n42UFgcKCfAGJJ92g1YsIMiKkNg+r
j9uBmf9IE+DW7n2Pj4AIbE106Ewe6+Yg+ULcChpJQF4Uwu/fwBW4iyHmqp+5di/H
m5xokpxU2vTAYaiLkvwMwi98qX8VIyYYEkuGzqXSP5BzGqw2LrtDownHQWwxp3Wo
cyMWYNLZHQ9t+xpjbr/nOP08u0eLXSXh/KkxK/agEzIDXYxOPQhgp2d8KvNvC9aL
xmzwnM7D1KBnvHcRUOfTCMI6/6IBsIdTlfWUcF/B8wXu1odRzxXtKBIPwvC7JukL
POO0wvuUG8Ji5diQCr9IyBJOIeYIOdsM7XKyz+98Ht9IWIDgDxutiE689Usz2dwA
SeELoVPMg97vF4wYWGO1kbsgFjZrEqv6GVdlofCrZTQfZ+BnXjFbVsJErhNQIZsd
+p243ZXMgxc1cGIUdQu7hqMNiBr1Mqx8vy2r7KbOLFhhqbe1R1GTQTMLqC/xTY5Z
VNMUc1Z4xU6JdqHi1xgQCQM5Tzimf19okFD/qCeYZAdnJa5sMh6GvYhGP0pxqR9+
A0VLUgatmmkOyi8VsDcFgIuvYjAUbc3TTEq2qnLRabCpQ0z7qXc7reJ2t7htWfD8
hmWHCNw85apZEiT37V48/gmHmFbF1+Gyz2tDLKBpE5SjTPENMfbImQlgr7y/+wMs
oEZJChKEt1qO1mqHxF4TUdrWqYdXIJjuqG+apHcbGUhR8ivgrDpsJu1DhstDIRvc
Ba+SkjFW2eWIgAmUtSKkHiGTEpsFCHC0U8j5fy6D5N6PXGEEy7APCB+i0ykuVjQZ
V9bWVRPQwkQXiMqJWsidNCGSs4cNB/Yyd+KRLl7ioXyk5WLlD7cCkVgdJXZit8WZ
9POMBaEm4CIKkJwJZ3OWY3CVJxGJqUF46kUEK2l34f3KXEuJi44cwX2MAWqJog2X
1kNEkdMe4XReHHkgYECDUQ4W4XG4rW8SSCeq9S60DdWCPmo/I6EcVnpL7vl9y6ve
qrtwPhSSRRltKqnuHF1AbCViq8bf83dbY/BYvCY3FeFqbVK+SsP0tn8XHwnO4dyX
6F1KWEnzXyUucrF6s9OeND4hvgUB7785/uj3JhzJl8kVlh3qvio77IhBvtg+Av/Q
QMwNR28LGOBxm2N0+c/+4wf6V202X/N01durnOk5Aw8YrXPeL/J8Y1DBHIsGazRh
4HQEE71/rLz1TiYTc54vVzbwgkenranpfIL5Z+/ka28eUQ8SSmSJI5ELYX7SfC5A
PIFBN/jX3lPUSPl3i5jvI/KVoZMQJKlRNOW3NZ/e9eJCtUh7CtDjATd7i2057J2L
Iabaqq/wVv/oLYj3rUUyNAFSS5aG0obLdBkGnJ0HTSym3MCZq99+pfI/4a1DU9F+
T0RPgaMcNIekma+dQG0Cf/44lSDx5UY14SXoVr8waAshIgyox1TxGDfejoOdYvy5
au/NF8QQTO4S7TFVkpGaMlotQH53tlsL124V/ZVtSS0qwjmR9GBOwAC+W7NWclUP
hJlKyItSjSydDhJHQK80ZplwpaqorunGSaGiQap7SNGckzrpdgKhOltnO2FB+D5j
P1u6KxNsn8s671MvBCYfLLQ6PHz4GkuPlDHUiAv7putAwD/Q4G/LhH0BgTDpCaL7
UHy8CU7M84UD0Mk0B7Nnuv/MLZBpv59I0Ozps3FIZI5D/roCQNjULKQyKQ0B2LDj
ToL1yEclYZtS/fnZzXCyr6ERyoxkawUS0XyckIwUCeiSDcNTHwyoYWAjBN9SaJbt
5HjfnXC31l0a5OgdNdbQqOkxEoTxNgXRPjFghVGT0KrpVS0LS+aByHWLWn0k81xb
3VP7993Sdvfa3VxFw6LQ3KTvVyMykghOsyZrgHPhnRRVqzC6Gpf92ejFMGeBHp5E
twnSKCMqi98nsmIyZ6OR4oZ1lTBLG8j7qToMkDZSDNZKS/yy5qLHPZ6XAxM3dep4
hG7p/gCqmolM4+7GzYbNHysd5AcRcAvE+luTjNIYwk8XhCQ70f+nS3OSgNyDP38S
ko8jJKC+qGEPsk9cE/TARnvCcCSMhwPcjkvAIWBY91pUjl/P24AiRYFusIw+oq8Y
pgJrLP+M7VEUK52lcpS4grToqd1GwVCu3EUeAYitv6oRRZ/yeKXslx/E/CSE3hkE
oGu3U9f0pid8ac3LEASjVyfyd8aLv4jRFVPwC+cnBIE0T7bZ8rPKC19/H+CsRr46
qu9JX176T2Alo4ZHjXG8kRaUbpDzOpv6ZuQq4xnagi/pSa0X8KU6y1TilNGNwed9
54XuJw2vDsmbyWrwZFRc/UtvlnJ0QseVNUqSlM1LXaH7Ur7Y5JIzLU+SC8RtDgkS
ohlsH3f1dlvNsiGOSovW2OSP/SUO39WfIjKKlwP44ixNyNAU/knyIhu8MIAS/Cx5
6ek48gEwJjhmhPaxjZoLlGtwUKQ4C4QlPcOfrlVZ5f7cHeO0UN39VfBBk8h4N1Eu
Qorb4d+84FvgDd86+c+gZ/sFUx5WKlPeHIG0zxw8PIbesP3t6BpDLxo2wrcV1lvB
amwQBAN2wPAiey/Kbd0W2y1E3oPpoAAJ7JkTrWqYUx664f7XMqBGeZKe0wAqmrvh
9NQI7a+q3GG1HPM5J24i8MdEdsRBzCcbVlkaFWoHdriSGByUv7DaDu3pnZmKDt+3
+KqindWs3/l4tXrzJ/Ly3tjENzv/ZgROqAZYj4POb0VZ6ElOkbZIuu2ukqOmEp+Y
BanZ8UbNH22TYOtrSRyATAe8atMDodqKRkGq+50AR9yfcqnspzepXYhf7LIWUf8F
y/Wd1oqVhQM3H1q2jvj93RU0A3ThJNJMxtS4CMhXOFuWm1zS5imcfNZsVRQK1qAX
rpHOEAH2bEXYuevWFEfag4Pz74utZwBI2oCCw2k1eUIjU1Gs/Xugp0jLG0Q6b71g
dQs/8Wg1zprm3KHBg5q6XvjVkFed4EDzdxCVpPbExkCw8+iwJ1zLjs+VVJApHBau
6WAnr+33dJ2Fh/9ZgMsDQn7IRLmfs+V47abXV5trvLD3w/C8RuyU7xQUGURUwoAq
5cin8tLOXkyEuG0lKbbU1OWDRhmcJcFMQNtVd5BNU64x1j0IoKFUTHfoXumO9Avh
K2LHFGbKvogw7UqbRCEHUTCjDOK+33+1ArTZNrZ3A4MhLYk3gibaA1u7RRuf1sn2
XhFwVqW5iXEdO5yu85Y3AxVwe8k4nMMl8lkXI7diayKWUg3u3D3IztLLQro+PUu6
79NrCL/7+sU3V9JyLjwmf7YANQ2tdu9Yf9MfSxIHtMZxTY+SXSAPXD+nkpqIzbbD
06oz/ZvQYj56p2+uRc0NfgHd8cdh6l6fqVVhTRANSqG80qYRPc8KQabddSYa1Md/
EcaiI+2K7ZjYjQZllQjYihjnogk0Sw53rGFqMXFjJ4TDpSfVcmQfGHxDX81ehpNY
bDcprT/10N5R6016GOW0Muml8vc4XLHZWGpkqBJawHKmX9fk/QfWLNUDYEBjFLp0
Smt3TmmEP2n3f/su3NjeWDGt5jvkS4XOpHuByfyypJd34vwKqIfeeeZUSIxZAQMA
tjmP1j/LTvuNdaYHydZgwHnZ0CTw3Xo8o6l7BVS42jqoQ/kCDTI180l3Jn4w5yrG
Dyy9Lh9he+oFRSeObvqn9XZlFJVfV8FRBlz++0gkeWFycdF6MMAP5G6QQRhF1CGV
MZtGYeELQIS2EWiBpAgN9XZwQCgn2COvs9+gkY+O4XyAtzg/eLompIKJjccBTwhN
AA0p0RLboUEhzbt7SZISroOnLT9hnibz2druPqDJa/KQCVAHvLH+sFnfcBdD82GB
EoXa/9mObvq2fN5PGkkK7mNdyqI5vT9eeK8BG8WSrEt6U2qDhXNpIm8veX7S/ibz
chLjIvDvAKOS4rhXhtpyMt1HLMs7icdIsR155gGPvudSKsyXZ2dpOpUw7rBgFc7u
C4r/jsFA6v8BkPxF+1Uj7fiXz1MvshRnN9bRcHS2/INuDL5XyoWgdYd81rDOisAF
vhCgxErUaioFXVyKqhSFnYmj4Ao8hOE5q5A0DittNdlInjCVfFaQqs4QoD+SeZ2X
QCsbsHm6B39EjV48b1t4WMSVt1VkAYQftm/tAUn+MjLRk1s0XLbQIHG2XSvXGU1f
+iX60m4hV9+ALOLmar8jngTd1wCXZ5XbEByU4AvTwxRkpBWnM6B0Dxj+bPOZPzdQ
qnjYSAXVg8FPVEXdHfPK7kpI/nwTPdjfcQ/MX+7LzTMkgh0oQ6wwYl8L3aaZB/RZ
/Sgz9wMdJDQJUVBlil1fgpSLjJZYXMkQmis9Mr+lfuOka0aiyaG3/mrY9BkOjAYh
/RFAFnaK5u77Jxgc7+MxwWtLBQvicuNadH97H6aAO08H8GVnjH+vHUvORQRVLIgr
wWwKn30B8WblWqm7k8MoBSvpiNm9AUvTZt1FbDD6mk8gEwmTIbM3ObNmrRIqvNdP
/Op7UeHxkCOQi+S/UpibjEzY4bLkkhLplnZ2cdPKyAd7n/hHiCnQ7QHX+dym8qfW
pVgovInTUdDSFTjWG1vBdRTUTl8Xwjmr55o+iY9ukPS+KE7DY2s3YQk150U4xl1R
M1adJjBW2F23Omy0lBiScPms2lczahWc3E7o2bUFi7YdXz88rOk5wzjT1GLHQ7I9
Kr0SHYmjJGLyuSJ3L1sNWggUeY/cuUZbFXUcbcpayzAPH/AF4typ1IIuPrF08h8i
YwwEtztYyfV3S+zbUrhQmCihK3Y4JoBN06dPbiAxmRJ+6CJSThq/zRRsStdaiCEo
8VFyVEARK+tBUNmobYdlvJ8TKV2zZeFHZjG2gKd+50LIJppHnQcYKPZ8JUKihoTi
K7eSOXl6I6Yv3+HeSfCpLOdmQJb8PlcIKpfQJ/mScujSvMjozavxIpnlAHvusZFJ
VqK1eSFyBNBR+ShGKmNFInXMq/R6+081an/ia53IexG9OuDRTgnCnkJBTN6TUFiW
Vjg79EpU2ieJ+X2tJbLpoBrQqvrENed41g2MyZM/bqFN+UEM145QKLzA8vTuakp3
kHZ4YvbZBvjRDOHdxjGsgwcohvTGzpSuEyDGegDlksq8XLtqUuZpWO5bFdHQtwL7
5vC9Xp79KYDgDTVAqP1RB4J8fEHDlqqIB2tiT72JoyXb6Sg0pV8CvVakepBdCYzS
P964nDbaGMe3/F5KTxTqYh1xU/yRJuwUjfJm4kJ6wlGTURpanhFNDTpiIG9GPomT
9lTBzwnOEhCPmKKFWlrCd5TIjjXIgq92wZfkQ1SExv5ozPK/uCVg7X5bc46Mf0TB
xhNfY/8lrj5I3MSUigsfO/wK1FVCfB74Kfu4byp0QE4Lp2gtIaLJjlDh3yArIbQK
MClQSEFn+tZspt9TZLXOEMEv21nhLOPu0TsL2Zii+CZ2v1Q1NK21rMosXyo5AQ4/
fAcAvQA8/Qokj9V03FUBfVNPjOXj0jJFwxx5NkeT55BjeoJGOHMi5OmxbZt1YgI+
FuUGVw7OwuWEc252d3FM0/1YKaj7grgoH5jg4E0y3cNBFl8JHgmCNGDNnSWeCE+0
E11pHWGlhDB72x5FqBzMakr/zxpUt/WR9R/WCcC2egrW5kg+JJdR58Y2MgMGWlzf
1wThP0FDkBTfMO71KI3HxP/4+orCw6uRHPce6sDmEYQl+/6jxgoeGlfkO/I/Y24Y
JS2qAS34HG+LiSQd4kLUGLxTp2j2mbmu1J9KIa+AufCLOlSMqRn1BU4Pvu4skleI
VcqNZsgpq8eMDbubEbZY1+H9QwIr5RwxrIo43eTZSEJR+rbNejvQ9iUY7FcBrQkQ
yLWyVlU3KdPduhQ5fVRsyplWCoMpUAVwJVG3fktmSzCSnZFXB1HY9NQZSiNlQGVg
NckVcp4KHF9HjI9/OAh78QCFV59HDSSY+s2b/kxoIelQbTswBUzcRUwMnA6Nw3/a
6Ha//f1gY50YDx+RVNM2g6JqsZITHlHh8sO990oJgz+emR1QQw3v3/UOQ+K80l0g
TcdE3+6QsaWbadwRdNu/gRhnfktvu3jzcTOQgGEKNrUI3k7Wy7+BkF12YalmJv2P
AtSgOVz2+YHJBl3xxJMQCMtpyaZvzJ6it943CBFS4/7iD7BwOhq23lAJ/D6TSyAQ
WSD94lU96LNlzWQ0rqcHe14dicgZ5krBkeZks8ka/Y6XNHk0oayx5OHVhoY+hDrj
sb41hjOuMH5TliJ+hAt//G72NkTrs1u/xk+N1iNA25X/Zf491ibXKZ7HUzyaEzVX
KrFw1O3m3zVsUYRXlioxizW/74jHIS/mRmYg422GF6BhFSk3837VhSdJpsFEI12V
FUqv7Oxtchp7u6PsyWyDGmf7r9KUF2x+ezNP0cxSMLTabD45PX58pQnNz5yNeeIe
1QU+E3Li8LNTfccRA3368MmjK7luszsn2YyhN77pzVrDr1zZrwyfNYW2TcoDyrjp
b8UB8upk1oHAaIlF/qIetV4LMmDuqdG9kyuZovPo+Niw+PbP5vTtXABLxTqUbA5p
dJEfj6dt946V8DxCPGOBM89TxyMGsNux+qvYno/tw5v+Bo4Z+d09XwdicH0cEAv4
Swjh3eViXFubvH37yrzFEOq/Epm9L4KuEiT4L8MI+uCKTv+nGva+/09orvuJRne+
LUV8OlCiN0A2QQnmCuR7Hwp7eFFhqH/EIqrrTVkXVzyVYgcjZ+KnioUB5F8PaTdK
c44OQpjNoLmFDgYsRgzBBzHwrRLkPxXqY8sVo4Pj3mwGWfJz2DPrlLHc1j+mAHVF
kGLs5zrVFyDOAsPJvrbl/oczR2pK3UtaeGKlmXD5mVsk0tEp7HjK0Re1tVHqGczf
HsQieW292r0Fyi/COyLicqdMbKYKXm16XQs93EgvwCiqmwWl0MaVfnr+8ospGEPv
h8uWbFfIogBjHbWUUmAhKHYDm9XLMl8XovgYh92CqLik6eiC6n3GZY/milGFANDX
AW5YsiKzRIdkV/vcorbMjcDsaNwsuyImPVYZtCzadJEoh5HbJBc9trIZHdwTpDKc
V7kp1lspegmvmN8CgTmW7DJeBR41GJVvzUl/HL48hT3IPhsvGmTooMVeHZzFk2AM
ZYPFweGa0SbIcd32tDH26Ripdw61AJlrTorMrAtStFCF3Ur5y2qEKwPif9k3uoQP
x0Za/PMhJAaHeGhYEX/zeU/wamQ4QE4BAR73LTfjU1LCCbp0r8+1wAOnr7YAxP4s
RUX1Y6ahyocTv1HeeCZDD2Nzs/U5Ou47NLuKho3MFmdQ1hVghmutpx1e9cQIdeA3
qqv2S1FWgljNA2cHJws+zoq3CBg2X3Mch1mO30SeapCsVnWzxqJCvdzS9bfF1lyl
O0tkgyV2T2WjhKiKWbcX2YQWcnSRWzyJ+Q9JRGbTo2Lhh1Z03R2vq6mPsIgRRIxu
87FLVPXWBmlWaQdFQE9zbmHLVbxKGR/w7l2RtTENdciGJH3VeKUuPt0QfjLcYFxh
X2EacEspi8C5FnmxWZiG+1P+DUi/gdzDGwp9lPe99o9yEAhJrkZpCPJ/j5gTaIry
qX3+amhqCYro+WOnoj/LNumLmKK53MYKf0dr//HBmi70DwL8mNY+HLZbcemv0C53
CO7B8Xp6frDhnc5goiGMx4vdrj8Xg2WM5ipsYONZ+vt29Vrz2seqwM7ZbuS+4zpi
YQK5ZaCLm59mf2c8kkHDMPaIl9OSQcU7WS6P4ID7KZGd7jjBLC6yGyNQJadGI3bz
gTvx2+ddxqFRON4iXMWyPfKoNTnJPYS9wbXpEOBkjtwsmUneH/Dzd2VEsn+Ump6K
A3qGWeJxB+qpIazG/cwDgzd+ycdEBu6KP4UFh3SdIgow5b/n8r5FdtZe5p90LwL1
TxdPQN9UUsJ8xIffDwnFGul4a/rZN4hfrTUMvb417yAArXhpYnGy8/cTFeARyLVH
WWjtlbVwPYAeD5OR9ma+XEjm19PsEvdMCvz7e6Qqufk78272jwtxdMZp/uGaYOtq
QETT4QoCPwOyLuEb1qWMiIABA3aifqqVk01/wOWYhnqBx8p6CUU16BwOOk1xwspz
SbEuTiSREel+3zXXvDwD43vfZtruJXO2GPrHG2kZ6y+BBrkmn3Zh4Q6g+l8WuPH9
sqxGpc1qCJ+Sjc72o/nlZbWl6oDQWaureOPAyuu7WvGf6qEWhE+3AkhNbPU965f8
hs2lZ56Xf7QC+/ADxf79n3SH50yv/Pv7c34TcMetZHECne4OZ4iQU6l8i7NjNpS+
NQE4VSthBUOm6p51dzQJBp7YBHT1uRPo+tuT9jqjPAY4bKMhoqx2gZyeJ4S7PC67
i0eFVt8rgNF3R5i0NBRGjq71SPuprVAB5xkxoqyj68iPoZg+rZQ3BDPm1i23Ne7I
/tNAmIP2KSCp+dl8KFJrfW8ZOUrp3jwNNzcS5UWfyNlutvbUqGiVZnPIkSlj4iIL
Ki9A4D6pBvUGJE6rPRkDpNgHVTGhxpkxtgSH3gQd0XCaoo+awII2CmP/VCbeo32W
GHEpYgB2iiwS9bcMqu2dol/lXyMNVPUcAen5DZCPJZVTnW8nyhTTQg2rqj2sRpns
26X5IieSk/L6xFe86PEPdD6Ty9F5KVMsMUybwrvQC0uxnV9JPBucvfTDDqYVyXH2
B9KoaWK/ptAK7zTIdW6uTFFlVvbXhMZBuW9ehyCivX6Fod1KZBdLQkbjtP239lqP
Cx+K8jw51M3IViWYofj4JrvfM466KC4ioQU+KIRitYPSPk0C/Ne41atU/8n0D2uv
LX5UYk6dfmVdXXs8XSNx5Nkeb6DYkhdEB1JLaECLYKorStADAg0Rx2yLIz8XW9gU
7xwNi9XxSY7Tk3C4vTuSCB2MUpYyunrMImgIbZKU84p268rvSdLzbEEG9bkBAmJA
jbcFKPVkCDY/PKWkAAAMQSX2UAvYaqPWR1N7CH5eqc1V2V+ObV5kCBbzs+vSKoSy
y32zRSv+DeQL4wM4gFAQtUWB7a1cxNOdQDKfnkSPGT2RIl+jIp4TJAUmWEBIVEc6
OGE5TQF+NEnQW/ifHCFVGyCET2+zphYvIL7awrgR2gbITTGvuhyLrK5WNu5shfEh
bXDCXKlSondWlgd7JZm/btiUHqTUv9G9KZlj6DwrM9hxueeTVbMtgt7El/xR3s/y
hAlAla+rObJNoa4Y4Ldc4PP2LptoWAmNVcjUu4gpfy42nv/Y1ngCoqKKxhlEDLXG
RqbbsUfjvIZXJNoKNqmggnhgsuvoyFJ07k58ApYVPjebIhcDP82kBzFMSR+fAIgt
1OycHkqQMvszXwo6Vz5PRd5Iy5Mli6AHI/asW9N3FS9RCBSGrPWtu29kmn5fXb+o
BVTVzqZEDev/RsRhNOCxdz0eBdZYTNWaDDP6MCorSMyJbZ5DNWxc/R6LlB+KUpQg
DcDg5vUfi8Esh99b90J2/XS81opxfJlfMuGS0NdyCC9/aS+hCx51c/EHGRD+qLTl
h7pIcDqIIV5uyExilTifihhCKzU7hHfNMYMKJ+VobZj3UXXtoZjx94ggQYGsM061
CMmqOlgtYxYPyIYGo411mlCBVrGOxl4PZBO4k8tGqusTlo2j4ZETITTHieDOKlr9
VEg+O5tfulsVDsi8dz751YsIf+TTK52sdTyCBd8DWa3W+/5GjOecOqnvaZgFiz//
fygw8iirMYyJOoCNLSxpZnBzRaM1jRSYJbns0Ti9yVcHgCH+CXU3/FSxJ/WTsdUQ
KWg0qDJI0USPC5Oh6DA/HjKyVeEUQ2X/kYqqWN90uzEtQwD/8nrR8+UeoFE2QbjZ
16/WNUOpWTgj38P+lr6kHDcShpC/4KSgxVzQoqL4wHdvX4jVguVYjNSC5sP3RK+Q
tDkz65D7dImYvDEKhr+ylSImBzKbslYl2seB8W5xhZqCgu4ueR65uW7mL/AwGcGd
GD+xYdKBaw7JYaa1MDOOc87xHlgbyE0kccc+Ga08qA9/YcyrB+3XodaU3ICFtqj6
2oNnRkkNQaLeFDRdRUEX0u6oLd5Fjlb/1o0SA4gpiwmyfN/Lbsy+4P7j1d/GzT4x
gHz+Zq3VaW6xJPI9fhENYhaxl/DVs5wI8nDczsEA5/wqzTm2o1O/OfzhixZJYEKO
a7zBs0uo61G/6yvPaWqwnsM0F5bCq4OwWjS8ZQlk4ma7erag5h5wlWhtif5lRP26
Xnrd6emm8sON8JgVjtAvMar7/8TJ/sdiRP+ty0jNAhaIJ3ZI1/XFiAUW7QXb0frm
x7CEfrh0NJpzv12udfx5xrI/pCbzNOThtOHn85aJktfaxLmLSZAONEg7atZAYwbV
GAqDa3KQ+U3DZ9FSjza5Bt1dsKj6T2qfCTP5nJZiNIpIZdPrmOBrs1O3RnX2mDiZ
MdB/hHeMobmkF3GEz/fq5rIjdeqBLZpM0Jw225l3DdgxDvXOTAvMOVk/vJn3e74x
9jJyCSBoI/CpBGP7c84/DoqJtEAyf4gRksle4Va7UnHed3vedu2ivxHFCh3WBhM/
ziNNR0amyxfP+vibaEafCxndrgF2pdLFCeO3HdtH4bOeCWII58g2DPNKw144xjYg
cIewAFCnLH8rSXRbCKzetKvJzUrKddaTH9zcLkl1Y8CgcFIJGOBwb/2CPmHo7cfS
zkICOdbCIXOmL+vQ0i6NHZ1M4f6Qf6Lgt7bHYLATZCQq3gzFDn//ab2i5/XoyRMq
ok6ZWXchTkvZKBRzN6frnzoDvswPYqlrpl3tt680YHGnquPdAPAPDZv+UQeS3qsG
d+GMwW3+pSa7kc3QpLw4QXCieuPfp6Q6Q9vLC9TczzBXjVcdmDPwfpXs91ReO6DX
E4GWFgacJb06oT1rYt3kJMfRcLSfD8Hg/Ip76eKPeAiUjRvKWFY0MP2fCX2qCGhd
ku8PIfPdqEsZ4S9pYUUUvYnUWcr00U3Aok8dq93DYnb3WtlCBEc10lZLTtBAf8S8
rnjrsjFCoW0fTfK5V5fJWXF/yHBKQdatGXeOFd+s0tiJsJ4wO+o1LbG5qlvd3hDz
73CIVvXaI2eh327lwPkuW8oMDgdzIAswle31fivlOix0JiudTKKQHxPNkEhagohT
Zue0+HFmfCfnjKDXT74h1nWVo7oI/uOeWskGNTC9a7IxuwUWCl0S11isp52C1db0
2x8qp0Qwoej9f80wPIgfnmMLXjFBjM5hU+OUoYHLvPtCAkkGCupgDWHdYDzv3hU1
CMNvt88J2LdZ2a1m8UxAifBgY1vNvJCGPvFSykLf7sx3vsWYKR4A7yxkbY+CDG5b
ZAVdRUNNerWf64tjndmV+lsgQvAetI1iGfrbMil/7W2DpFcqzib1p+8u1BPrtB5Q
q5xhIOZhltpkk21nY7PyJ7zRiqsG0pv2+rW+xs0huypUiMK7tW27x8bwuVhr9a0Z
KxbV/Pw5xV42e1rHPDxhZ8vjaAAax/ynonGGGKrEuqK2EZqv6LwzFwe4ZWUUieGY
UbLevklwafM8h/TwBtD9zIfLeZC/3A9mKAR6/Yfi+Qm9edyhqecghVt7qvjEUYAO
ckUj6cYo8oBeRJxm1amJuY+ktMBTLgizRrn0LSRkZtT6Ugs91R0Ahzd39jdOAkYX
Zo5vJeDTrkE6PtfxeGSR0KezyMu+yH2mEzmCHgJUtIlgx2Ebe+gJ0p2VQ5zSobiQ
95f6Nk//aZLc5xQlCrIFGIpT+jYSDbjndnk46RaqnAE21nSqqYEMNe842LudNwIy
lS3vEzF49nFJqqIwLTi+aLeTGPvOR/0GgFvQozI5I7dxYwWTasplFJKoC7tC6U7T
BxTt5Aw38mPkzRmeqNpDycAXneOzsIDUvWZpGmX1levIcEvtYmVVuPa1/ANxhTXJ
toAiSsw38oMnYxLMr5j7p9tX9A9YShccAsPmzPcZEWLVUuON+6NG6XpudGkFTeP2
gtCtE9GfF0cNmB4cUT/wz+ndQPGEZXBHUOkUvlI2zLmblMQyH0ks6UnnhSGxim08
kfekJ9gsfg8AgQLhAd6J0pw/e9fB9KFBK0d0cs77JBAbiSjt3OkjMRBHF4hSFja9
se4EEfPLUgaFn4N8I1pDhTgPUrvXJfOJv8ROFI32eCoa5TY3ZkkfMP7KfsgzUfN5
HraCefhNEN+HW+quPmZTYWrPuyfvQYNR5vjVWJRAiGfELSnHJxAo9UnZFgzKq+wY
KpurECQnUbq/+yZleK0yyP/8o2siwzHuHDsp5qD3WJ9SP/GfpGj4q3Br8Oc43PIW
2MoT7ek/YyaP34hHEfQKJApON/6HZVFi5zOYIoRv3eSt/6fMIromRZzJ6eVY6Z7f
sw/BDp1vwZp7WjrAdT7aXSp+6b9aLXEkQKw1gk+3Sn9/MbzQ0HD8OR/xgVDWQbtL
UQqAjgc5pr8gpvPA5QkXcfg8+SyETf3OVlLAFWt1xKII2LTDrf05BYulnwSzlflO
wY3Ehj/Ylf0fSQrf8Dm/0kZfLGI3e4e7bEqu2+sGVhkOhQTbcqq2wr5myCPd0bFa
62BX7mMbpCNUJGOUGqeKeqYQ87Wops0nonVSqxw/IvFPe5GyDW28UHn8aogA31Re
7p6wti9fh6alfOHbX/IfNdMFGx57mPACFcNemUM2h/A6onhJi2EaQGSYGObYl64h
MpILed/CFw91NZNHD2zOCYlcktqJaRGijStdMtoz6nXDjVdxOdVI8KmqXOQvh8KB
ZpP/ygh06tqdBpc/mJTDOxT5jtR5ZtAHgUV0QZ/lcD0PdRI8oWfNi6kutTrnsPMY
8SyoR3od0vOuvYuf3Dwfq/ZyLX7vECCETPzDGerBAG2qjq4u1KFNEBsPNn0LNrtv
wjShNHonr01zUFCYjuZcMBS770E230hVBLYN3cy7hlLmFo/kKPB/5osgVexDFYQK
1QHF9d9TQ1htZRUfQ85ABNfdQlfA55VQuHcUh/uzXvDupH2YUR2JvzN0LYsjEIft
Og2dWkMaC9tCBMHoIzBe2Kg0hU+8LmjgKiyFCcZPNFZX65qWxtxRdeFmlRdNUTg3
44ICHCKRpMnbYspreHghorQmyyaIh91qNdi14JMHVKTUJuj+uhn1xdoxmbtTppXy
Shf0Q+aH60qDN8svG0oNK+yAEuvNMev4JKr72YtkSaqu6PmW7RrGBaO1FJShYx0v
Dp6JV7pqaiSd8HLHsBEbEkWvX89WlOiVez8psMpFNfiTyK3BLgyM60y74tl1Dmaj
WXtTPcIYreD13Ys4z/Hi8X7x2PMzismIEIJO/PzQk57V1Pix/7jKJkssw1PYri8N
qrWCcNkwYdsAGSk/NxvwqkPT++tHf0zgojrh9xgM+jdAvDjzgZKuPK4UNIEt5NQq
37M+2vuuRJCWvyTJC4MlJ4IUc91s75qGkdBoQu2VCtQO4oP2c9ZdXnkFylrEn3OJ
QHIEUFcnUZjUWFAHfk6OTF0UCBr8fuJf2tKkRY364w4YOpoTj1PK9l5Y3gup1SJD
8Oe2aD0QiV4hZ6+jjVqs6XJreoEY+SxO7+WofuQY7WLnJ9o2t0PsYg8WQ/C+PZuf
xEWKh/z/aHxxiHBvtDzEMbggMUyzAw7ThhtDFhDV//5LehS+4yba724tbDFZ+tTW
wnMYMf9MMLW8kJ+ByMkE9NQ+FV9qHA+1guKExWvo5+FiWfO+pk6EDHmtfWshNgXt
RMTxTabXXokL5T8yb1A+DyZ9ErhMVTjaYneTLDQM9SFOIqtH56n15DqEMuxEE8cr
ydufHkBcI0pVwNxOP+HVvslheuFzFWji9Qop2iT849HggwPaZ3rFVGley01PW3Dv
gIab+Ft+VM9YBSId8ak+0RAL/oW3Csx2ACkgUi8aS189ei1fV82MXjruZ4Ftal0E
WYPJNVWY/BFIjY/oyacQA3vZa/PsQm2AnYju5X3ADtGdBlUXpy2NEbdEl9mbJ3Y8
Q+jmmlPUvwCzdi2Hnq9W8pdkG8J6C0zkkQKHf5oQjnByUo/peaaG6Q5R+hukGGw1
ZYCClbvaqL0WcNaqeA74+Y1lr/mXgxtirmUw5WJbd1+IPjMsb/MmtuMiWvhgZwPP
uxkSVhykETP04neFQVJdFYSHE6HftstkAC5fKccaHc3/vrftJe/95Sge7/nweBYV
Y3d0cd9zhAHKEsPp2e0qb9K0qzPc8svHwPSjxNUjHMz3ux6L96NTe45N33ycCmMy
PKdPaq2umZtZmaSFFK2MPcydUGm53Sfwd7aTF0RkESi38DaNy1D7ppQcT0/0y0nk
bx+VFWZWj18WsU0pVxOs8IhtXLkWYTI6x+aSp6dhmqlhhMNOglrdI2+8nyTG5qsa
wN2rIr90/hY0CWSQjIu9jp2fkkyrOUAO5rJs6sQQIxgcTo10vbHbNClT7PQiG+gV
eK9n67tvwpdPWq8Jz1aVSEENSRKS4YedY2fRwZhQA1f+ESOF6swZ9jcsPNOIfni2
Ivrh/acEzTzt3N/8akAw5RqZdWbXhxQnlIxWQPrhuqMOFWWQZNPW2LWIUNxklEX9
wmeza5Iy+5sFwgS+2how6VOLJ/RsC3Ih+vKbIp2RkS6PrF+PSWPN8AndK1l+26FN
xTDaKaZFzECC9CapAJPPXOT9DvbPs79aQGKBWZPNRyiHjgs5uQ3HHrKF69BScDMG
VKrOsTONvqBU8+4IsO6dxMsJ9DAVuU39y/3YP/yEgCyss5hCvcRWv4QiVGN5URne
0qZrM6yvaQjCI2u6/EeQdLAmpp7nuRXKQ2T/xMIeEpiWKSHDRtmnv5yNmcL4qpU6
Nreon04DVnjowqvuvtkkhQjQLmT7NVPiU4XK1UTTwJTQ5HjGNcIXlGMVy+62xFZu
tCshdAEUdgBsnIzF5gO0KWPjfEmbK5QdsIY34dUJlabEXfBRkp3J4eyGdh9A4Q1T
1BfI8/5iBLvjXJ2vZodPTrztbMFX6ZgUOkiqb9JC9DcmnEZTdTb5Cvgzmpz14AM3
rAgpjP0pQQdIOaxbdIMwALTrSLi79thT9DahFNApZBGa1uPO4vJo8xPOeiaghZ8R
Eg9+JreiRkPQ/wxFbSGsY2WVWp0i42sdAG+egf4eEz6JcMgOSi9/nMQWoifX+H3x
P8mhQUfFm0EktYCgueYvl+SNDz7BfzlcUw4Qru0YQujPKquy/3YCFDaiRBIoBLzj
yQJ8ud1hFpfsvdceP5itLbvha5CYOO1J0XP8Z1hHyJD68giXAL70Wz5U2VDuWV/o
yT63RnDzmmbLoyz/abmaPIYLDxq7mgDRerNhOK1Sxb0lL5nmzwhpXB52EloblaS+
xqiWtjYTFYP8D3K8DUaoNyexHpT2pMVqERjD82BnSuoUGsweAq4P1pUq15uvKIkv
3JR1gJE/olY3JOfUiKWEW9ulb/sYTo4D13ZzZZKjAi+KOO0Bmt+RQqLNyBRnu4Cp
wJ64FKgWpqT96au72vxuJkAAyx2W8NhhPUpwHUjXIQUOQS+zEgaNr2E86mNbbJJE
NbQT0hYYRsoalBLBL667pqbMQkfxWSC9EF071zZmo1votvZpImGvljir0mYZXMfc
BAnXN+4pCD6eNz5VSBPUHrAdN0f77XsX18/bycJOKf0Gij0cgIFH8B6OJmjw6h9s
mHwwNuT9obxwrlQILYkDV6aBJOj9r8xi0y9+n6qYwApdKBHXZ2N4OLP8oFQpk7np
ppLbnwev+tbJdC+Tt0A0cB8Vo/waDJCUKIve8+VKuzqQIdt5iy2RX3EtGTu/fxEe
k3AyUzr+gK4jH+y0BTEAwhDq18333G1sDYTwKcshQIvhGIXjFovHhkRArCh/KbUT
TlxudbCDbatLU4nYKdBWfdHSRhyLFGg+o+BXDN/Co+SJUPG2outLDMLElLFplyke
aYunNozqTgrvflx15aby6yMuXWwMG8MdFAe0q+LlH9tpTirdJcTRUv7cV/M4q3XN
jTI7jt96sDsaPmyrkoo6FRdTNx5o2oDQsq3wMQKUMxBK7vofSkuTFVrUA/9nAL/c
YElbXEtHoDt7JHuNz0eSXTuSpqh2FA3kBSXyDi9Y4NYP33qWHOPoRwE/oy9Gi/KL
YNJ3+AdqoNAnAc8yb50DjRBjka/pZjUi018vi+a3W0ni+QAJ4jGSFYjtKgbvPRlr
hC+GF4pOk2shIbiPmae63wBIcMWmNMN/6f5vCk6jDPBMo+eVBGXIAvJ7lV0Mkhqc
s1aYifQJHworiPJZcieMJ1rZkJCs7T4vCCbJTyz2eaq2HkbpLRhkSzCTMhh3ih6V
fyixhnA/zRSCzUdJcTyFP6im7voOy2H1bmlZUexK175pHrUjRdCXBgYvluEk0G80
gJ0JuRt1vlaHC/NL4X27RntHeuAPgZZHwlEYPdoGWoXVbBsZh3uyI4FtP86NVh+4
fmI5jkFcWx6XYMiEgjspv9ngpLfUwze4cYb+S7CdUEVpVS8mP77BPlvukis1lUdm
PoHdt0vZKRo/qBrZ8vW3P6vlR6NuY3ogFRzLDQ1l63GJ53MejGPOMk7S97o0p5GA
PJ48GlxcmWtP1+ceWy+7oiwqP6sZT89pTTytAV73g1XF+DHCaTx5lAWDXce49SDd
26wcw1sGCccDjnes6BxzeXmne9C9HEfp8qguut8koJCBjN4Sa4bvE4Cp/NEOvV1o
LjwBeNGKhLdHXxX8sp18vz4SKsgLEOOFk6zfCLunk3s7jIzzp5vyaZUyhBZ1c5xf
oQbmGwbRkcwqBdx/3kwPtvoebbWfsdE8rhzhx/Vaw9zayeGL/7uPHIah7kJqODQy
S/+19usUgs+BxXtGwYYrOSZnedkmU7+euQcZqgdRGDSHt79TfC5+HvWu/sglonsn
0uZbn5vd8zt1c9/0XBNmdhxxgY09I1BCtQm2tosJPnCD2LJzhVAr6L2g1p8cz/i6
Fjokme6x9FopEhhZmhoFqnj/SCNcNVOJ2zlCfaPzfucDpavAWrBVbEi5wrt+cT/1
OptsacKNELy7OdgvjI2cty53qZMUa51ePf51EfzmbBCLhf2UzKYpiwsBikmaAVms
opy/t++7t9CkjFBjf9aFDOJxMnlaZKKIISaD6MyT1qYN30/M7vZoo0O/fBN6zGy5
Bie1keKMV1rF1Jeo2q55JOHcY3Hn0uKvpZNlEgLec02vrzH/DP5HhTTRWFntpZbw
RVLq7gUiIJ034N9NwmfLKIyryF0JMZIgqeiHB1TpfHMpr48LewTe0TDdmDzUEFRX
jslvjXLfC7WSUTXK44qCMPzgdfjHqpGZyWrlTGuyanuF5NvhJPjvJHWZ8c75wcFU
MgqkIRR4nGjeVvdc4LvKW8eYfImG4QXkYuVxKcSW1Ri92qTxmwcuseDLi14r0f6Y
4B02n9SJ9QMHx604R98bIz6e56zrrDrscu6+wXGJOAv6k3cERz0MkeNNQddzI13T
U6N1jSqxJc/qyOLMB1S+SuD7bPRXwvdZmyPNTaoI2/8jfO+TyhB0JnvvEHFY/3eI
AQC+yOjbUC3d1VbuNmDOovBt+TZ2+xZttu6yyrSGB+3wvybTday6TL5Z+cE32T3C
WPA+lMJ9EbCMO33VfG4oMac5eEffDJAfGZco345kKdfZO+I+JOZRCaxLeWVDJjYx
MbvzNUzArfgBxrLq9fgbEPJg8WXxubzLQMOPQQ4OPAKR0jVvY0+EPXt70nk2rWqS
yKJO4ySeXjOdXyyWAG3gantdba5rzYZgN8zm/LJYP8aCykr19nOIQoGxrGJWxEt7
7zvbP6dlst750kCw2Q8/usFnZnQLoLNiZJ33YnOlca3/TliNbcumJsHz5UhFhYfG
9RWBv993yJu+83o3XGJpRQwLn4lYy1BGR/7ELUEI44C0XmLPsg8p1pbpZ8l2isiT
4jeZ5B0hfr4pFD7VOLLN2P8iF8xyizvct6WdWc3XWdoxzOc8jhOE9it0bNGXvekL
Sppk62+h37XRiblgwbjuQPvtBgkBS7LRZ4h/hQtQS5sIJTbzgQVOjPdAHErCC7NO
4K+H4u8Cbr1c1qZkLyjGkcJ8HGzmFo1jArXg5NPgf2zppj5hHWqXsBI3Wj8+Ph46
b981AZrDHD3e07Cc+bVoWLP2YIp8/h+XaUg3qTCfURAW/iR6GQCq1SiFh2Hh9JJI
1pHqLw8cY1Rg8sguYiXf/GV9LVHt7h/LjHbaSSaPcA6nlprvsmw95XS447CO9xPN
rPedLkpjrcarNRUE4bEpxdPiFSF+2Z1Sly/qN0r+oCNZA0tABvz9zwWVHuMb4xSH
NsxoUQP1A9mRR+i2bpIouq2JsSX1zK9b0jFbeTBJUeviqrexHtovvg+QIAkM6zcY
JlvYXP4NDQo40efyBffZyd/l84+JqyyBSFS6F+8YYkyWEKjF+cvDM73DVgbT3Uys
03CQZxvrcwmo1Ni83PjnW2FyS2gOkeynqzHn1vL8I+xDUnuPeQrd69XD+Yejtjd2
F5I3rt7gamSpPmlmqkmWxvoM1VQbF8NKHmyPTCd3RoasAORH8/kXP6SFQsZpMm/1
YQHacVLwzCzyEJdhXYZuc68cqCq0bF3OF6vvL3k+D/tEYRPUX2YFNn9TNFAH8gYX
RwiNs4oUqLbWx9QfdT5E9Sj7akPoYMKenqIpY78FWjCKFqdT5/gFjIiCI5WjfjpV
IbsxQID+9997Rr26Jt9OQL+DVhqVA5iJnnZI0UnwoTle9lQWAkjLZCUSVaG6IKw/
MLtIcrHSgKEe/GzsJAZb+/zOgR27/BgzyvYFbL9bpdIqMBlpLu08XPajA40MTPdN
bbNMJlGMYHkA4Wi7PWwOeVezQvt3rwuXmsahQYbMGRQCvlkUC1QJxGToMushEREG
7Mgyf2wBR3VfjotZCQBZsu9C9uJg8VY1nftu5krklN7s1v1bB4RGg43Jgo/ZhUKD
6Dsq6bjKolryVxQ+VRlER1/v9nC+wFEU4Twsnitt2t2JnyzH1tMHI2pLw3m3v9yj
cwekgnT4gHaIU5yG887CPaYROd/bRwAnYZ4amxwdhdHFG1BDU8E3n/+wtJ4tNRCc
bJU97Bm6amHADbyB7LvMPsDP75UzWTnhgi4+1M6MMHku/4Ncs284/mxUxU/c678j
WNienAzyoBXV6qjg1uMwCEDwu2hROj3vCrUI/nzRzNPKZhCa7AhAx7Uk6L7NRJDo
VY8Gt3Jj/qq1i/IMHo6AWTMoOvLCCdjoXR0PduRKxpzqczz2CBQK5phUaArcCzpn
CP4dQW/Iae1qI93AFUMFArR9px5LQAeJkrGofvXZ7V/vskpWX9SRb+ccoDQatdlK
0aURuJBh1YLWp/j+LwENBrQleE4MP25NkQu3FGvHatfiF86GU3SaIz0V4/UlMv5+
UD4qI6fJ3vjTB4icd4NRisCRpO+oBt03VDdI0YBTY7pAs2OPgt+3w/Wprb+SwPkz
x1OTxoWzg90qBavzMjWMiASoUevzWnvsr4IUM1LWE5J7XFPcsqYoD1iJu3nP7vNy
q2yz0lrVlWCr8AZVhbL3NMjCaJlekpwIHxhGS0YWt24mrnLJl0pq2FeSEetblKN4
xzmZszZ3TZBZjYMUlTG0NmEODbvRllLVYJJ+y2rhy27kwHn7egJz2co+b/cGNNHJ
UWbKUI5fv+tr5K9tEmJ3y+96Hd/jAs/rZawNLICtgTvSBEBQmBFYI97QvscdyAcx
U6cO7z6DM6TiNvak8ivp/KVEKV45WY2s6wIW5cYXlu1zToOWMewEftu/WX4KzJ8f
bykQPVBoNh1skuaas/JWVbDWAiwAHLp73yJmCK2Xv6VF1TLa45gzvZx3X+8X9bRM
iWUbENltQKJcP8MyBbHup3jqlSBLtBtIqgLxfHhxPai8C7rGfbPpL5WhmAIRiIdZ
zk6q+57ayDinXPAZH9H1GR/9tUdlfs7J84yzpriMZ3uv9E8Dv1rdoY7eEK1K/wnH
4r1tyZUOq5eRan13cS5aSMIpxNy3JPoNTNaeDcj3w66vIYoz0P7KQtOhpbu43a2R
bQYi/B1j0uP3MNYEWCBryAt27/AY12yPyh5p/UtgJFoLHmHo5C6fdA1ADaXb4bvj
+HbZe6jRlyXjrif2getnLPhpBMuAcWsXBIc1W4ZpunzMSfBN0Oy5xwNSf3csso8p
7JUghcYaHkkYUHkwNdqa5AKqiQai6XkfejHZ9Enr2QKCEBs0mIqQ4h+CyQf8LvtU
OEKX3tnI/2bE60IcFDPR4HJoGyPP6YZR8Qx8j8i1oab8zbeG7IKDePUavjDUVgO/
w3a34rruwTxhzXCtqhiQbePZfYzYcPfcovDswlQoHhH8srDV/NvLbVlSP71rETWz
U8wzeExL+PJHoJzXynmIGrCynxTf63aUZjbsOchAWkZ5KHFm188bRRd/sViOf49w
GdNsgqJUseikRu/MlIK2UPVUR0g7E0MUFkhW+2NzfmGJG/+4bPgA7iJoI2u+XPIW
XukanhSxTJtFMv1Q4XhnDIa+j1PULD2cLi2ftI4D13LsnUwEKtZxgRsNvYL4lsaa
x5jbQl9sOLcB7qALp39u8e2gfxjLUq1N7nYcswBB8mNbDx/TYddYu2C9005zrLnt
Sb47Q4AlWOSXNMF0ro3Kt30aVpkeMuHp31Y/FL4BDbG5Mh3z7yhWzJS/t2x+sg6B
7TNq5A9zss9uzvLhKaKyt4nsRhpG6K/tjPHcrKho3I+Xlg/0hUWf6KYFNcnJd8Ww
SH9VXJaXW+F867tZiat0DeQD5LwvZHTuSN0Ycx9Ice6wyKAJJGrHFpsY3FJ9LAqF
R1BNpBCO/+jCCx/QEPOJT+slU7GuNQvIZw9cz+ruNvax4ibXcpoNarfDK1+2+S0m
fjvl5q7bvsHhuttYVmqAT+GiOhe8w2vXQbKZtWc0fshjEgF0cecL0EcaUUSAVfBs
/XcnNU5ko6W5Rcloqj76rHPj7gnjo0vIfEqa87hoH9UCw1PZnqGeqlckqFdlbf3W
tO6UO6bwRYgaU71S/RIaHW6FxFoOt3LIV/nAmgrDZZxG/ebTeoSfliQle6eYtKRz
XlQB71bF7TpFTfrbFt1g2VydAa3oWxvLkS52gvEZGSLmcMDWLRNAMft3LqKge7Py
r3S7I3NFNzIbqyAHA29MhG5tUcXGzv+4+idXqiGHBLVdwOOaJpAf0n6/Bgbp4Jjr
q85Qswuh0V5DOh0JiohsaaPLL0esLnXDKK0cjPdEWA6Yh7MZviEIOuViK40NYCeq
hVF9x/v/jU92OyUKkogzdt+nKxrDtRgRcrzq2TWAeb8p2JJolVgPZCqhhSlFgqY5
e4YK8bDkF2CNc6yIXsAGVB3OmZ2YiPdI/ldIzA6G38kpnMmUEyOVn+F7PXRmzi7A
f2QwSWD4m+SuKvvFv9k/Jc9f333eTwge0YLd/3eWdY1MQrmCxUWdV28HntDKdlgk
BFBFnCsej/89elraQBovGrdRxYkbeNpM3WqF929JopzCoSIVcyJ5LBgFg/8up/7Z
UEVJDn/quMaB0udPkXRSCK2c1uFoVo+tdEZX8eGK+N8RjKe1N6NJWX/OIiAKfli/
ik1sSVgYKFTIN/1rdiiqvZdwUuvdaj/fzh8ucpy9UhrIcQmVL+vVM2mdgLhcvNqk
TE3bhbXWPIY/8G/nuNG2vRUO+H8NUWXKbnnjzf/8sNLHEJL4I6tpvvoTQYBmejt5
hjyQeag7ay81Hry8Xgb7cvZBDXisXc13PIGkM3v/Ev8fE7pMr69j1iuuDsjbGWXF
Oper2X0OgAz/J8ktYU1dS5gpju6TWDvuQXRLp0A81fTBDqYcYYnMieYMSEnBcclu
QjKK7HrWcKdBlRhfxCWTbTfq8n9gVbRQXXPAawBQemx3Ccl3fnhk7+DQYK1K+TC9
mmmdPIP/gF/d8iZM5qYzMdOwa78G4+ti4TDKhuNDoyt0GfR09+KRm2P6TEywozNF
HC4r40AvNl8yMuw/Vh6K7n5NtxPNGNhyUlFRaYprbkgM5rd6MyTXVNedMyPhA8bi
FEU9/KuVZeKT7tKr9g45gtoS+4FSfdHhXNJiEg7jkzlidv7amxvMofv3InHl8ErU
po5sj87u5WIMHSHlJfqGgLN7Qub5UcuOvI3tBVV8wfuqgOOSxS3e9xoYlNrLPtUL
5Vy7trrM3XfPBq6vc+Wf4ie32hvb84W0jxRAinEyriD6tCeFxIiB19yk8XZ5haWB
P0IucGe6wSSKaQHYyNy2Ahs0hdUArvQMpEmWim7PVDUIUsfFfTZXtNTBPWLnWX6W
1QpmyVL2v9P4i1PzNOJlllPHQU2z7rzIqBLrbTqivEUx6CcjGHSW3sS+ryziXLme
xIbHAtvSOSGyJv+HKIiVjyldvWhZuz+6pP4p0gqN7bZyoBiZ5m8zjXZKcJVmmz0U
tvjYmiak28CUgvmJyOOl4AaAap9AY23OY39wX5ACqvfbNbFdJaRNyu3K1vSjucI4
PKOpcM+s7KaS9zvF7eixV/EjoUf5cWVuN/flqcbEevirtkpBnnFoaeUrNzSnGo07
ZiI+yFbP0cLyXh/HIc3YZqEzYZs3INwBKvGF4od4/7QFaa7BETaJ9yt/skrlJLdK
rgyQJNqRpAJqYmn4xKOUWSlzu/ArXNVlCclK52horbZ8PRAqVnobhtcqMKuMF0rs
d6yzXQtWzknOSiRv9VZl29/o3lHar0Ui89qpB0fKBYsePSvHSA2zIpMcc1pTF5Lb
BEI8vT1BX2aCU8dm4JoDbTZH4J721AyiXWRNeZFoHnBpJGbNJR8rwEd7MSnMo1QG
m6eVysLaZRuyh2Ph3FZsLWzL2I5ODHM2NrqUGvSKzz1ZyIm92+RQvLP2HmovaH1s
H8h5SSB8HetSMyy8Xce43qO0KjEEqruUXJImJeoMNOx3A8x+w/efgY7d/s/4aCJy
HEQsV9Tvb0KY+/KjXNAwFgkfuNVyeAahU+YhYjqrYtTadBM/AaibFpzenpoRanHh
P9Exm18CtZKG9qhPv2aJPIPczviY9KDFv34EwDVLZdcxmeXwCqNdIgaReKNWu/1G
jWbi2UY1LXk6XARcyE77fmnJcB1b8iUBl5x8JbX3X3fMQg/UQ5MRhHa6BwLOPgOA
lVwruuA/hU3dNXuVR55ZurMd83Vi9IYPlz1sshndXQ9Ty9H0kpuMEm7rstLVupka
X6HEcXf77FTzln+dnm3Jj4WcB+R3NIJj0gb9UBKQgdhU+wtPfsMKkYuzXUrorBH3
8docxfHQ8scdW4w6Pckwx9s3aST8xgNNQXfP2PpsNqYbRvX5CbsRrV8th83IqK6Z
5JkQHeBvHFKnF3l7zqC/Zcv+wWnkuiQ1MNBY5zR3meEMDE4YarRjjVCPHt/OVbg0
wEi/KXTpuso/l+YF3FVV3ft3YjRdqmJ/1u+SlOWVl3rFH9pbw5O3NY5BUdwhvoPi
bL7uAXyhdKAHSjmJ9fFGYkN0Yy/4br+JG7V4Nn8lASw2WnpI9uhFlFMxaJKxm/S6
qHweL3aNPqG8WlUran39u2VU9xHg/L2m3p+6mfJE35cz4U5MGUs8xwJpBHx82jhy
91FUHl8vf7QX1fsBBe0Un7ixsp0uyvkqt0ZBclXIcmcNdaqAL/Wnd4ZHGNvZBV9B
a89MyiP0YBrFoynX7Z25BqA9MKv73HdzPJNTcAedihV+/4ditJb8odsA88u6zMTn
cwOZoiHwqiS/KRK40AFL7Fr4QJM11VvbfhrtBsNPt85cQsovv9vWQ0qp6w6QbHU2
z/LgV9MIcHJI/SKWR6vdPf0X3SgH8oWlvwwWngitiXsHttXCcg50tLaUAIZb3C3O
4HZHBeg+6jpliDeP1Pm67q8l3quY6Un77H44DIQCgVQSAIrcJe/6/c3Se7hRTR9a
6qzdWI1c/P90Zb84lWr8WbVxESpdhMT5eWsyDGatm31dKbHc2jG2/qtnW91VoNL6
U2x1DeEUYBj/3c3cdGnGvg7OvhDoWMCXO6gOlwSBngvsa3UdC/Anu/wZWwxgZwzW
pdW1nfzZ7BxNu02RqDnpatFfku0ThFttyBXzfzA0xOP8sB1LDhllnB9EXXuLrm2u
Qaka+HXmgPTsLi3MWP86Q/OTTPJzLOadtMyV8ExkMJ9ShneELfL0IUFkQoFmzS/j
wwXm31xvTJbKpwdSqUWXOAgbihznea4l3vXVHa80kj0sjdQqmJi9m1F6vfvL0yiW
lyNvfjQ9P9TjCReFgbbz7cjP7JOuy8EJhKJ4fFP8kVguGP7I4kHeMtH606dqtGom
ryVySU/BEJvGWmLO7unClIGcynEN+IIIygd9xSQa79/exNeMXFfaYerVDI04Wg7z
DMH21D7/VdhUVliBfoQs0EhzXKGXCtB5QC9MFKtea9IJY3HnDmZsUwbVC7w7IV0Z
+kZB9LBCDbhxq0NTPkeJhlszsiDy7Et9IaAU8hO9+8/jfaYhDACUrSSMPgS2sMW0
nS2ZEl2bNApbYl04+y2qfDO9YrgQeLpdaJuX101TzdLqVBW6m7bR9GnHp8S2Q9R7
Eft6aDeLd4dyc8/iiVM4KUOtEKpW25PxAG6qMTz7rSBTg9ZIE+jmw0hKWdYC+c9F
tkDTI5jYMURcJPvXgYzVpojsM6bN4Wmvua5PHcA+qVOTxHor5NC2aOvtVFr64y/W
1crOs2qGvTjRyL/4ZEDqqYh8bVwc4If6dSm8gHwsZ5ntv8uzj/AQKfo4xxXm+7sI
LENl8abrSR2SLH2yPW34BGODdh6mrR5jm1S2OjTZPh9k5wFQ/QJikM0GwN1d5qXi
tW9NNdEvE13WLzK+FweHkyvKYLnNDRZYDEctCjXq1pIKn9JJ7L38+78P0NH1RZAL
C55no51YmSojXZhH/9IljUl6Wuw52CLMBgAMA5VOWGaUe6J8X8zKYKwAR9DnTCgQ
A+XYsxifEfuLiqt4qRjwmmlNo1qH2EAVarr5zvd5i7+yiDG0m6n8xFEolQFt9b0Q
XE4hrrXMtNEV5vlB5YhDP/y9Wmm2cPnAGpdrJ0KIl+hGdJkUPKeIbkjxJo1Zwa0F
tGuRWDyK5xxMC4CRvMwYDw1f0EgqWJHvfzCAXixY065+Xtk765q2uNQUEbWxgw2R
90NzYE1rRzShOeC0HHQsRq60JRfKS75atzeNmhWMpXBOeHC8dfxc8Uorv5FEfpx4
5FSzSeEP8jyqWHDk0VT53WyMpvXIrDcf1LVJyczg+1FxUoISjNXcZYCXc4K/c0eX
EoLOuLNrmaF5X4ctqn9uQlMgtlCwZtGdyFN6AORZo9Ao6iYAa9quv1qzYth0AYQP
EZHnVFRvVEiuLIWjxS/0OWVzEwwC1woV7ZHrMMXr3zgPBteaMujETB9R1+cmazir
VSmRhAiq1EjxLdMCeM2CgkWnjIyEEKqAkEW5QO2H8uGVFPtIIWu7puvufjg/YPIG
YTsbFVu/Ro0zrhxxF5klyu3GMtQP+VT8GA3ydzRVIr+Rr6TfJ7hqnrdwde45VNsJ
XkE2pSP0zwHA6WCFEcNoQyv8D+v2ATvOfCc8M4KgMgBDX1PX2WK+GqoTc1CShvay
BhmU/ZbPnu7+FcOlH63mwcWcmyDRftSXKJr3q8atuy8pV7966fufJZoqYc0EzcHs
CLgBRxmSDZ0vRBSaG9lTcAF3++2Vg9wo6M0Q6ybfY1ZRw9dGeQgG7EMFW072At8r
U7oQKbk6M/wOGHuqSaYTZdnaB1R3Qy8VJmkcnpbR0G3qD50xnXG+gIjpwgSu4cHh
hz9764yp/3ZsmGKrqE2eu0YHRttSdTjXUCduf3Ku3kXsz5qyVL9MP8A70U71N7A9
76P2Y3NwTuvUUB7Z9mgNWptXk82LaEdrYvJshBJrRPtncTU2v+ODTW/lXUVlR9Kz
d+s/2R4ttqBNSV8BXI3+Ty+TfZIkkKsgjy189QMiVS65TMKxfvLmjxNvwTLjiSv2
QM6EGJVt9VkqB/mfeP1i5H+Y0yr1/4gE+/M9GV1cXv2PGGGPXIvi1pSm6A6xPRPg
1CoAhwx6W0EBDxUyqw8OreyJunHKeFvk3y7/FZjAcgEQt1xNy/3p5paJ5AfZIG7B
+Qf76RjWw5aTFk6TcRs+WsCC5oVTJ10KiFGgfLFE3SzP2w3FEruR5dcrVs6wvY+r
7k1RzOOAQPc3qCe9n7D5U9jxy4bW1Uwz3OGqP3+135qfYuaFVPqiktFLNbmNamWG
7fOMXmZTf69fM2Fl++5f33HNBRfs0l0hq9CTYmqYNIQ9imovk2T4EnzJFaczaNak
Pzo4ro07Vz1tZokaQRqy9Dkd2u5w/KR8qDUQenmRamWj0HeysqJUrSBDw6pL3w36
T3gdJypYWS0BZEKAQMdO7ermNq8Zzr9jgkNCwmIEJ7wc31/eVnHCqxAVylnpgJiG
mO40iSakOcJFWZ6tFqmRBJ3kl253s2xmwGQBb3CJKoehllaCRl7KlzDX+e7kgZTv
AxJhIa0HeYogDeOG5zDEX70nkKR45lHOg4tGXGcY96xk1sVOxvXlMuE3riv2Wnd8
eRHn7f7PltK9GF9GfpEbQYTnF4VYUfiRscr1ZFgNQc60nv3ZP3W43fkMGyNOSbgT
U/k/TwYSfu89WV/bpxsUaNyDFp5MVL7Mh0687lrMpB/gzQ7Q3NR+9pYCMsSr/zen
Q0bLkAeB3WrTB3VMwKkfXMlEfVDQHgRM8LtnZvH1DK1cp4LMo5Ell2D1R+4jyoVr
hHpP0S/4d0SwYkYrwR8hYvlGFKZFo8TMS0l77FTU86c7F09yyYg9zE1k/TPFstFR
9FBlwWYmlZPkFsvvZOPUv0FSIxxpbIRNXuJ4fruquZDS9SgPtTJ1EtrGu6+9kH+r
HnS8E7ruVmnq41QdK2VxBcc7uaK06W/3E00AHCrWXdRuynaMW9VcOSUZYDkHQ0OX
+Q1QsZZ3PzBkd05gVIEHRrEplE8UW9NkHBmYqZ/Ni+8+ESplXIJQ85XnbjPWhKbm
f7VKg7EQP4RG033ylly0T4TXOWccxPcBQjqI3TkAProsuuieSGZfJkeH5AXwcC4b
CTyoA6AXEdeKKpsbVCKMBZrn9scgOc7kFtzQOyPR9ibyfpoG/g7MjVODsO23QON0
YaT7fe2gSQyXQ2fk8NYr4QXG8TLymzBvPsQf/h2gVCVcoTvk4Ra+cMBwQMuM7xcF
lo8/AFxXHzjbNQWMXv624a9mD7XHX9U66j7XyZrAy/y6e4QqqNKjcN/P/iMm9zZV
Ft7kNlfyCYYNHczZ0prlpIuFGGqX3WukUBzTrzJYyNvJ1xpboIfuvPHjA40HtxOn
Cvw9N9RSUuuYWJr5xt8sJoGkcnwA3GL1+V6ZT+frFpEESReB/cqi8hiYlgbASb8s
OsqZAvsgCqD9h4GqkEdbRQP5IixaKKgv89fT5oAoYVXTDlGXvyyZPeCdMiNuRdVM
rIja2AlL1EVXE+/8dNwkJLeZlYDjY9GVZPTuuGndPvMutf7EmUZwWpuUzjnwHgIl
orIWFPIotQB6ku1qNSpt5EbMFeScmNONuMN05JLU6C+qjEq38SoovTedk5zV35st
8B6xPnuZgpG48NZW/E1dUwDsi/baG7Fq4m9JqFS78tUw4IltJbJYVfAtjS+SF1OB
AvpOAOy5d0GKvu/f6YKjNgKyetY5vWWoOhlPjiAdI/HLUSPMxCxS4pcmBpfQX2Uo
jkSuQVQg1Xrz3sNLFkDuoxCNKWmkXA89QbY1Ffo14+O4Ov2By8NurzAHHcS+W8qX
Bd/tGGMIsIjy3SlyNbV5VSJoZ/6pSIMFZIFlKLdDiCmAqx4/8lSVYrQjWnNCn4dB
dYI7RAbfd6fKXqDkJ3bDa5rvuk5Mwbh2fukWIo3UeCNboqXYCmVzyOBgik0N8ybk
F5rl3Ui6Wz9ca+HtjEaRhCWka0fvKbjJA6IQaVybLYLBHcjl5QBBCzMGUuZeEma6
bp6i6smoITl19vMru8hRaM7R/1Ci6NUmfxHKJbJF82cWkpFfbI0XLPISWk7A04tK
z+zy4ZqTq2Syp7E6sgrJFwSjnGSjnoe69sAoU2dWjPHCOhe7yCjVeWAcyha49Un1
8jbW7vgaoCKocEPE/UhrvOs7hscL47qUIewfmz8tHA7dmwhv/DRjwBCNU5QGmG54
Qxoq8YhEhWcULS10GBijieO+G+kAmO79qxbd9pLPs3ERdu87l3dhqrUCW9zJH617
MhAZdD1CAh60Q7XMTAC7OdcBBIfPL1Z5giiB3Pdjw2m9r7p4be8t3QxbvDjaqOr2
ifZGi6Zwki0v+nCCpLZlABnKmHnPndDhNIxym0on/3rpxTvm/xPwfMueoNzjbqOT
/8MjoJUwlDQnx3XMIFCPuKF/+RWJbXoBMx7zAqXgLSB7DXzM0DGD0KMYyZ/fJKV/
QtOQ4Fl/GtRK9RaQ6Dh8YMv8sWHoHvySdcWrksePUVuqMNFoqTWH+YptHs5u+M03
If+zVekEoaGNaG6KiDVXki0oq/hj6y6JYerdc+opIOkMLIrIKmoHWABYGEXkZZzJ
EKlHgGLVTtNfPk7kZjZ0VkEx2xrd2JE0AVrqufgPWfpj37MEV/T/6Siq0bMPnxKa
ZbJuCMg6M1xbQeoJJs4CMG438SUKzk+rd9407h4QXI9LasSaC04mvyl1dFvva/Lf
mj6GRYz1Q0ALBTLFa9/I/rUXK6qU/hcJtRZsL2RhMAA6JU+IAsijrEh/m0ISKLQA
yP+r9wTCqBsW8wdAs99OmzPSyWaGdRERr+A6sFSGXz8QCzlhjh2Izrk+/raAusLw
VEESft/90rDe2zo/tvwVnQxsNN4YzEu61p8cTwlISQvs7IugrzWhV4ZVBbOxag9z
1zhDk7IwUQEk0z+3wRWXcdviOoY70GYguoLQI7CoDWnAdwocxjWfGU4nDSruXtzA
QPRNaD9f9EWW0ahHSCcGm3c6lQnPZ5bqRZuMRgvK6y2NR1omuLXg38ziUmbnFUlD
VbktYDxelkLeHrfvAj1JLOH+AJqU40K70s1hj6ObRzxJkXEz6jn7kTAt04Fg3eFv
YmDkhoqfKF7xjyzalujP2Vg9F3mGK3E64DyBgrY9h9TpFym14QSr4s2yx510c1bD
ulFCeRd8S27SyQ7M/Qti57mRRl6Vf5cyNuumGak7JGMjiEyuQV6mDPR+nXvX9E6E
zZsmtk2AnnpU0UVWjfsZAPNE7Vq6kqyRcELkYjSvw4Bdd1EzmeQHc6gq4KgRL0s+
A1H6oeaAuKiFSGSU1EiRYec3xwZLE4l8iXlROK9QN5kOLnEczQjfEZ2SuLqiHxY2
V7yRKgBO11I9IR4qm9NehVKMgxxF/EA7rXGTNmLMJF2DzPe0nD4AkOcDHxDZpjTh
ibLdUBPMGMKoD+MI02ohc2uJGpvGaWiFmbF6GTLjMupoWpLieEwNLuWve32zTD5m
dGtY78tLulbxOS6RRu/UF/pFjufwG24r9KjZzL9wA4I0vApIhafZRhk/oMpI0kXG
KYksKxnyO0BVL84F5joXCWQ4aQfIKg/9JKtbIWnIXdGXyhYwGeknSamj50l0Pe96
0zT+bSAFy8HowxIvbtfhZdJFuzwVn8FRtKcMLc8meTNLL3Qm3+cH4NTjeXZWHA31
MXOfAs+cXT2ma2kNE4dQtYvMnIqSExZvNK8r9baDlDv0z9Y1MWnL5E86Bf4OYGdy
E5LUF2lLUAE9i5kQYeFouvIitZqBvYTr2vtqzxit63MCGbR1PB+lj/0v3vcfyoJP
f6uLpywzy/DLUoSTFCX1zPqcoBjICFsc0msjX0kfe4tumnApnJBrrBatpISLygtC
/UkcLd+J9NU+Uz7FHltyAJhpjgBVBwrRjk2eN9ZYG0Nk3rhJPcbCwEtf2mC9jeuo
pUS2I1vbLcusVxjQWm9fExnqrUtXf/KsIreNPvbt6VN8w26AEzs0szr0Ktu+9m9+
fEUREx1JbsdYoQ0qFLOhaBlufQBFDZQytb2E1w73orpTCIAxCSL8sOmdl05DAjiu
NnYjAK7omzkP//OKZ3IuMnY95x7KYPScvyMCWRWkdhjFyJO6XQCVDWNXGGpmNqsF
JP//oH+/9SvVM/UTqmRcjC3aLuFj/9GzktusJxg+Jv2/Vn104DbWL9QIDyv1upUA
qOXGoo5JmczqK5CYw6pwz8WCzydUACW6MD64NsEMyoF8BliyZNXfaanu0ScfKxw8
wAvYVDYWMb72fnF3lYLjv7Twxh/eQLSZY1mCi4jy5BQmrb4MvclLJFJnymtvMBn4
FbibYjfSzV1QcFOOFIcnklGY8TEX+IJ66l3bzWBwqitXOSk4QBfp+2pr9IHqLRda
DfUPmvqpku66/dW3SwfXFgsTkAFLv07M8C/3pKcCFFZKOUSxu1XKZH7RNS+byrRC
pWit7jU5lhclixfzpGJAelPr3mokZ0qcBcED4Mnd51OjP31MyneCeA2vyqua8bio
TqIbPL2VlrEMArjc2Npp92GT7bPbLm+Q+lMQsTbenkMgx1covkHlQIZS7O5vXQsB
N1dn4j0dnD3xaFzsZ/FA+COUVPuBPHd6otxSib/g580mdQ3PVWV/JAqy6frPa9J1
djHJJnBjScwAnm+mez9cM5L0+dfmbtzQN6KIf4BTcJTSEwCjt1eJHPtkA61VuKse
SE40xrKASFs+H3aBVqXqTEb4Wo3GkvGnVCw2wW6d4NZKHVwKsR1Jr3GY/GDzXtGK
+1DOcWFsP4sWxqDtvzpwlUDieqkdEMP854yybWYHt8fhhC3OhRQoutsIH+YkucLL
m8R7N9X3vKVX3JEH4+hKXkhtDgjnfeRADM+zyEo4iJJWuORM76/UpJE0rLD3Ms64
2gkrmIO5tLfP6DhMo/puHwcMD8ljc75m1a42a7k0zv8pDM++42zdrASrPqW7+ufo
lOxm6gpxypY1QT/Q5qTP5VIIgBib8Pdij0CVGWi9/e64cjkXQB2q3MoRJrR7ViUM
aRsF4t8PRGWZ7+IXJVtfsqyAGb7Co6MuMYT5ur3jWgUqvHRb9G0yhP0ffpHCh2la
+1T8/F9bgL387XsilLMaZYohRsCMmY+yCytp/dnntEDVdTnm8QdHaau8eaJO0D3X
wOGCvletDlP6J2EPiWcvMojDIVXzFIjVmhHxMKVaw0RyDL8PMcJIK8n8bH/kusrO
nreHpLuZHOXzwAdtbMlRo0w1/XSlBY2BHxO7TwJnpzfFoHVYmG9sn4OtgEiUmyza
bLyvAmG7+5easlC06XleWp/8Q+ufoSkbxwVhlB8VaxDtpGWhb2DAVWAclhW43nPb
GqMUVL8MtWbzyn9FIrqWcUdc6xOuAeYEwkNgUc34eH7idlZpq+axb3INs5Djp7+8
oRsvcEaAU5AF+SfiIhFSXtIr8tsBtROOSk22VQr80/ji/80Rr2lDOEtX1/5bVmOd
OFAwIeHaRJZTmjZZ2hqePw29oEIxhfIp2bUmEI9yt/5OB+s+58NJ0zdAO8NQJINE
UlHHLCiww8J+uVCiyY391DaiOJmGY89IIvuj31iDXzsB6Fw9jzuHidVF8c3Fpvqp
rEZST4c1nl2Zy/ZEgWvrW1IS91eovB3/79C5pDE+kgVFoRou2RvNk/Y3biI4RdHS
nWWGCvAjHbS+f0ImN0KZg1OhVEwwhtU14R74Y6yv9JX5ArDImafXRNZr3QWmrYAe
+lRI5sFTokTCdr/Azpc+BXRaNFtguOwIJ/rltxeDd+K1mYPpH3mIYfnsJon0rB7j
0GGEPYQluY7tEu0TFryFZomjuxuXwSvSXmbn6S6UN0Yt6atQzYoQGLeEM28n2LlH
6qDDXMe0HZNLXqHA40d0dilNMEH8bXCjmMlXcLYqSg5+dNNNuTACJJEPALPkEKUV
if+HRveDPHPAYBo9qYSDDKL1ZXbcLx6CZEpKe2J8vrFy3Dh6RgpA6XQqGVbZ0L3A
f3DOl+qKjnSABpA8FcB0BpfRkvh6xb/0OKmqQSC/uZNbeHbaiOahpDvV+1jnwoqI
YvlXHl8drRa49n7vQ6RK3wZQmRhV7QBPkN2CDaZc1pqw2qUte7ymkntuoE5wPOQI
fmBXsw/O3TG/+rMyzAUCRZ4nGbIr3I54moJtatXEJNayb3k5THV9qa+YKUL6NmxT
ouOsYhb1vvRxOMlPAnlu8RpeBVr5heGeuUsDEks1kEOWyEqhWz8laP1KZ95TDr+o
tDrIS/9JYGcGUzH+tRon0dDw/uIsc3KljO0+vvLQ3VfZNZ1yqGimlh1u0NlsRHG2
5tLkRpxX6WuZFiOfBrtTAd6qaowQES6ZGXQYoECaY6hGaeXDTidfy0Ro65IHKc4S
X/tjRZ+3RaEQRaD4dvFVclCdjDpZxrHAPQwrSu0zXR86IN5dlFKDjSZoQGlNd1CR
agWH5METan3COH4/2M1UFB8Akccd2rrYF3JX2tANTzZ1udKwAbRKOjgWS22Cuvun
wPYtPfyW5r6SCZv6BPatEXjyeAkNjOsrScYzx7GpdOh0gwBGZW3PkptN8glAMHvP
oPZIKGgm+fz33Eu22Tb0K0wqigxikmyDR2f1oRxjz5iYM/8ADRse9WGOYCPI2J2p
zJPZfzigSbgsfOpjqQK27vPO383Pm2sGaizo86jam+YArpNgp8lI/83JYQWZkJKO
csG9kX3nV08GtINfePsOggSAmnmSEaamISGtyIFBIKjKb2VxutSSiTiFS3qWGJDd
kfHFlM8ubFhBU56dQu1h5c69SCWsA27KSvwKypz7tpa+ZaNNrYrgk3Oy9NnJ22k3
LSTi/2tduYLv/EcaQ0d6BBo7kWvJ5Twpv4zw80a1AmowSoSAV2tsfQqCU+I8pVvz
FtPBOn8gT217kVpyKGX+aW8KKQSRj5QMw1L4gMv1k1xdRoPaHZXNM2ZuRJxtwudC
FNu5D7krbkn0xzOmooApOrF4ghraLijM5q22zIfY2lTSuLvP5I9rDJW1+OSPBqM2
E5rMUlSpbT3ZKjs9SaVJQMmqPgvkwZAfPNFij73fkS9by5t0hUuWte623gpkChKB
4OBPOeq28gYAHKuce07qqO7mMT6SntV13ttgEvcnRRmMhJFUF+soESZQr2EQSZsE
xZs8SDrteP9lEt5QNT57O8Dll5aGYDTjatTKm5ix8mMb9wQ3Ak6g91BqLQmgeMv1
COfVBgGff9Fl18mfqCHBSxUBUv45iY/t3No7vZOhebX8eNsTgl1dqOq9TFO3Wc9V
a6I73K4gaHlJrI61B3tzB4AQjh9zAUViiKAAc9EijA4cXKqNcWxv5d23DKD6p+2r
bil5+9nOh5yCujD4P0fUKUy8bJQWKWboDRymGHxfOIorjCRuw2prIMs+fD5Ssher
2GaN6KPJ4nRJVD4fY7z4wuvKczLew6tlbSEYJr/aLAUJdjYZjAAvjpG+OsvklbzQ
58HNI/AzjuunUT33F1Vd+ayl3QvyPc/8MyN9SFRSW2DcZ+GQIe1FdYHciteVHDHJ
Of8pNVMWy9VJIW3l/Gsl7mTniikbyuLHW/qddjNJpTpCZN3vqZumfthe0sxLX2bW
bpY5aSkNkd2f0HtqTFooKN1/H5Nrc0Nqz/HjBWzbQpFCeicZzTgR7OA9SoSbeXD+
9qpUrDIt23NP7Y6RZgSaWxO6pShiMp8jnjyk5HB7GeaQrd2R4BllSj24fpczL1sJ
1gcabcc8L7IFy9Va+3K15rPKUTxpAt/3Lccm90OCkkxJyyS95T9m7IEDZLmxBD4A
mObbir62HDUC72yDEJQ+lS9VymhOTVAzndlsaJIIqyjg3Z64w/gipJ5HxBjXEZz+
8UNU+S0ImounBiH16CxbOEE+H2gD2X+BUxj5QX+Pio7LSD4olzT1cVCCCaL7S4Ns
K+0KPfmkoygJfyee/Vip+Xhb/Nx0yJ75Smiv6V+cCuBUqsvnUanGslt2buG8CHdM
NPEpvPnyOINHOai2NJnJYoiNGbVJ+OClmznumdNMyGMZEdgL2syCAjTnR8igfbwb
Cn68tA/zKpA3YL4ozPokVXoG0d6m9ZnXcLOnX4csjQw975bUHRBqAs7CyOQUKaDb
dl6QO9RKwvLzSXLhGaClqwvk79FfYfz182bk48GITzCan2sLQ+tk9CLgcnXu5rKP
yfesbl8t4CYFjm/T3j4khPlSxEzpj5Y/A/yGm4+pA2jWIjq2s8ndSKsudkfONnYd
c9RAL9HB0bDmElteCaBg3s9uAU2H4BBBIorVhzq6IhlMTACJ6Gvb8mKOFP2H34YJ
SS1aDtS2BAVYfjVma5YR4x7tSVZdIT4QWi1fXTolFKNC9sFGCUC2eiI/hI6FZcT1
8/QDRiBcqOulkPTvyTInFM+mbh4iPaEFWkWp+Wc8efIrS5mU9b3osg5BVKTDBx3u
RDMJJ1MD5Qn8xyGtAKrPc5i4JfVbTzLtsVpM7dnjocO1XqPsRGmqrPceeDSWDYo3
YHwXKZi5KxEAdiff8sQWyU2yO3CIX6pH65/ZpMZhLWnD1AsJTQUiORGLgpJlmEQq
XNDoyDiR1BMIb7y/vLKAFH588HyaDqWWJwmJ6h898QBwZlv/DPZuCRaL8zLhPGTn
3u4tlZmIOSM8kTnQMn+LUHvie3Ob5i7nHI9mvmAcKYgoIh5tQNvr31TLUbNBJ2dM
KA51PiLgURor/CNipPKch2hf4w6nKGemRkllhBYkiX7ktsAfmdaleZGytlh11jEM
HuqaObbmVgXeYCn08HRqlZ9Cx7KhXxgN/jaWXsx37AB1kGZsS34dom5d9JUslprV
ScpgavxQgdzi1YVCY+y5Pg5j4pjjrtw2sKueJozMT57q5xumOkdkjCRvCuh3g1bG
rarwiVQo7fn1Mj39UfR4DHfmPIkorWuumk8s2c4d96QUxtXqqWJvWKlhBoR3Kmde
Q6UUWAzBsE4DKUJ9iKAL35UQjarcNrtMe94DVvK7KvrQx6XwBllTzGWHMM9hdFyJ
+eD9uIWzn2G+JZ2u1vc8qkzNMaXc9k06lIlxWzROPXL4QjNI4CjWyam+Iqwox3Px
5FEdsgd4fdYFACgh4CI30F13Lm2zB6K24XiuoD+UpZszK2vzgrfQ4+rHq8ju4CTM
3+vxl8oXsH5ZQ26OapzexYcX1dWLYEsmxrxl9FXVIpGPTwdcZkocOALNc0jtZE7D
gr+hOCPQjooeFqD3nSWrK6wDD1M+myrUTZXUz92XwXzIbK7uG2V+XCCdPJ14n9n1
5wFfcGqzvlAjujTnzU46tRo+WjHDadWs2zJoz+/VcPzsQ64vLBZXfq6tL1tS/WgS
L7/QF/Z7iXKxrj0VyfKa2B52AbqiDaCgKndivImyV+3h6AEzZwf/EpfwoLFE5R3w
dHrsMk4jbpMP83Dp9XXcJhlvDlS9nRr1bvXpVyFVdNZpUmNxo2IACMzbCacInhrW
XpmLIW6OOXwhyIgBxDDaecOwQ2UJDH2LwVyTttK28jbx/IVYRNebRXpqHNL6yfkE
TiisjWrNCc8pJlW/EQ43e4pGbCGtlPvp5Odr50j0x1wMd8A2X6k9Gh/7VyrTenvj
hqsQrkIRotL4j8usVBXCqGzH4RX2YORYygoeepNzc7ugK9Gv4it/y+kg+85oa+Py
g79faZqCAINuuv6AV9P7mNKbYqklTu8BihfIZ8xG7D8ftbXBdtqGYw++ZDuJaYZM
KOZGqH5lBzpmGkF1Ed4y3h+R1jaeSaEfHsDnwX5jGoNvptX47ep7WKVhanwQHZCL
4wkRW86CSBwunmaqqZaFI/G1zKLa9SqEutmXV+K8jn+yQcLNUiC+gydHZdX4+xKT
xTW/ys32TX2OMdVCNOqu9X28gttp6BeDW9zPNLGnRZDgL5y2mvOE8wtF5ykrU/f0
uUm3wNUv9HBcwBeKIUVZY3NJYQCzZNqHlSoRiFzGKiomUU6l23LlWHQSkxggfw5e
c3g+hbxyVap0YUClH7SRAhEFxCP1MwOSEz4u7xARyeragNjD7p7PPgYOnIbAH0T1
83hWX4dp1HUEErZrzhO0JcZOtt6eCI5sU2Ju1p/EyRT4NywtOrbGHNcMZEifk+Vh
ruPnqyFyedrpPOTZrNrRfEgAT7HhW++8Z21iXfok9iS+VttAx5jpeVx2YuPGeLhi
tQl0VsGPgWQhUKLEFIGLdH9vPsCxA3ihSC353mCtDhNroE/EyUc0alWfnvmuo4BI
VBZojdanu4i38HVwo3xxSni4rhOLcQkopYBafWsaDOivzWY9aoykaDK7eQ1fky2P
ac0cL7vjfevaqHYuyG/wnfssJGwgKPdsQ+30MN/OiQt6cIqtcGYxdr/421cANazJ
55A077nzKaM4W7Q+PWCOFvr88KmKWZ7sUUmSyYozIYyR+xvvHKn31mn4OMLuMp6y
XEBLZR0aCLTGNRwu4loIv6XezXq+qMb/oI78WphYrM+nei1MsWGQb31n5EdWVN8j
KgBAx9NZ8IpVrysiFoPZV1MDAZJdbIaeL0olBj1LVGZUzCwIfIRWiYPJHlCaLU7h
wUci5EMsE2CmVTosjhnaqMYqt2FgSVvPOVzyEBYnRpOA9ozF2YdXuNblsTK0k9Rd
VyTawdLtX102ZNdbuVv7Nxb3FbiGQB4l67dbvO6W9G0ryZXmEYWYtieDwr/MpWno
9jyJyosoWnoTZaoniuXrC7Tujll3lwskM/TeGBbnVARPs8A672U5JwNqY4HLg5R9
WoMrFJcG6Yi/QUpoZ6uZk8dHhfy5jXcAztUXnaO1uOBjrFH6qtSrHaIH/pxYfkKV
pbhDJbhcEPyECOUsUVJzie/tPDoagzCDJxLLT4ebvrdqlccOX7AVzitm8bwZFrKy
6T26gf5xh1niBPB5qAckfMCdc4slgcotKgJfWSIBtZH5F5TrJPHn1p9FawcyUdEw
1oizDsaSybur53YHOlah6Ki2UBPSzOXUGqqLZxtBMgS78bVim7mQQ6uOWIi1EpWI
agiqN4qK7QlZgVj1jkDKQ1fpc+DjEb58z8cUaHMvW+7I8mCmg4qrCyptWhEg615o
3wQ9DFWOBND2wuSPujhzzA/KrFAa2JVNqL4hoN54dISd7hNci/K4jeLGiyMcGKIJ
0Ehdytmmo6NU5RD74wEgKQW7Yt7l/Kd+cJk9A5U33nTd0J4pR8+6I+UGP21cegWz
T59fIdPEsOjgr9UCk/r21jPe1Sn5aaTTCtyBpIb4Z9uOVTgzDkwCiw3SLwPdBSVm
oXoleyU48ZoAPL8Clvix/jh0hXk3jiurddLz1DEfyRuBdOWrnu3WZyVNZt9mDO3a
ML/FHm3UEnPmfkhC5ixWwsGX5KlgUDHlBZGDSUrpmsSusw24A+Gk5KcofaocJwuc
3ue0iFr+3lHTU1fA3MJxfmcm+yESfZaVLWs08zO+N6EVihhDpspaKiOvDX2s8yZX
4KbeBXsN5OREn9pRC3ROC+aj2wGuOWHzeAGQgXHrPgk4yc3gkEJpjCHcyb2Dw6s3
VMmC0yENgCZDPBfFYGopZDTmtAI2Mp9kbH51BXRq4syrWAnYTPhZBwEknCpBQ9gM
NuO/NIHoDdrfD7QYqZ1tWIMtZvceM2+4ZDN9AmsXAqbtXqrGM96bmTnsfL4Gh30C
Ph66CabRW3CYLzUhsALpIwdzoB7t6fhRh48m0ZbXE345pkTF6cE+Q+ghFfj3h3Ob
j5YBq48fsq6yW3/wvGZlVT5bDKVDZhcJFforc56jRGsxXvap1DBC/PIfLThmz585
/k07YOr64Z+VyRBYTjqlRkILLZCH6mImSXMi0u66laxEbsa8k3aRob9oZmn3JSWZ
j5lqVSJoDA/730cMLTuzRNXHoncX5hZpGS1nMrkdbts+idLB8gkqirNXvPLax1rq
wJq477Zo5ERR45eLtfg0RiI27a8/e40K7zmVhhBdV8jV77sEMeMSdJMCjtU0Vt0b
fpK9oDcIZ5HTK3vWUHfCqAtf84Ep4fvQf/c/noEV/N97vdI8GbC68xNb4dqRg7Zl
pb3/PE141vamuQu99CjXfsmTWMRciKFS6jUFclrfOSY6nQvx0H89v+LdF+E7aCRN
RVmZRRaiMD8gYAOHa+ahTzNUBDqdaGSSDtT98GAueGVMj1pZuRJgK0E1Rr5qFTD7
trkmoxc3S1F+5eK5eEwZF6kB8H8vk9RV0nvjZvJKkZJxz00+tLQLWI3B45yRWFXI
T87MCexF9FRAedgn42hbFPRrzp3TdmL89jpgaY62n4f6DKbPi84EdlECzHGtlOin
Y+il1Z0ln6ICRuFMK7zAQW+xrzPqAyjMqe22pLhBAX2vBDlRLFjy/lxHdJ5X4+JD
22kiakdRgZulzz26zitw31aoZMPZZhi4SW7CTRlcyBRXFE8qzBn/n1DVHoIf1Tfj
vYEELCHMXsnnH3T7t1LNFo+Dq+1rAVs3WVj3Ddpr+AamPXImliO3vFlxYYEQJO2n
Zz3ipfTDnfz20wajFiHcEu+U/MRJssFUXZUgL8JMVkGmyGMRx9/4aaTNRUZ45FdD
nQHvVA5I5+9ETHu54O/x/Ei9eOu0tKrqY2QP5L0v86Gi0d317+pY6cCwqeduPXE5
VkWSyGe79AtFPtygK1qvKMVEeRzaqBoXLO7vQ5+rt/RnwZXvOinoeRan1qj8A/Th
DnmC+ebrOakCHUAWMg19uR5cCPifYY0RWaRvRcf/78PL3ghsNHsmd2f5uIFB0M6s
EgioVxsu6ubKjdYZbFo53Gfz2+IsswQTHbccsVJSzUmucq86qDNA3lSoWJrA7TVG
z0c9yiSL40Z4QGwqmY7rjncJHBLDd7+XW26xxfbVa6BUbWr9XrMcKyLFGJioxQMC
D0924T0ezuGFfEBMz7rz9SrshHSRXvdXwg5RJ7o8RbNbs1u0ZLv6OO2BP6PeQISB
2nnZvc9QMCF8nYdhsfUJKTjNGi1z0S5PQ1fS9jGWQKq/FMMOriep0gWxIEQoAk6f
qTmyKld+aPeSPG90wL2v4CgKheBSVyG/7w6oTiwmEC4lT/GgA2BkbOEa5kkT/yh4
UEpRzbGerEDaGvLWWrgoBkZ2UMV+W9z5tprcinL37gpaunczHRVj6cbm1BqJjuYj
06mBnIJCGjy9Z/w8iSmYKTSqxEU3/1hG4DQsSP1Mb8N64j6ppU2P/Q0XtJp/y5vK
EsZaCS+KlPt39mZ8qAZYtp2UhMXS375J+TkyuRpYoZsAzsGmHtL2H0Xq+9ZL1oo+
fBi/hI1CZhQ5m37jW2kiSWYDpXNanphA5ny9L1eXtCRelxky2B2GsAon2sG+5CIm
aXURkg0hdOPUNa8maiwZIFE9MicyVvg3XSgyi+JezP0FbJFPyv4DJgiZE0GkfMfP
23MgIoHb9RXWlvTypjBktWCPwy+UEU/w0jOlwMElGSU/Jvhpg5Lm5BzGczu2MXi4
mPJtWeb6kTMv1XiWTcqjD13nvt9BbJCaIyGr9AZzdJ3Yqz2IsiOxZbMThSJ7KcYu
jzMycoExnhXQqLkSFzuOBhqCEkscUyu3ebAwo6G+HTwMraVaPb06bGRd7PewhvEb
qjUnZASQEd4zNKw0aD6fXWhhHHAPUEcPWVrJoyCTkaxUePApdm+4i5jbTj8rCy3t
Tr5xT7wshZYeGYL2P08YPDpX/F3FBx911CVdELKzd9XyR9yWgTQIZlJlL8d0uOBt
ysy5Y2PHCUgH7YZKlPhLjfQfbXjXzP07PAV5lc76Zrnhf71i+dvojd5inUvcwsvQ
WnD414uyf6slspqB2qcOOt6/+OvBC1EWW5p1WC7NEiKsa1xPm5PruAbK0b+pISMK
KRKuorDJW1ZX0Gh+NMdq5sLCf3KhXqVk1KxlSTRs1mXBRyZnyX/AqyLkkhV73UMC
2cEmVg09/jr/4yJGmvE00vGrH6oQfAaUV132ltJVpDj7oHDY/16358EVS4XDmDgj
C+Mo91KdlmO18bf9+ZMwNcCW5OPEyS6Mspn4Votu8OH+T7eL6D3pB1JSfgH9+WeX
r9pB0gl3G+AeVIQnuEqN2S8ZW08++bnwJM4Gtxd5OJTIyfHRlMvMjgsWXbDJN8cD
yfcUKBA8cfnJ78RJElHFfLjI2Kb2rF9tDAcddizibBQdPdDHZ6PiNRj9XKpRWNIT
d9+1FhF1AJrANZH+MwM3lbjgIG70RYszg6H2H52HXUVGj6r71H+ifjH7E+TfMfxg
ovdtj+Fk2f6zHitynSra3vzXN2mFsI5BEocGolcPUKHuLXNxnhVW6tZjiZMmSb2J
of8aiwck6K45RoUj5w8NusDxJ9skKYeKcAK7MoaIqdGoDqYlDE1dm+nqA1G7GhMP
bZZofs63j58Pla/DtK/XAeKm6QBKXcei338KB1xUL1ahdmMXTCVR7fGzjbOoewkJ
m8/BUFuPqbryhqkufW0P3TJZ8S+uKsH01QQwpRyFqKjRJ1iY4SXDYhs/t27nRK2V
yJREXKIu1tL3toQ5e9uX2+x0qkgp5Wzepa+1V/+spCPhCSKA7thguWV3A/GvZr3G
bJLTMbAK9G6pD4EAwr0TBOYfxO3PtaE9iIHp9XRjwHsEZMJ0WfXlswAiMBDEnTbp
2Mj+IorChwtZjNJj5kHpuuOMS8/HjVuSfYhcy1OH8gJbU5WyUwsLb6T6hhOW5qIE
QjDZzeISCX4pdMxs9On8rIKlECvp6IO/f/kSd22noCQQ97YCkBrQsUS17l23YnUA
unEG0KtahaENgzcUBosYavJRhzyFMOQGhUpCN/wsPQeg0NQhmKquIUvZG0XuXlKR
9ye4OAOtE/ZwdDCMm2WF7cEyjvCq17FuOGOIbsD94Ki1hNcWU8KevRbxCCluTFLC
7dGyM/wKR0zPaQ2BzcitWZlNEtEEt4a0N/6LLDXvXYoA9BbjcYCu6SHY3WfSVq/r
7r8SyPiR4u4YByY+vEkMJ60oD19nP0V+tT+zfCr3NWne89pqGQq43uY23l1+6KZj
ZwrKkjbWlYJJUCwo4+QWLlLPdKvpI/hrJlojG3m9bvRD224ssUhAAbJaDzY12pmX
4zR/+2N0V38HaR1olYenHm1mweLsfy8QE991XDIpQenN8ZRE+2RxGQM/5SDNSEPv
1OUM1Xli6/k/Ew9u9vNjXwKSHDk18ZHoDaVgRltBDVu5+ew2YKrqaauYHwfi62X5
evzReg8f+Yo1mbBpMqenphsH9xkoIvTQHMfws/iGPnk1hqkq09Ga/Z9bB0grXam2
lLT1pV3u5JL70Egfd8k4sZGXlZF+1/u9AoWRgwlm1nAeT7Mgevp74J61O5AkcKe9
Ec5OulNTq9AkdRz9mVAYmhgoxsUaAqepDCDuej5pDy/qlqICrB3+VleeOie8Qi54
spcABXonI4s/Mb9NmzxrO4EWzxp5EOVVJxE0XYz5cc0UEfJ9UMqEyCqR2zZdAp4E
GJoPqMcqCI6Oiq6VkOJ6l1GqnitTtjv3UW0MFwkH2VARc5I7+x0ZDY7GhoeyBipu
YKmBhFxS8U/xgZTap2vXooc7vOxJ6FvyayxRdHTeebnBel0jeXQGJN0piT8r8PtF
+BwTixqZ0o5tKRSeW5UhKaqX8kPUmDhuWZWt14BtzzxydJzSiVUWeeKvW6ySTi56
DZNUSy8E7L5Uo56M290s7sTqMcM56eR89Llun9ZscuAumCg90TO8/+xszjC3g3Bt
jap6J7bpY0DtulWe2GtvmZ83iPlUZ+XaKGCABfJfZKb8IStTRjSnXu557yDKYgLz
9vD7yv0DsJhIzZe0zYMRz58nX9ltXQ4OoPWbIzPN5bp93f/lci2/FYqx8p9GQwQe
Ieu8UkOaoUrKZ7VZ864UoYc1tJIjXbxctszxoZNd8kQ3BWR7xcRktq6C1FCTM/wU
3oaj/Kle8qHjs5mnUjYM7yaNFO+k0S7J6cpNqo3Um6R66ahfFZJB8FseaNGxlUD3
2dzeDda/Yv3p6pzgKaL7CFciodysON4r+bh0VCcQHTnLDQm0ocX5uXgCLpWPV8pE
iy1IZptl9v8/xKOPziisWkvarjHpB65uFR0AQPMWLh31vfqWh2HFyGiM9z75IIF1
we7RuujLUiyw7jnxoK7tRf1pqbWPqK+9ZAvwEfGQjGiq8qeKuf9gz9p2iGU9cwhT
sa9akhooR6vBy9nJDkF9R00eIQ//d97UDtjD7PQjTSB/37hGAPHJm5BccN9sOOYn
FzNJFpLCc1m4ddob6ldBBAmnRRLLMAhxF0zUm/qPvbht0BwAZqFINw8sxzkB3cx1
o5NXrqtkhgD0gZr4PnMywtZC9mdI4HdfFsef6YbtV3P3NypGTsN5pXFvxFB371sD
tZ3A4+N6rBS+My0ocvh2MK62d2Oi0uBTDJx0W1l6WoTIAzM2hFDBF4MzU2PT9BNR
4ghAn/tx1nCQCyIWX4Z4X0goHDVzZeJAbc8iofMsszJ0rcD0AT6YCrrXxdE5ohVr
kbj4zw65Y7JFD/M5SMkU0Qdcr1K0Q0P79j6aRQTYfCIiPYlC4FRnxRBXpSaIyfdO
h4nR4NUnvkUcIpl60YQNc4cqdNw1Z+JFNSFG4kDBkCXoOs+AvT+pzKq5Y0bL85Op
ZQs3gih/peWBByVYFmYo6791yU7G/Dc855FnGoGqhK3O8MA+29Q7U/nMNcqQmlPw
lMap7HUlGTVxWmcxzo49hzjnuFPIdqYyZg9M+Ys+ej0b/hkx3lg6XK/j0lJnlnMA
XmaagGxnwCo+EDETDLe29ZaZtMqiz9f0o8QWVP1+oAZFKnC+AIWgrRJvlku+Kz+W
aQPB8Ck2pKR4d359Xstokcn5jeEL1P2q9EI+f0A9OQl8lByr8nU8NVcaBojEIn28
SD+nCA9Ti/qHc0Ea3Wj1JoVJJgQtNisunUdnFQylsXwlghSEEUMmEnWwGSAyY7GV
of3XY/L2KWomaskleod1ftbA0lDg8J7qjPYdT+utKkWvxxthnRE0BQO1BcQQEiyf
9acjJjauv4NpFVn+UNGsgNFIVQewnwq8GBnjBERww+ZTZiEKT95Ug7voNIKesZoI
uTzF7ne3+LdBH2qqHBXrUxGD1tjNu9Mk9R5Z5QDYFZGRV1JWtvST/v29JjgpbwpK
Q+s2eQS0AgvDvub6mjAs1dqLdMv+fJIcsUF3tabW3QuIxbkJi9xGf4vn1BjuctKT
Th0kOykc0OSB5WIaJTYOmKcDiERRbKqLATryC4JhbYZaw3lrs9VxXEiSTKxSku+8
ZkfGOCX/Tiu9l0xMSf0MyXp4qR3B6x+fNB2Gqy3Mk8WmY/3jgltURYTFSK2quotC
GXYhxUb31i5SGsc0A/e24xu541b0BjTiFkjO65KT8QijM9EZMTfww7CoJZQ1V94X
ee53Rp2tsLnK8lmYRr7v1osBQn6th9SjAB6YUDJfrJipq0392Dx+ATrHni6/7gdg
Y3IY1guWbjKhkquFBXbCPy8rsymJ+FotXlEPVCW1JMB3Jt7M8mItYvW4w4DMthbm
mMOlsjHLPvaDtCw2VI3UA5pIf1eZ7mXfxRndPMsuDU3RS4NkGPG94QcT2ub1KIVs
mKWi8CX1NQs4MKQTHqE9smUjNxq1XhsTPV10SIgIWwOVFMQLnyM/AYSuS8iX3A2s
CNV8U5D0+QmaPFgHXcpMuIPL7b3oVAtX+Nx7VY55PwcPBQL+XcFIlePnlD+CXUpA
IOZCnISu3F1qUN1qmpLJPUAZLD4E3cAEATAw1g772Mzj1Oc2l7axKxO7cWugv1u+
wwAu/70h2LqrvuZ7fBiYLUcntSjmQvb9bHkleg/ROBVpEGvpFS13AB7Bs0oycTFn
NMMY3h4OnjgIgySKGQBKmL/E6wR/TvbCJzFOHHeXSsFG9rdXuuJS26at7rDwbtun
LfmmV6acynZ4NXBu9YqqqirSATRhtIAiY5uD6b5bEjih0KGGWS3a9ww1IWaNiHqU
Ezi+Ms1ifXtmXvjYXRbngWwhupeZwI+KUbC9sOzS2tlOBbkGwo7AqojAGq1SjXeL
F6V97zma+7S0F88OmNPJsbYcR4X13pt6P5o/vMkmoo6e598USdnxrjUdCYYDH/pU
jB8eQ4sPjtteOvLbkH7hn9znjz1IaFQ3OUTh6lVJxosM5SjViH3KeQlZFTidXZ+e
b4MD5Qw4Qe28haW5EavKxiC0mLd1w5VQQ8eMipQ4/kZW/meUN6K0kRdm8qPZlVc+
wxPesrwV2oNd17TsNgm2UEWx7RkNSAYiYZDEYA+gGqpXpIc5HYHtS39c0vYQe6vk
QjJSiYMza1LqYufViAwf4WKHIAn3tD5NWNbHstV8kkzRj4FyR59e2fQcG0zuSnak
k1yWoGs4PdWG8xknnWVyZ5kZRppPzx7MWEdySNWF1VzDxZtn1fDIuoL7QwSO3ZsM
jw7A83QPpxeZ3mOg4bK2ef/4NG/QMOjWONvIZgOWv1uULtC31YyxgUOvz/qIMwU0
n0r/+Piunx0uO9YNmB+3A3N4a6kkmbsgZEfkAvpwL6XPp9S8/yDFa4HNF8OXL6HC
eku0rLQwX+ydaCnyua1aZwHUQZBNcpsvUkpwVdS2qeIO1OKEdn7wZY3M0ekVmc+g
jkeeqHk5SyQYn33Gfgw7JMqwXXnnOg2abrPzZco3IASAcikc0Hcv+hLWOaey+EhW
+1yfFrms1T5ryufevg5sZWPF6N5io3x2ppxmh/DDPvT8JegVb7LAiPJTwRvPFNbU
hzz24uebkCxUKZN9coMY6VeWoJ8eGbnakfstKt4Ds6FYgYQE5/ShsZqd7mHhdmAW
DAeTYEeke4mx0rd+LrWZwjn9Owukb3nZioWbEwkG6rPC8uTG/6vtt1v2iv30Eo8o
WS2LthAutg0stLjyUNZFI7df/szWfbuMxw5wb7ctVrG1OtRuwWdKrrJ+haByCVbu
7EoDSfBwHlwrC+e1JFIyuhmqqpCFc4DQmxNtLjkMarnNn7XsHxSz1aeRgHU05hsE
zZ9C4tzDs+rksDQLewvhxQVTlnsUAM05jdh/tYqsv7I/bQOXTCwyjoVw5/HdPMNF
NP0xzwpzSNBkN6ODdJiGHrV/eCxZR3pewHEEVA43b0ATdLdIxwf7/vZEBvhz7Fyw
8aLfsooK/P9zBJal/j8YWalVJJjF6NWI0OYB/D/POAPyeMGQhXuWf9yn5Z+HMPPo
n5CPseA1ZuzP5A6oOuJmiyA85WbqTXZ38jLQ+fW/iYf2BO/IYWaW3Evn/ggPnybX
xiRoFn4EQ8VLDiN10htyVXISXD32FZmpedrDWAiH3qy9awGo5oZX++AQYaIsd3Zr
Cc4bC2KLns6FZeNeSscz0urnmMKhvG9EkXZUlCcV2PPzY6H3K4BZmrdoleEUabLD
BbSQTsmMuMxSsFG2yyMgLR4ns9HjmJgLl0818sySbXoJnledDD7GeCLkDya6E90j
OQcbe0Czum1krcLN6ri6YioxX30qhTsjeiTC0/nCOKsOMV5sed7/QveL1LmB49RC
R6C+Eh3scgs76pSrGezIKNoKXl0geLdnvAwu46Bj1pfwvOzfpMSSoYsTnapb+J2L
Bo0AEssX/wpLqjv+GrbpIdCtKiWYsoUH5AaAt5NaDi4+oTTwFoz5TBwkQJubOOuc
8U2j4UkVPKzXUFAWysFAl40Xmzj6mzD/a3nVWvkBN5SEFKchuT4Z+LsYBNp9OcZQ
9PJhWhRXXxerqEMbNvh8w+KBRX3sMx9FfH2tDB2imSsETHnZ6iDbTfnusKQCP3Fy
g6jMGlrmAIj7rKmQE5iL05G8EPNCpG3cLcFTJO98VFPzeDyz6bsxQENSDOxH9ND5
IGeouc1EienYeVtsDjGnmhVL7sJpzH8KJ8uKpRpPX/DvGFbuSrMb9G2rKOW6k/Xu
CCjQR5o0HLWIpAdkDYfY3ghOFQ+xLn9H6hYlkeisKQldc2nwLQPdIvVL/TKnpjuZ
jz54WY0hRAIKXqZVfhZXXb4IflQ4IKcEMJVBZOPkz5IZ/yl9orYbbxp423T2mGvv
Zbl3t76ZsSOhPiGi5qyp59L2oKMEDqvB1Y/DrA8EU5yuNZGHKUU4KIZUa75bHEft
34cD8GB5zG8mP7313n7RAxlxF9NNmL3qqf2tx+0bf2935+pXu5DVR9CfZS49nKNh
+69fYWtcDjS6gVv2K58faAA+5sS8CK+P7vMzAksgLjah2Qf3cHPAbvL1onxd859T
mbW289RpcDw8uIc1FTVIPuwq+96AOcuWkaADhNzeiTkLcM2UNZMUjqBK+losbez9
vQ1s3UsZttq1imhjVMoeJIRR6jnWmxSVoPaIe6v6Wzk1UXUK5AaOeINX1YQtRYF0
1n9F3wXSOQUwa/i7iy10YkVxgdd1NXff4/IIFOp0PUjneVcQgfPFG+nki2sJyfG7
EPuqk1+bUoYiGdhim1zSakP0zZeP6a/XDZlzn1ajJBCd8yjTk5iIDyj/67o1JqbY
atJxaaq7KP5jb5xQ1Gk1dmsUF0LS3sNNcZUzi3l0mALzuuRlqZQpn3WK2xGbaAGO
XmhZmp8AsPJV9AerIsrQQTzaS7bCUqSutBO+8dAXYSSJs4qQWxN9W3eCEzuwub4I
tFMLeZ4BGbDw4PmmPjBCDBqvSXc0Gjzmw/BuJlMB9ykADgzUd4LPdQeNeM2SDdit
R/uKd7PJ+8jEEF/LEuih4mdxf9fg52ohzVDtq12xC/ffujeb97+OsV6oJnKHgQ0h
G2Jrznh2Ii+78MTxTGKSjeTIwlW/uoJUlCWpUrnKo9+D2KZTypsy+x+wpa4IA3Yn
WgZ3KucREcAv2TO+v31qrPQUNwNiOZNSklVZ6vSRv6lYj4RjCwAFWSDNScuMUDDd
+SzV0ufcW1a9rjqPxWpgXGfc25lM7j0LGDNrtW2LiH4f2DVUYVXaR45cvuPY//CY
CxBv9saNodw9SfUZWywM+sEdZ/Zn6PNOOE1oB3i8NwlN+aF4Nl7kVed6rv2rGbrg
HV8jUPwRhuoSHF4u9nICAinUjGro2fol/cLkSH2zmHC6lOT7dzWsLBpXLxhjiTf3
q1lRbOpkq0ulpJ3wEdSZFbSWAd93mHV+U40W8691zE/t8xxxCHa50nCBn/m4uRGo
2yOceUKRZra4uLopAD779nZJ3Be3nskcBgboKIERV3XmU5gEQ9bj2T8ZuRyZyzPy
Ria88y3UjabWkkA5L7VllWVYYmQlKXALzyn+6xNqc4oeP+t1/WLVz9WT6eGJwh/S
Hx36ooucIPiawC9a8q/xL3Y718nd+OV+naUclfnRJ45cu49U9B2mXmjN4Gnr9QRJ
47n61zA+14l0KcAhhkirRjLbvErl9fWp2AXwsY0lcnBv9J+GMyu6tlnbvcHfzbZY
YryxqMbQLuJaV0Ea54/j9vw/jGUfO4MydqxubsdA9pGY+QqamvQ1nVYS5h661XFR
EdRtSbC6zCxqI7geuJvNsEPUs/b3k99reOBPYSLyDZVD38qNURRHXOa/Lb+KGv/D
dLy/YQIZ3DWhsIMdtBvpRimMI+UoKtU6lsbPxQwpZRz/MEnHD1SvSEn9cb7LCUcS
2mzbhyefGMfHnkE9AyWYaqBevIbhJz+uTKhjwNzpOuuj+xo913fLHj3XmYSjcxiB
Urrr1lyCV2oj8rK1aeNRhnUSVGtGgmQX8nzaM+ZJiEHgohrwSZA/6mM2CnK47V+I
c7kwVyYF+i88tVglRlE35/VTuxgJEflDv4X8ch3BTGULcCtTLNLdspY45KjKdANb
+Fc4Du0m4imKFy9VwuAiEaOH+IYufv37yZlo4eOkOdOOU5NiZoIQ3tKj2kPDtiiO
W3t6+qZMEAUSJ9x1RVs/eObBQHMgKTOPzxo0Tna40aHtgwkWmbUaKNbyFxUG4gDg
RqBtKIohmcu9Ku0kWsxzt28LbNyX2JWXpvoRGDEWANZz0tY+PgmwuEhAtUDAqqsC
7SrQMeJauOMT9dTNfNmApNf8KdvSzn3710t+CiTRu4Vl3bgtjxWcZPsFR37rYlw+
G/hlxTIdnqwtxk1L5G/q5SLnKX63u06+zO2i25mXu01jPTAOXcobNfPW/RX2fICT
ls/qo9lwnd02Qf/psV3veU+j+SnUvBDPXhbgTEoeFZjecm2/FrcBTSYe7Gd2QjSY
8C5SigSi788y3OopjL2cjHAJlMY8tvLMsrIvk8gV4IhN9mh7vsETQf7Cf5NeScgL
sxMo70JQ1EPpDS+59bdGPj4q61USsRyIs7FD83map27yW1BVpu/wP6sVP73qUWDu
SPK4a1najykQIv4gmOBGyCkmkQWqDYoH4Lq/3HfpD6JhERa35rSMGnATxnOk5XOH
ov5HG02akBIUJSli3v1Dx+x4sLf6Kr93kx9nY+ZdONohyP950RzTLzb4LYg1wlMC
vnAkdNsTbqJj3Nuiaa3yLJjTHPn02faa2vg8ESok20zPh/9VdIYK3bI6br+kRlmg
d+JBvWnkEEy9B3ax62ZzTWB5oqmee1L72Jfx7CGsnwT1slJKYWBd5CO1RSknw4S0
J+WsN3PmT5X5BujqFu7ibZf//9mRbTFBEp/jRO4r3eZPcnxQMQ83T3f3uZ7nAglw
ioCSZpjuWk/QZI9xz3ri9vi+MdeXGnEOZt5mW7XKPSInV4o62hJB678jex39idmI
elGJuITiJpNvUmGvTwlMjDhxuFk4o2Gf5InQpWo01OayXs1ZBGbNkMX+GkLwA6fb
9ui6946WnEJmsAwID/wS1Oeli9pOI6TKygzeeFFqkmeuElgvkmSHcR+HFEvdYqFi
mNeKeAK9Edl0AsKUC920ITcP0jwId4KyD6Zd9501VeDtt67CcIEHTH6VqrMVSBEm
+M7onH86Yx5b7lj4I9qw+VroH2RxHXTaryzPF1I6rxHuYcjV+YEYVHtbicyFUTtu
PaRTDMTkPAoqnt9q4ORDtGLL7VrmX1bpgjXCo7GAA6DYudfM2naKi75OB06T2/V4
sPkhGj73EU+vxwvwQ/Zw2mwtimzTRSsL0c1RIjGXPPDynlFsStFADJ0jSH1RVDbX
fW03aeke7mNXWmK3ZivUBLRVtqMs/546YC1aXw7QncnCRHjVPMmV/iQqQlKCiKzz
jyzjAGMM8TvEdkNt3IyPZ/Zif7coByzkb6ULuglRfCqJ8ue9BOk6K7V75uZe7K0u
n7z4T/sof9lXYV7bb9V35FxEZidMfLo5RQkTpX3/kr7Wx0pIQxYkk4PJZofBPcCR
Ja7IIgdNK27u84pay+z7d7lFdOhXEPimW4R2b4oW4OacCTgH4DYdh5SEoNRZvocR
1OhoXawIbvJOQNkXWcTEASu4IhGzbhVBu5b4uTrFm07UVTzoau5EPJH9+QYprINw
wu1bc4SNZ5ueRQe+/JYWfI3ASuPFVmx+Px9jeAz/Ur7zNTYQCWaQf8l6wFf9ctQW
IROKzC09ZL3bQsNOd+5PN1RZDjr3lkSddRDiiu+FqY6KPqyYUeNgUSc1ollKtGFn
O7iaYjz2uPbPBc8Xp5iw4mW/sgX1yXyICu+mnLJfI6ZgqFSNaeeOGl4J7cEgWPff
kGzC+tPSc8cqID+hczfVwX6Bo3Ln7TzV+5yLGVul8k3A+pOUnoMkUz04igMFInIj
BzFvgJ01ppclAP+/W3PN+SmRKEC0oJVZyX/eIIm+kNpQcJtXsXax3z2DXLNlyTKj
kMIPUKNutGwJbA+E97QhoMI2zWcRWeFIzUVQOM3vAIizNb3HA63MWEZXbtNyjTRk
cc59vuupj36v8HMpg1f4Zz/59Hmcv1jr+rWULvOJI07Je/rfWUJRmmReNKht28R3
YzPDRkenRYlcSP/gWnE/N+XYgxtad5CRAHgYi8KOToeS0fY8Duh5BjI0V2qiGIA8
uSw2Ko2xzKfhkIsLsKdueu72/+vPBXhOZX1yspSLWVoD7GnRkmjqgokQ8mR1v2mc
sBNEXuRHmiayVZfiiKVeUWCy8iHaTaAZI6snioRUL7KZRsJU+SF0oMy6BbYeRnmi
CRmU6G236u4Mnox2UcDQ5t8+Xtv8qtBURVfYk+jiXhHZ4RbCWFq3qQhPqC10lrhB
N6JLMsIdy6cKo+AfeJeMH8joVn6LHkpTtfgnltPYaneAN6VZwnfdQutjhA8YBfU0
xylUrROy6aoFSDS+pYc4rLprJgeJFri9onwhnNxX2thZz3+uzG3MFpGlBFA+jqtF
EuL9vZbkn5+x8Iz13i4H0SuCQ2XJaMwOoCo8XvJI4X79oITeMzqTyT09SeKcmth0
WV/JbyEPMXhXxsgIwxKt4FSCwGUk0YLQY7vC8iv6HTnt9Y1yRCOeG9z/yoiAELFh
f30zSNruG6fENNe2a1RxW1K8UMJ0fvmyNAT+vbRXnfFf5pHXJ48quKBBK6zlLJY6
R8V9zMN6vv9rvrToVBjbUwVMlTfRIRhmTzLSPlnkeSp4F7s+TGl4F5Qyz9SOOfk+
mUQG5TkuRNv1hVphimPzouA/fUG1aifELSNhLpUQZ8+OuxmrXBw7tzeG1k+4wbDn
o9RXYTz4fcYKhKj9M5XIDxa5/YECLvTeIQpxEeOmqvNW6HLQIDjn3siYmK8QqM+5
8EuSNMObg1C0M+XGs8bAz6aea4ck6dJ9QaljJWXVaK3vVXINMESkja4gAEsYQ3YX
D2tw51+Ex8JZt9ijw1KwPHWYen3eNfDm55zWZb06i5FG8WVwMlY/s0z+hNMTZRdO
hWraNczyvbAQs2rzgVHlSDHn5iGI5Bzgfj9dFJTOlFKD7AR40P4tTxS6tOQBWE6k
VFsJsqWGqcyvmo+biPa6mrIkgdbFYiQxfeSPN8UozfmN6ObGhQ0rMJl9Upe+g4sx
DxT0gYvejaINY4pvYr6jfpI8+QIPatzLen0M6W7jFEUHf9cUnyvKJjOOxW1o51CW
fDqgQOMhUPPKJvl6wNpu1B3fBCsB+JG1IT1RWzmFOhrOtG0p4EP7UTDTxhaF5lIH
isZrSMOHHmlzKorFXVSci26Z2AG3A/XTV4vkLYdY1k3+vSqRjTqo41RJH1I6f+nG
oaZDeftIWOQIQ2kRGPHoQLr5AhbxjYOaKkN8M6BCM42U81dqf9CVi3C9buxp8zyQ
eL2+G1+5MLvMah4oG7aPcprtJqVbo9sfHLCH8hlZTDjdn173YNvxupBrq/cTzqf1
CJL+PwcsXUtgXVpaPG5FWJP8qvB/wxM5TccM56i8FL+cHGjoeLGTAsFtQzg2X5cS
dr18LYd6nDdqBrddUXaaXAVVdoC+GKQoFznRJkZ/KO1tmQwNdOUYdHt5Mp8TPsqn
dbzlprNoYeL82cL26mNeg6j8sqQ6Y24/6bnD192lGRg4i1ciqTChU/5lncn4mNuc
YBB1amZLsAnRAi6OWLqnO0G/ue6OVHrEasnXw6Q7Eo8ROD9CV8wu89x3wHtZPLUJ
BvGnqNe+MtG34zinzk84XKWlUkT6LCyUhMdmTlyGqPKxMiYF9XuJYMt0CfHhHAd6
I4sl1OuyCXLdPRViYsnI3bfmZaCbmZNjMnPuiJ3U979BEUPkgLKQFNi3zXO/Fooe
oupyBJDj2MDo3qhf/4hHjQcS9KDLfMKX+2jc88CBPxMX+p/uE2EzDRRaK4dE+6ff
hgMbnbhiDnmUGhjRxba5abiLFr9aYpu/CUFWoeXn/GICEHqSYHb1vyhITGQ188Hk
t6JffWgNxAnIsB3Ke6Xah8g2oYSarycfGTj+DFEfG5Q7EN/U65Bmgaz/TDFdr+bO
BLpO5LSqk7xNb/6YCiwBsEktV8FXkMpdxCqPBuS62E60aOmLBIIjeemshsPHvJYs
p44e2Z5jhQpZoOpCzH7qN8qW+UXrQOWiBLfLQ8femHVE/4PS+I680xi5Dy/gTdVJ
ULsEE2IvzRPZxOUle3QV+U+jWrtNKeuG+rZvUsruqTCGRnZqnwRCHueV5YoHc5in
fqf55s9dt2ybOAcvy6jZF5E/w8P1Da+toq0QH2X3PU73cK5KmRZ1pIi1chFDGjFG
aMq5LOeyoXAco4j42LNUMsXtM217svpn4uHtWJXXhQecKHNBgR5W1RhE24VVDXnM
GfxaBeoSLJGSB3tCdIYNAuGYLF6k4Gnioca/jxMyZg0sQ1Ug5KWHJ9ARn8YMIkTU
cjNIROVurW56hypY2lfqwLZvgPPnoFY6U0upTCd+QVZywzIu/BnMz9ch0KnjAV//
MFKKuHOQZ22J+HybQ0GCi3Y6sHmQTIjsN1zjeThOUjFPD4xapbup7vzuWk3GEP7S
rETPPbgfGWtVmfAq3zKnCaCJWLY122bMEuMny5qbq+q3wA/OL0M5g4Bqr0PjxgbC
WEGytNjPE3ZsC4Dk+6zdCdl5CIl/zYsH0YeLyG9ZIzBK648fbtCXDN1IXERUJA8a
Jn40f8Hz7rRb83T/inSVDQVYaUWQ+yWePsQqViYUYEgWcby7BvKa1Puyq24KcVMC
bzSBUoeeYm64HSDW82abbbhzDxFiaGx4bVlXM2ZjC0AoKg2X+dZ1B/f809Nxrkzd
Bfdih7ZzBAia3TW76eMp++sYlDtXSwF4g3rkS2IRjUWMNMICYIR/e/cNsve0l7N9
2fcLjftJTalu2htPPDm91V0BVv3P2EpbCWNQgqv8YN41XSzZquJw71i0SQD/VNpa
j+CF8oEI/o0ZZtTrnh2D1em8qxtOSuLFyE5Ljri7uq8P5waCnYDEZ8uFd7u2Xc/n
McgaThSbApg85kZN67z2RG07J30VFubuHO9x9lJ+DjLtieg+1f6DfaHFzxC1FZAG
/xcu04pBy6q+4f/hUv7lR+rB/urSFQ1o/ZnND0deQeiuqFSkziG1001ATrDwKoMV
M7Tuocypt81VSSohOy9sTxxUxBBnnUYug0enMliHoAH1LQ2aLoUg4jA7vdOXI5jM
4lU023TEmJFtVFMkJ77Tny/aKa64rrt2mJOk2JbKfoufTIp0MKVcSt4P3raXAzjs
dAa+aVOetrEmzi4u5ESlanGkD7JbEz2d5OfnZSexJPrmMFNz/J4MPbfgV9H13OAy
98VuflXfkOIyrlpnFkEbAwdETB9NXa5s4Q3qJQNmY03zTSY6irigG4EXDoBGj4u3
DDcgu6KPhG0mdASn+2Hzu340t6QxF1RA1BNOqb0xXyIPa3kEj+wctSlbMKolzaPw
Yqbt5Nw0lPz/V0ax4fbEuDw8W8djXeSvLHr4CjuJLzx/7+LKT0W+zlLweRZuxqd+
SEq65m2dh+Of3fXNEM1URfRvS4Vif+ZQYgCr51aNI1gTwez1EO9J44GX+hMkzqkC
qbAfjqYBQb+yRo7iZn3/CHEHRX4yTCrnV+X1kp6aCjl6sPuqla0eO25cn/3mGhAR
vs9p+ZhdLtsDVwxlm++ViAJx5AbwZcs5AryongPNt4fTDyHKiDpf22XACSVM84rd
MdksaojdfkUTn8eRyiD3WWG9VB3GJJbLc9odjJGTo4U5wJGnzTNwYKDxRWJoki2e
EFkXNKVw90QkdjMSKoj9nQ3yQxk48M6/JidOt4P79jy++3e1At2aquzY1/6ri9RY
4eHUUDqWa1Lrm1HNHKHxeYWD1UV0lPhjCl7pz3ENq7D4+xfWef4rKGBXEu7ZoslG
VFEb/FndjM1ginFh8wnbm6DrcLHlIFRCTdFwEqP/ejzJQwJK3hZKeT5IJTLU7m4C
Mz6kUhJe1lAGNk4zQIOzAenp0Dtjh3UrSUdoZvCLkRIC+XCfMQyza9xGBxwrQ+dU
AiK8LpQ+uVYx6N1o33TaWaiaxeOtIKBk/znJiErPzmU7F3pJGJ9SNOeT8SIBFuV7
9PW5905eKVaRcCgpYmOjwv5DB6rCeFV1z34mG4bHAhj95pmJfJtHkxSM497xhLEX
R6X+bcAjcdOENwXcxkdxVHhydRwBxxW/i01msmTWrB0u4bCMeeJndLJUol8kT0Jb
pJyGoWdP0pN4gjihZa/l8OePSkcdWCsdc7NrwlyHCG+XVyOFHGwCUxfNDBQutvdT
HBdoChyK6NBvTJ5tQ2yboQi0wLjZFVtS+UNmI+nOCzFHt0PFy9+WQBXlXzoXEnKx
DxeJhn+RCg+t2lCSIMm4hFyfpc+nXqVKkJg0DJcDE+kKFfy3vCJkchsu9Oqn85PD
zR/royvP5I15/A0WJTACA7T6SZrTnSCD3ciYolH4W7iADoLgFzI0xIJy1fBOQRrW
LK47kPa/EgUQ9VYJcznj51OsV0GJ6styidlCVRiv+3os87dVWBSyIn7Xz+q17JmB
KhdsCzEkODlEfPnSlmeVI53IKis3hkfN6Yj0Q06XVLO3yJMpPd6l5tycjph1rCD/
YciUIpUS48S8aAqvjKWpKw5UTg5kv7I9b1fnOQdttxL0TfLGDa+wLSMM4na1sxze
m/7n2T1fznf9H++yZFmPBCyAo1Z0d4bwImLgAhY2jslkfxk92N8N1eI5Q6HYwOkT
sMmQ8TpxZuviFeEI0EOmfXNacHSgv3qC7BJHbEX0Perpp0fe80HncBgxD0oItETW
NrgbTmJXkKGTJgYzfxCuxw8NxL6OabOkkmzojaa1KFPgzIMKXMtWX5Qh0d3XX/Qn
zsNxtE7+ewLF5Osn/KxnMKQaANHeMA2kN0mZgzqEJ7rX741Ze2ZV20TVFreJmt9E
Z7evP4mbsnFs10nhqz3pGei6sGSrK5arNXs/f+W/FGrxaiovJr463CWQRnjxwNiu
yghgGXpE+/UU6q2JlWBNiLdx0ssY85IEvs5pqkPMzKsJGjbdTREyAx17H+LgmdKH
OQ1738h4cT2SVlaY50Y+XCkK4P6JNa/1BKWZkW57KoP53BD38keq/WaNJG2mQV5k
+zZu3Cr460e2+JBMyi6zKR98CZBng/C9LLURRbYVssOVOhA3vj4z44DWtTPT1STJ
6vNj4RkK+rHXTYf5kRhKtguTIrTzKuMNlh6rn9LJkjKuYRGRZMDLP+/HNh4CZbSM
gwt1Okx35ZozTCjQ3gQm94CUXhAte3p/pkYWC/17rdviLZvkj17Gl+8+1E6C/YGa
CM0kKYcTmO+5sarqmCf3HocFDVUEmPZ/3Pd7QEtXnvKIoA9U0gQDPxqiaixcBXgV
fGiV7MATWV0h3Pgi7aDvEoGOjUdaVBDBKQgzExtmT+KHQS4gohVElGjHOdUSdYeh
J5RbvL56QqhexmrZWTscUISYMVHQ7mas+iHLuZxuudIuUnqN1mvN4DdKybuQpGG3
Eg/uZmOuWLfQwCGyV3ThoOUPbaoWXkWOQN4WEBvSeudhXhiStwsA+UZ+m/CqJyk9
PHiUlTXKEKt0BkIiqsUVSb55Dxc6Mhb2RqutWAoBv70CuCFZz038QrUmwCKPfftn
tM/2sjoB94/86mQnfQxQg+uPqm46Wh8Ix3v6NUbKbuMBRx9HoeG+rUavOsVWZMsW
1HxkPKRA1N3yN7TuzC58t2Uzmh/Pn/MhcE6ifnQZD+XyuSxnf4bXDEGe2Ab4JbZB
q9hJpKQAfOu8acVt8Pv8IpKcHLdYOCRquAfrY02GTrSHe9UGrxUmBYkscfvWFUcI
qoIephY2hdzGZJ7OoagWI2nKqBqWLlw+ZWfq9ErZ2cSyfXiBu236IOtumVXTjUnL
SQYUBb3gviEhsMLPRo3zgyPNsDZmcLPFre6p9/gWillGIAzgcshWjATqJxw8QO8N
Vz7LRqFBgKeFqxq2N6FMMjZ8/68JQMSILwNdNNjyF8+96ZjE0HTm1drg7h04HaK3
zEtr+UGYDBaPcgsGLw49Dw7arg3WXApoBnPqjL+FRkgg58SZbKHIJu4MgQzlt++I
+XBihVUnmVWy2t7eeLjys+FTVyQCfpvmYFkV8pQtvkDQ6+JjjV/ITROXPmiWd5sE
bo35zBR4rHy8ZnXAVgL5flb/mmxx/1qeCskhY1fbmQT9yrDlCMmrdkXMoXXnoc4L
c3xWznfpcQPNd504iDC2L2Y2byHAPNky5fvsJNjDY0M+3MVKmT+D3NKWOvdemZI1
NahYGHhubZPzmw6THMV3fjevA2VQcpm7GLyiFzioz94HHZWUtrAdcfdxR+0ZrkrR
xdtd36LBaMbgaRTQ1IfcXUg64j7/IuQQeK36NpWSOgxKvpK2rC59g3tofjNkDajF
/z5BsfQWncXzP4+fozHim7Wg9ahONXNlLm1BhJJrKV4Y3oub8V3KzFY80XsjDwHW
SF09Ykmaxt8ORuYpcvV6RN8KGo/J1Uhx880V30K3tY7Uid6Tsm4yPy6mU5vFCgTI
fCFsRt/afjOHPmGks4ufpYW44UHfGAmZImYiUe6jlJWreSU4IdkEQp6pLARwduGE
gwqWT+0KKqsV14a38r6y+e0C+Me55CEohDxwgS8Gj6Art8S0MDiDP0f9RJkfVVfR
RTdmGI8kf6RW0mhR3J3gvkJBb+o1/bS5GJ/h+mR5QOzxaoJGJ0bTbvEMmn4EV/pE
pdJ1ZiqZ5lSxcAQnR+C6Itom4bOiuIEhY5z7HBBeWBjDcuADxGQkQQtdIQFjQ5ib
I2S4Bn8anpqkgkcDlP9W77dLJ+PLsRU8K7cUslMJpCDy1Ihig2xU6Euy4gdDI0/8
BbTpxgEWY5pR4wNKmkcrkIYBgmm9ShZgh/iSWFwxGOlhXEsFQ33Fy7DQOjSyYlSw
YSC8cKnlyt0dJZvIqBVzaOCSmHbx6P79H0mdXGJGAIyCQ1/Dp/MWVlh4K7pOIwiU
+nWpIQywqBGFelBd6AccQ758RHAaA1+MhazMkU5uCp4AsMjD5n363udL6L2hI+9k
tIJfteYHth6HHcx+kbCIJV/kEPUpM9rOBgMFPGE0VRfyh/uLY1zAV/rVpi94tmEy
csobjFicWhAoaFHOtMBD62vWIbe+KCBeJUTmN1L87vjdvOWCdS/4pnuvbpUqc6r2
QI1Lg2KSL3B9SbdTDH624n5UrgyBczxVLpTKBqQmbQedFQnstmwgQU7LGTzur4PS
37tspcIZkoco6rOX0n5fuuxPEB5F3RSGw3vtZ/gzHbFmgpoY8EYEbZa92z1CiUWV
pEnK+1cYOEbF3xWVO+Bg1sDNc7kmSSrUsOgBMvdGLSebLdD6IrxNsEF/FRALUJnF
ZGHJt1y/If1DJpLs26eTb/LdoOu3GmGEqPiV/+Nho4sVqaYY+flo95WQ3cHk/2LQ
cljavs3UIr0Y9pxkeOKbxAWyTm6/frLd1pktrFwnZpvm+wAkHrNd9XFM+S2DQkL5
ssn9o4QXt4iso3KG4IPZMg3PBqk8y+F4xSAEpU1qQPQ8iHmQZ1WtZhdq0enoFr+T
Uhm1CDbme/YAEJsdr+/7sRKZwtJj3wZBaHh1UUZlu1LZQUBzd20qUGaNiGmd1jQf
DKpozzPnkrm03dEXD6C3ydW74SnDQtmWQqQQzo8P8ULWmsqqSG1ua7aVDddgIYtP
s3yjsbqNDwj8DndjdWdU6+Hzbu2DowfZu8hkuiEwm93HyqSsVX35rxxHvk5GSBJ+
CdoS4HVGT+HbF8yQGoqJ+9nqwZVGetu5mJRtkFUdo88N3iVL7IAN9BVMvcrQ1wV8
UAQwEhRZI/u4fakU3Qga/J+yPwB68h+ogQXyHBYmnRFVbKiPgjYQa87Gr6D8RvWH
cMawFzPdM0uz6xmXVJas1bFrOEGglFGbB4DfARCfiSsyB9VAT1ECruN3v4WTFI0p
KIB5Wu+5xunNbw7Xpq4sulydURExJHNNqTlxIj/EtbDn9wqmLyD690Nag2TrMnOR
ltk/Dub+sO2I59X9MWTNUffww3IBsYwTB2YU2Y9NvDwIx3/wndN9/EuAZ7eoDb70
Ypcrb3zD/DwSqSdat+EVfcH9rOBlt/IKThh2BwGAytQQ+9CYojo/7FewsYU7d7QC
P+/Q4CZeBS7gzrEFxZMml1zxq2Gga5WYezVyWkTGs+QzESUOfPM/PM3iUAlAVErS
JLfqxo0VflL66gseZ/Kc9e7dAZaQJjrD1z3r415ykveL0qONqB93laV3AX/1scoO
hK1doTW+eRMOFLnpaLRojPxq7cm5ROnT2nDo/8xuRdrY7xz/XP6m2+fkRyHWey9f
085h4TC2A+CclAqeNX3TDJFN34aV8n+Afr+ywoEZ60GZcTOiZbju6Mtzm3Y4Im/F
1BYWzGDz+bRD68DV3gVra/nnlQz+fVOeR9DF3bp505FJwppp/NMBwQpKeoWaiDLK
6mVMqceuMjCfeWD760cJ172DPYjLzgV417iW6B0iHGuesaUlqDtHefmHcAF3rHvR
lCEYoi+dcR/EIYDsGjyeB80sxxRNdW9rA3UxH616SGfsWar6BafHkuUr1cM/ntGS
TMOCbt3yPCgLhjhBv/bWTdpwuN/ms3bZwa9cN9kLthjdDT+ADhBg99cTsolG1eVZ
+VW/ldiYkU32Bgef6ImdT/Nr+UN5xJStqWW2O/zXhF2xtRFVDwjJo7b82wVB4r50
LXzei+25JeLGFTMemJEsxsv7J9iIJZNBVAAmaQ88hzvMx4lq6Y86iVwELU+hXZeN
d9CpT8+QZvzw+HSRzWSmQ5wwpjM8+Fv3IBWJKn24N0Ge8W8UpnIdA5ufKck3Q0fz
9pKVNZcRIzphWFhHmx09owJo0c38Lpk5EsQCyCLRVUChHWHJO2oMJqNftlanlCdG
l3kguQVHZTF9ec+rDWY1vEyT2I6me9l4/Hz7H/7payMroeQ+mYWu3UaONLEYbNU3
UbetpHEaD8biOKCBFAde7Gyp4N4jdF6pzZVJSKkZeL3R7y5nDsqmGAJ0eJHPNN0z
TU2WxZIw3balKGDgLz7lTwk1PZrS1FmL9XTV+srV+AuUi6mP7iK/YaHYhybsP4yZ
TMlaCrXS6SzALN2mvr8LaL/wh/tncMoPiebx2qFVXs4tOm7Y5WDW6U337hyqghXA
AyEO5lGCcFWanXe7IdydIKnkmdrVmfahK8GN1+7RH38qX+vMMF3lZAOvyD+Sz8iT
HDS9am26bPmVVC58AL+bUSidR3Tky5nimRLKFKv9vuSOV72UfcdrjvUcY5YCjsNu
VSx47eiwU9Aixxuui2yO621wh/N7nET4vvfJt03fLYXJ/04W+OQGCOpFy8vcvKID
VS9rnLeOHaM9vrMP1vea1w5+zEbK1RzFO4CYzlTcfl/FjRqnsfZf3ZZyjjrMq7hU
CV0C2zt3seOBfm+SFq+818Tlpoxae6LSBP13mZ7D2n3bOeC8HtthMGex8RHB0O8A
rv2fshn/wn73y5bN46DTxB7/JeWLUB+e3tZlboWcBDUBtJOKUmj9K8ITtsadswLc
XR5xyWACjCyopplIo+JfncLVQcSMCkrFgAyfY9xdWjwikokz9GPu0qAugRY76/Dn
2ofxrrBj5pjIWaepHNBKSCBxmbwqJ3F8IPeMZXP8/PBXVjUoTwsIe8Qhh5cFI5+6
Auf5OGEhuu8q1cac4+0+r3ZrH0e1jF65LQb3u+//7FljQQSWYUcBTzdM6DWbgvZ7
ZzDaDEEYPL5M4YC3ceqjnEdM0aSfJ7an2rgsEMQhJBWek2Z4YKD8GvaZ2Zsq8Q/T
1bBk4Hs/CnWlJSOU4El03MPBRmjKcaLN2Ej9ASMCbmNoZzacRBh8+QV03sE0HahP
ikLEgUI8xOvW6ULqp4tX8Uj5rh0FpSo622/bVYFNs1i7z6OFEjEdXhuPqRl0dxY1
qxeLOVJjCeaXekxOcIPPcwWpZc9tZDohQ7fSiL0q4nyAP59zdaQFj3nH7kNB1zQe
bDbCoK1z2juX3eMtE/SFOBMSIjDWNKtTcWpu54/nlY31gG0IgHLmRmmlWvPY31Uy
gIWoU/8cWGuAigs3ka3hQOljEtSpwg2CNeqmJfMwMdUhy49O1Jo53mgdx/FwwVjI
znSIw9aLK5cHbh8cuAksPqcdwb96EJTVp7Z10ldexGWRiGB0wMMugtg+j1b4ZkAB
bEVZY8iUtD/PCfvltGv1SKZOx23t0Tq/VaUimNulX56G5XqecmrzIp7j2hHVnlOY
k7X5DERNJEAzR8dvt5IOgzx6jbK2dnhED+mS7zTj72Yj5UdIBnUynLxvGLHkBkR8
YL4bjmUJHmMkvlEvL/vjgutPbFLXvgxT7fhoQPmDfY45grG0KAkq5/0FcZ4Qb1DV
waaBr62wM7rOauCOGP+0QQc/8gwdPTVz76L7n1DgAkQLEE9HvbxF8n23mHG/vHuF
lKk8ISA9vS9id40lthkDu0Maqno55rybRW33/+jHz6/LcST2f16Fs42svwiR/Bip
JEWwHyHOU8yJJxwaicm+/AR+96HDK7NO3NpQidv4zVJU6olerudxb3+/I0i1Gi19
g9Wwdzfz31xqYxZGYZj9TAfTztP8K3Ya3xNYf+Nyz85LbRIodJsLdyIDfsZxYYNU
ujPq/HLaFGw1sGud+fXlpgl+d/NoyjdxXJjXD6We/FNRrR5RhB5wAFBZAjqwTbsc
ICzlhJIJKwruf0eqFbfjlscZkKJUYVGP5NDkMgsvm4+9v+B+jLhfFPe6LwQg3JWo
APpu+loeGByQZRVesARHpi/p9UvSjaQ3F93Z91UwVEc1AFeeYhSR6ZNOGSH6Zdoj
ZISy0h4pfv14FwwvpdisvWlOzFwwaPKWfixHAdfeKGUrCl87R4qd0qJBKqqwCDh4
g97kguFxAi9OS23KhDEV0Wa8rhI331DC+Kn+NdwxGW3YwZhg3/TqPTil9j8/UIvh
1TDNi6PGjGWGWKy+Az2/9FIZj3UdnyDXy+5EBa7DtnPHCiHRb0uLD/NqfjYvyH9o
apyI4WIfdbiFQcY9uk7aO8sSDBHGjCzIyvluBxXDhHDAV64HGQNIYVOs4Pn1Kv7/
3aQ7qmeTNW8eL+vhfwlbUTFjGJ1JUJzpMdJZbqvYveRehGF+QyvFpU9IC9zxPlEE
t7CvUA8ZCZdcuWki3w/psUu+chWS37O+WVs/48uiiZpw1WLgkVbjIxbv9SdAXwp4
I7PZK7e2FmdUaLoUxsoyxAdCMincK1Y+Wrqj/QUlmV9o3WH9buCE/FTAV/I11tC4
vvWgOJR72qWXiLqGTYF+0C4QHsNpQrkRwDeX19O4zkCno6QzZ2K1sUl6Hx3UpJlj
Qk04jpB9u8VXVLMgNCk0V3KRWPVMsW+SZu+ic9zpDLXTeAynN3Xh4JbrcjLoCOIs
UUzK/nyTPcLjSb8/4HKfIX5v7yVSZ1haudhvZE/QclJ6y4vm3pi9ixmL8gpzu63j
xkoJT4geAZnO+3mD0iee6lRVeCb4AlT+gTUieRn8hIziI4Gw9hRsjv22IdXG7I0G
Nj1/b7a1Na3+DKHwCEWW93vbLX4NU9i4AGYjXSzRNxIBRhl+Cw5PKMXFwS7Druih
KJAgfLHTX9fSxgdjTtnDXWvi+WVtlZHiSc1oqSLMWtCSsByW7FicXhnqA8CT8DpJ
Zy0bepiOIHTUdBIWKQajaK5zMHtgNmSJ3gBXfLAvpDkUFt25wOwuhMwosHm1oW1S
/o2za4UGr7tZBeGzznFslDOpP0j7c+p7A+gthJWM2+OT++NFiYnyAAjt9tEYkUre
O7JpeCYygIZAZjDDLmSdTwpD1arSU8VRYbmk1ILi3g/Hp7CN8CsApTcGBkNX/d51
Z21dalVX37vSLWfQiL//MJPS4YREhpFAK1hkCnDTF13OMh7/9jnmA9fNxjQmwVyG
wqSLQM72euOYS8l7Jh0MmmIqw2WvWDq8MS9EFu9CypFRH3T61V5r+RvIdyXwUZ/p
IV6XJZ4bV5H51DeCGhTWLe0ILNwwOVGGMQfr9PqEOgHoX9E/ZVBlKoSEa+HkPGb9
SzqXNJXm9PUJp0uOes4xkn6goqMCzIFN9x/m54MJoiiHGdZ9jFU0LstpLOPnclqc
PRk8xrosDkVwDUXzha0hGddtfwRcwqOnae5MZHz/V63nP/vBd/QkQxn1qzrjDq2O
0spt4sQ3mdOCy2CrGlsfUax5JE3ETruavVKzA/a5gT42FhZoXYkvDxo8SDpyviqq
QPabs6mLJhb98wykJXEUPiH9v72HSEVvaXBUkb2Bm6HEKFhxDe6HTmXB/abbjfPY
wq2qz+GSaWePgmuGa3CuTWABqq9g7DaVmVPyeiQkNvlVg78uG1BdMWjwNdrtilbO
0XzFFCbvbho/vUOe/Opj1fgC9fwVZdxyQXVoQSRdc8EHB3TSEvNc2aknRBBuE6dj
kgShEKuyzmgSRkpF9XPoaNXYRpALFVoEkUzWqRbE3WcALm/RToSi2uxGiY+PxkxT
7f6WuVFYUNssj9bQrOPIVmgjWpYiokNvLHLGNtZ0LbKbZ41UQqhASjCnzFZVYcEs
K87myCKFZZoZbn4iEzE6DofW1FUe/nSGZbMIyOm7JaQahErttSDZfhUHpVtpzRCS
5oHsCI/6eCS0nMCpdYXheIoIltBIRIp/bUoY0R6oNyglAc+C3aewNEkYlvY9Uj5t
HiscSp2/aR2zYzs3807Vq/UK1aYza0wYfVWiU9l0Djro4ZFWW4s1Br6+AH+zcykg
qlfjVVetnaEnlThm2JMT0NvyEBPQ2PncVxz15iGVlUEFvYYdl2Lb0eup0L+etyHp
gtjthfYPtwL+UuaUwrxFkXci7uuX5XYruUGpZlEM32u7opatDpkLzKsoWUYqj+Z6
jlSivY5qWHT9EAT3LPT7CNAEjA72T5alyZR6lKT6XVnGs2KGTrUiQe7tIhXtFyjk
/03HS20IvlHYNhR6vlRaaekGhc6Zd/lceceA31EGPriiz6+H3VEnvW1sqMmGom2w
S7DXp9aOnbT9XLGHpNxOYEgUEB2YFBnoXPszNSFxq4ZxLwXxHe5MvPGna+v6FM2b
bXqOWOsp385V9l6Bc9qnHOamTIOUao8WypmiRE+sL5UyffFPY0VxfDALC/xeuT0e
TL6C/4qg0BbfRbtf909cvYm0Brih7blj2+rstaBN1In2VyIz7LfT8dPU1jKV6Mdw
g1BPwg30noit25yqafiY1EwxEBD60DWiqH1JrU49uPTMepmRPtQXEOF0JECGhsLL
6J1GKZDQpsynMzMIEaxiL36XmqQd+W9sFO7w7reQky0cYmBAsRugqKf9XKTkIea2
uB+jgKdiau2p+82QTpR0tTcn17m4o31LapbiLxxYro7qpTXm77mFjFBMhUarGZdj
sUab95WY8SDwLJXO7Uoa9//BXz+3qdiZHEf55vLnA6jpX0e76yNt1PIbKER5HZK1
KrI7XlO9SxJ+qUx8G7pBL0z2P6KCA2dukDJQeTjbjopqcPxXPeRw1tWjOinFCnRq
+jG87GwIZOqNa1sUNJIVR7qTaBo5/8VSxHa71A/NHoRcJ3rKbHYMG8n+nACqU7CY
czFB6TFe0lTCFhwV3vz2AJvAMiEiA4S9WnfvFvc4w2BgZh1xw+i0tvRJY/TJ4v/j
UXGaoxWYpq0yZyXCAalMhpN3LIMs+/mEq/dMOizDjOmo8eXtGxUq2x2BtOc1/keG
Y9uhMLy5OyJyfasiI1T4fi65BbjFXhq9Ad86V74NSAjRazawJYD8XMq4r+sevb9c
NNJ768vZYNGiAVhjOogjciV9BTFDHNK60dyZ8EhfV4YHvkXEy266dtFf5nPnDU3u
3CCX86KRKUFA4REPkp7iv83llXYJqCNd5tP60bAdwyRA9BzbXRiINRQUvQPNw6KD
8S5bTmxI+gwf5XE9nzHX+XkirShjsJ0Y2bQbVoTBGleM9IJsIFKvAUAcWJE0iFFg
XzphfLmCPfQim2iEXlTEgpVWm/xIguCJRX2sI9oOkioB99B/dsIQq1KiCMJSaapn
bLJftzq60FDkkkTQeP2u5r0abv+vZr5WzQ4PyjsbELGmp3Cp4y8hXsoLW/JsH9T0
7xvDPDQmN0TBu5nGO7r4iR4dnOQBXDF0u7bxQmxROxQxLZ94Jyk+q9DE8okG0ABT
NK9TF4Nb/Hscvrk4Htbxvz999IqsWa3CHLNkR3za5s0Y1ikKH6YUfPV291sSdp7X
JKakeVXfvoRH2d84UG4yXCQbKdTEJZuap+HEAEHCQHiwjylCeoM7+R9ubpKIJ+Um
/6kxc4N37BoDVYOW+l3FjY1Q2Ygf03AS81drmu5dqypOHeeX+OpZNvTdOBc9q4Y8
XhNJ4imZ7wZyTeI74PcF+CGWtPGNqfiM1dq2Tmx5Sf8xhz9r5SAEzx70bdInvYIE
KSV4Dzi5aqdtX47eXMwQscnpXTWLaXPegJouMIfoFl3lt9m1Wy8ATq/3VRSRhFX4
6+PMup9H8MG33dCV8YavH/B8ove3T0bOEgQt8r4Xr4mwl7UI//QEHIaX5Y8Nxcky
dn3N4dZVTVQUyZ8Teodnq/rXiXOakh51DvXr5xl5MOkSnVFMXXqFLM886f9qLdHn
0IPnM7+1hpcfFK55mvMEL9yjM0D7rAiu1SzU2X7+sF8fI5rw8YPDW0cYl3UzfyhS
hfX4b+TE2c6xanruP8APpl/DFmDgbKuxh2RCpfbCot1xaxUhvS2rSk9b5Q085Mjc
tIRaKuI+qLXmjhmHXmYXJ9UlksXsnlS0Fyy2yIHIhhTouQ80VWyQC5qoG737x7dH
v2UXqFHaWF+7ockYyFGWw5oQd73sWtGxK5/vzuyt59HozboRUhKvhWol7SI8RqVg
IYmWlGPyHGIGluEEnPg9ALLSw4J1LZa5PYxTm/rYysJapojJ50TJwKKLiAHuPBBv
7yhAdVft0lYf79i4EllAHee3v6fmsSq5qZtYrwQxO2A3jQ3n6WMAsq2ukSPjYZTN
fPZ0X4q6qEMhLe3WqEBzUhJ/23XEM/a9fD18d2NlgMaAXBTlxApZGfpSp00PSbDs
9kpDK5Uo88g3DIq6Ew6tJGGVDYkiFdlKvgdL2F0XpCnAGqoH2DvTfSeVCc85Vb+E
JDCKKOEgfy01DcDhowishTOXcEA6EM1iS6hIFsl8lCMlSwq+CHP9Vw7J2KIkzXU/
SxkkEef5eMVAUSMon4haMh0UCk09KrYoYZD5zISRw37HJYzRbJ/HRmeg6BAWisE1
+oA16WhXgnWCY1b0HreOKKBHxhNNgtmXfA+6DEBBPg0n8+gFTMPLtlhILJeT2fKJ
aVBj5vjuqxA3iHC+knyV/HQOKkAIuPCScnLxAdZGMsf2j6pSyp3zVYpr1UzkTbp6
R4O0YVNJocKxLVFarj04WH66ax8Qvveq+Dgwwy2HIvd+GTZOUyvExKPXDoA2MM+B
Z2vYsU6WQKix2mTXgGwxh6OOMAbwKxtS+zMWSwrJCTCotC+aIyZDYr5rhnzUP0rE
g0gQlZq2Z1ngweMwIOpt6IOlI2Tik3Se+6JkCOMKibehSOqcFxBBRzObkoYlQtwL
Sdys4IvmuhEbmJCBaXkfXNVMDY8I34+zdwDsLY2CY/k6Hx8zHU6mKWCFy8UrgOzi
Y9xJumL5k03jg1GRATVw0ZlKmMMk7NVcGibVyCkgsT42UZshZd9ss/o5SPuP90ux
AY2CHbu8yJMt8xaRajljZCeHbZvhUPHzUbPBrECw3x/jAnxh5vzWtbm6cIytZJu1
ZDLWagSRDPTNZKE4rS9txnnuJtahoub5jOxmYfSpubktKMrcAsUsINJroWN57Wy/
yeLE1tNcAqAvOpKMRz0mhLmZiVnY76cZGh88bMLdMZRtQGwBCqkNHJh1kEI9ixlv
eNvUw031KpF9yskVfy3Gtz/8+4XX9IFVhcNRw+uulgq8DSqQ+XrWFU8Jpd0x+1cy
LGNfW2u5nB3lUBMhqYXfAPrdi3M1G66303UFHmv6JFcBNYwTAs99yMXmvKNwAG8y
Ve8qv3PjFW55r21VZnEylbHMdLVBx4+wlJJBx8R6dTbXjNEFvakJaDDXEw7DXiSl
ds8jvCDjCx4No0t3/FadrLZKHfrY0repoOC32U1NSX4Z5ppWj1n9mIxmZ+N9+J6w
975Fv7YOjHr3mQXORolSpGofKv8/Q2+iYZhNoKrq3baUZwQeGmR1VRmlhqGLDtcq
5omANM7UPrpyT0rKXP2rNlfDSb+53047kLI1pPKa24CzqxmyBcSdteESwW+1fOuG
hiN9BRz/mYDbwJpXmx1Ova1QT/kkq36Dy2tgXoshhaCJuC8ZomKOW153HOG/TyUs
N6EH3xCfiJihaH+sIme3GrBi3jOuLDBW3bbSkilS2EA1elq0sC758qdPIDLXA4r9
RBkwus3atloQzohSMR/LLd4H4VOrGGOeJaHKLcW7lUTyunWMWb+aih3b7X3j1int
F6gOswIHwkRsHr4aDAWGZm1H3GDs+JqSyrZhdb6/zAKFJVEtaL5D4picGkbwWm3z
VhDuNiH6k830uUxyCSgjOvsacFogusmNry0LF9yRZAQ0C7Vh0yBt+RlV2u8TMIxl
koo8G5j//LvlXVplqnA4iwmvVG7vxxkvCUIkzjm7ou3CvUIPoeZlUiIJzaMqvB6Q
Cs3UoQceIAmNON51rf0ejB7gIw31C604Bquw64eEshcZMO/qQuFs5YRSGK5xGcQr
wSZoNsLWSRVaBpTV3kaPDVNH7kjm8zEX7FQnWm4s4QqqrOVtmfDFECqU9Ci5wGXz
BsrEE/NrkFbhJcacVnKE3/wBFUcucZY2UB9SjGHsANOJ5PAKv5uW+qJB5tTMz6m6
SfBmyvYYRyoCfJ8RuNPvqaiv+UfyesH2IEkUFL6E2KHAteUNtAgfUfpfts7O1z56
STuxyaYICglpARzW1Wg2QUtFn/7rPPoIaXdCiXcE48LvsnPt3eYoK4bmpaaO3Din
5HKMJS6kKffhE28o8XSPNMpEorIWeAP1FZ4fEwX3D15HU+o+JGsOooIfCmYgudJQ
gEE3U4i7bA5cD/3WBouur5rtufFdh306ezO0736gqqmgn6wUopJNm2yr+Q0AQJju
JGVdialN+8AOeXjoKvrbZ8STp7DK/qf7l//1xTK4NaZUPjGvZYKWVNWaOhCz1/Vy
RnJo+jrZ24sq2wVHooA5kn1g+oQMr8GtOrUl3/D6VK2yJfAFqBpjSR9D6FIMWcWG
9mF7R/cfYmRPut4ra3dLaesPqRdWgF9V+s6eElzeSYj1y3us5LbKpdjOsZjvcTUC
dmktkV6uLauXU6qcQ96yT+MpabhH+yCYiilq4aMsYlAykfC9MUq8KzZNTdYYPyCP
6UjNSBIZeGM5quHIdUNmcuFVBXwffm+eAUD7qpp+6SKBZ+N/g+t8jeLrQkcrvRv/
XQPwzDjcthzdBk9NujyNTHNCNjYm3/HwNVgeaUxlcnj2TIkEH2Quh4sjGItFYZdx
0dtEWiNklE4ch74iqkKKykzUYRm4gwtZfPwrkrO6zKXjUH93C13ZeKROwy1WlP9z
yoELlFAzbpYUfNuDBFnRQgSkXn3LCXoEfhxppMRuvFiIWGRnwuhhW+EygcPJsdp9
Ml+C1n0Dt5wnrLT6CsYAx7rX/VFqINAYBgJBAT+ifY60EQfGkDfxXNDJWLd3vpb5
ebk5x+WO02LhwI6VC/dziNCLW5+Zt4P1LotT9/ic48QX1wliVMl7sOIgiqd1SMku
rCOQvzqweZPmUnBBT25WZJeEoIlW9F/VhNMijjrTDQihCGWh9zQCG8CUqo6sWe3h
nu1Nu3+HPxHHTVMHKXS41hbcPvsOcKCOsWLiJhFG/5rJdlX54mljrmwz+pelhIz7
YR2/jprkVhHTkzlpgyNlkuk/S1gGKEzr1OagX18gibGca4ioDbFfX/z2EHBi5P1P
5u/75kvidHwYtg0rQf8j/Qn9rT2rqDmtOyEoWooR7zfvi4KQepGRQrhtqLwxCT2B
ShQ8SIGTVzHc3swWyhyUGaIJu+T7bSDEr8fQot+1AVNDxkE4otsM3gIajYplaOO8
66bkWmPJ2v0f+63Ik/LoVxOw5DGEPr6zDArvKFQ78Cglb3rdtXvPuphzWPVV1VT5
efXYEPQxWPGtBuwoabzBNPHx+XLgFoVhJLaaFM47pslW/h+bZuawtKfmhZwVSESY
EA4SRb1wMrkVTcdOQb6R/Ry8wb9EK2JRXahaF+rhKOpf0xumWV0JWoHp5Bmrw1fR
VtoqT3fxTJ2030hT/EMh6gOwpuDA6Ll2lwcPZTk2HnvSGZnTh9tc56DJxUPhq1O7
BlA68xkfKpbjCTaLIS6uSAKLA+oVZ6XAjN29f7fdARJ0YYIxTENfM4RbVyykygJ/
gE4N0KrESHKNpT6mJawsYfBihs0kjKCZ33Vzcpr7MjH/YOlfw6OOg6/qSfLluySa
Bqw7FKYYsrFsV3rA8o+hZk+OcKkqnvVzXR78RVI0MyQxLCM5jzo5VCA3y7mkKeC4
YcZciCviFmGGnrgE5suX9J3C02nDyo7oZnEsNFdooOYbvJi1N9y5Gkw7lwDG0kW9
wZPw0vfmOsYvNfE311ZtC+pzlENEvs+DwPqvfRjQlFHNfjngt1E6bp+HMg4OT/ug
/wFXUehbZ44hswqrUNZTa7PNfaLVltAfvdN78wfoDNzxhJ4/+cs0IS5VpIDwel5p
Hh+g3UxbdE6Da2BoB29f9dlbhxoIvzEFi+60+paI+7QfAfbZGiknf5zrN4bd9V/r
UsMdh4xCLd9/jayX9+4zfG9No+bH0gjsMtyrIi7c6AgJ+g9uc6GJiI0XCXYh/WsC
6Uy459NhkdKTTRWdqoVRd46qtw8OrHkPhrlhC+16i0f4aKgp0IZDF7b6hExCBbLf
GZcAoWTA6ZLBG/vfq16G8q1d6Y1EMkYYxP4/j93Dho6lzAHLmPczvOt9iZ5FGCzD
IFNyFv7aZtTZi4lfonEM+j+3/W13Nom7mDLKbBcfTS4oAIP3raI3ShrX/eQlHF/Q
ykHauuvIxoOsiqJA0B+CnaTuo1h2Kny+LM1XqrZM1Dp2EKshdKQ7rtHdbgONZDZr
QaH+B5Gd7BLK2o057bVdjJoih2vv3Lo2wpisz7N1qAJbjpXxVDd6QUVeH6y6E/Ro
MxkL5muIvizxO/x9WBNzX9TeD+fESKam04sUA3Pr21U6ToQ9VNwXiPUU5kuNfIhx
d7gfAv+MBBB3obNYbrZPUBeTUTEs8/6p75jvohoWDFu0Hp2h178FNY52+u06Lb1C
5u+h3nfsjZIzONHkyzPih7OjLiodKMl8QjRKisR5T1if+XwLqaJEi1tGCX9EqUzc
9AhVQ2rdDZtj6sry7bwg4U0NtiJWIoeqpO6Heo6zXwMcvyo46gL+N9qsx7op68DH
+wWTE178QBMZS55sPfWuZTDAFvpA3ihQ8Jsf9gDiEQ9I60XCN9JaO5vJKcwAmVVO
RIVONso2kKoLgAM+p8zd2QClfQYGvzGBZyLKuReQCQ7sr13SgloLqkruuJ3fLFlN
W4FDzBFVYZxF4hGZRe/+4b6H1Cqnuad0tbt0sOeNDM3KzQ4AhJHiB91t4fJr8pE5
pK7pGZXz6HV18fEXTz1/712j8BOzoNWdBzwJJsosAPUBmLFtZ8vgbnsE4YA6nWgL
WRvGUjUvlJIjY/S5xebxH561nSJPEWWi9JJxgxnd9+zZRw8qE9YSjo4iHwnZh9in
FPLbDfFQDQR28wDiGRH44AC9kAUOiSbCf6BZ3vUMVxcAX0vW6gUoMkM7tgeuJ9wS
2cn3UQJISmDXlc2qNFF39NMIO8mtPNtpavym1DMiVJt4KGrDau5YAIv+Y+RQHsYY
wWCwgi3UlUKvCdHlnOJaBzHPRyL3fsIY2GxeY3yn/oD9hkme8m7yz1l1Qdkk2INe
n2bAWX5W+8Ux+Hy8b/esgQWYnhLR9Q2N3LazTkAaDHfPulZoiuTn2dn/P0OhqRMv
RbV6ZbSVx57dKJnn+G7+XGzvw/B0yOjVtDmnTXluuSH6O1Q0xmFk0lr/XZHzUofF
lBGoh7UCnnW8MdyP+9HGkxkIj6iMbcScyBd8rdtGSKAYuNDXCfZuIHJuUry6W1Bb
nLockI8dHv8e/7tXK4iRJedYzBxnTnnI4YuNzzRhSgLEWOI6+clKA2yc1By6EZW1
XX7qWydR7UJf2Pp2kLF5ugq9aX6Z0v53uOc2PsMS3Uy1uD0CTbXeR5e4R34PvfLL
lFXHvwysWVgfhK3qqY41zD5DaazLnyhu2/ZnAqkxwSJZO9sZZRXxJbCFz4eYxAYu
wLFtyqk7Ug0AJRz+z3i0Gx3mtcxzVydTOmhpy6U3Y1ZFYWwxv3AVteNeSV7PfcQc
l8rxZysUkfzdH+fM7DHUvBLRKFQcIr4Hzl+xJrUGnHfpaIVUoUmM1MoEAc0stcE0
yL6a/tzbT7MfetFCbsenMpsREsc4mezNl0X0XXNYdOAfR+0Wm28FkPyGJY+6FRYp
G2mx+1Xl+hZoMm9sZAmuxVj4UTa+2Uat/VzRm8qqiKlY7+T2ngPTlm9/6L0t2gms
0OBdfBSgHClbzmJ/bFJkYV7EIArWltDF+TqLAk4l/Zx7VBr5gDkgkBd/fLVEQYjp
wqbhbZEQRdEXkw2SKpBoyEZvZBBBXUgWB0wEYwhZxcdNHjAVmjUvuTXcT/ilrjwL
OtNO//hPR1GfGzC+F5GH8BCj7FVinYdU7dAcZr0U8ct3Y0bScuUfOkI+E9tLkP2n
mW5UMmMNiYPy10HBNiQs01ZWU8RsoJ3gvDTf5gRyOYFqbyVB3mbF0drTLqWGH5uG
zEnnayY3PAGmxLsTGU4ozefKDNScalbsHCSysMl3woSC8t9/zPF0r18MTjX84ehQ
pXSkhm6YVLzTsgZ4tKLMOrkBiwslOfItmFsMiqa1Gc+LdkUDmqAHLEc1waKGcwNg
zNq5rhdAeGSPrn66D4RVSt/49hwx/yUQ9PZtqC5OW5nDpg0DJyrzR5YZZP38JC+N
3eMoVAzhs/Klg4Lo98FP3FVufHHzYF4aJ3M4EED43Epw3imVpSU513830Mr/BzkJ
Q+GPLHdZgTYSJABrgmhn3SbuHBBfynf++cu+tYV0n080frIUtO1CcVB1KdYXyQHU
jnQ5RdEiID2pzo2ex+zc7jlfGtm9jUhblzjLATPO8lWRcP1AXKwUJi5IiDkmwWh2
iHnti1o+Y+DqLEGevsjkgvfMcIeoEglYqfccTigO2E/DXtPzFZ7HVhArvI37xTQL
25+ttWQ+pahTdoOjoUdqA3YEUM7sGr2le0Gk6Q5LO2CvThcaJ99/bEex4/sv/fuu
JFVbEeRd30q0S8W1VkGX02ih6+a10Sl3WlPyDalsncuBWi43p1uAMzImCbyWclmD
689v6BkvYySRLpEku77juoWcaAq5olrnBxWOdADrEA9UyHikHFhjmOxN0gQzN3Kn
e6t6m5tSscrg6FmnAGkzoA1LwtieEmOMMUinVB2/n47h/UMqS0XwFoC/ZfLlVi4s
jWLAK3OzLEubKQrnjiidMFtIB9kj2lwYNf5NpU6D6fFhaTnzpN9hs8mWo2uQAj/h
y2+PjTGn6Mu+VGzRwV+9K239YwLkUyZ1L2UPKi7tIOSA7AGRJqrMqNUVOPVcfmeh
bpQtFQezM05B5jvUYd6zzYu3vYZ67oL92DUgzEkkklFMRPwlhijNfP3KoYOtLi5n
71rC8mVzL+lMmkxQCTm6gCigGh6FxMEBff8Zm4QqGk49ErEEHg9RFH6Tmzgh2yGl
0n2wnaewxqxg2Ej7jil09DamklnGTIBfUcakFkDJJu115PZxnTR01IsXbySZZUoI
2hV093TbS7KUYZtNs7G8iKeFsRxIQ+FKrSwDrJzY80FMVENOG7Q4mchDAEJsu7GS
XAvTCR4tuK3OVIIPsQ3cz47lIosl/ziiO5vUHXKeoUJb2A/YtUfJXgW/TrdIw8v1
YUY7G6DrGtQqiwNqOoZSdcrnd6FDacqUzyVaHZBoedJd0EDfy9Yk9zJVrRf05rRU
yRprjVlRAmUj1lhVM7XB9wfPbX7I4saRZ3eN6Ln4HNLoVeAG7jBD3ukNgKlNjNLi
TXpcrO4kyC7R6DXVGRI51NehvYBnJ+gpjYvoWLvk3XBCPahT2GKqoj+NmWhHOYph
z3KinDz7hyNa10hu1m5qInqqr1kB8C77tGF39nIEUegZuYDS2VsF8zf94ZvDU4mg
7fywk+S/nvDnuZvXSBknwhErdzognk4PwQnXChU9d1mWqx5KZPkX1SJO1OPimz06
XgVZ61k716VweaurATol7lVTs9VTl2L6KV6MJK0hA7gJQaJmDWuwiySJarOm9lm5
Ua6/PB0NPKWCkoX1m+9f9ehYjrAouWLVH997cSo44H0qJ6qaLLQG8J6+MiebW8cP
k+BEkBic6wfUW1YrLtg3Sf4s4mqArXnwX7YvomMRwOKePjKVxVp/Ac35JKiHgbpA
gT1XDPkQiM9RhBOyW0yhf7IV4oe8cEymMllW1aKqACOxf8SDeh6VBnmOFg249yqo
IMHGYPkGuT1v9zvYnkK3ce800vzhXsxNWo4FTVb9grOJtdcm3Q93QDT2vPz3VZEP
SOTvnMMqhMuzcIzRrDT14lcZiSscjgprqRM2sMxHynT1D5lBqLdM/ujAzzVjJ3aK
Seuedp4rTFsBF7OIO0sB0SYwcQtLyNE2q0RwKQOAma7OlVwVr8HYrakFKgoUk4eX
XpacKR7/cYwGdnh4jnWXmx2CO2mORSTAJqNMzjrWCojIXaRy4r0gs0xed1FhyZeO
4suZTDxA8IMjxByXyG9WdBcWXxQZyBY5hhJN1oW1rbCybMIMZkMXHzY0VmZBpoza
2l7SphVmVzIfTecIDbxHEXc5HRY4TKdJaw/X4YffGljaIUTYrRdr4avFUCgH5Hpg
RdblFAsBHRGvJaQCMgdpEqVuvOPNNes1XFB00T9p6QTYShusfK/HLVceFAGc4Nlr
qRtijUuLqUUUomsEz3q9Doc7ZAZGNiw2pSXZxiNxlWBbKW7nQpwMM2AMZzEGwUdK
V5EnAgU4Awj8deUjg9OBbtmTxp8F/2/G+64LMbuiNU+qtiU5OQA7c7uCUHKljNKO
SLqo0DVTlWx9blDpk1PXQSTE40EQdHgC+6cOzHNq0R1z2xJwmOI6cleMcjZ6W+Sf
mluV7qBR2YOnrQFI49D1wK0HT/crkQR/I9nn6du1kOqkhJUdsS5nom7HwBss8RAC
ERJvAf2FWd4iZetn6XXGtqsm1BPdWVL85Wh0f55T9gqRPdUd5/GlALHvlB6TVA5S
X9Wf+PdjlFcUgJag7+wXVQpcxBq/d1CwzuHPBbyuVO6d2qaNkWe4gSkff+/KT8Ug
D3CHB/8wQvt/aS83cRK5ba+Gd4RgxBGv0DUugHydRAv/DjpUYWvBv4YX7KnxslaS
mwdWujrQyhqTqJanoPkrYXWfjEdoNCPM4EVtF1FCeu11TsCo2T7ujhszMxLNS8c0
J4LIAuyQMtC6m7QUmpE9mBNSzDvEcgHK2r+re3D3rzOuhU61OUGvYj5LKc23bMoA
gzP0Ku87y6JeajLNlH6hmjNzspez27bf2Bb+O3g5V5wXWu10Nqpphb1NXPsoivsp
dsIhgGmc1R+knpv+xbtshWEq3wNpZrEDkItnz4Og6TAs2OHO1JDFPgfbweY9XHDl
7UCbEpxY2VkfALJsNRdss92b99Z91nJPqhmXrMLpaaVDgFxwn74q3s5dUScGUAMm
aHysfEhjq6E649AScTmwKV1BrEQqIuvrcuk7oJ4x/VCZzOPrdUuMKsxlleC/6xg6
3AnMVKk51GJQDtKrJr7fim/7KCJHZ10QmRdJHJKL8DBoT2HN9gp4S0A0gdd4xiin
KASniPS3abkbzQuXbgCBgOcSlfckU0w9ciK1p9NjFSqEtyKaIumYWdowHLLpw3b1
UlzBZeU+GLs+g7MqTgvmGhJ7gSSt3Vy9gJC5KZedTi/iv8g24ZVghhlsBept0iIX
n+rOPxpdTs25REkuVwq5cTF+5PioHzrzL1Lkao2h8rYiz3WWiTI+yB0pOgwqioN/
P2nNMOKfHZz/1vMRKbOLUM+e08N/zYwr3ueKUkdDjiCUbtBwb3NTDL6dk7+9n74x
fqSZ22D3uh4aukGOACydqxECCMOon09xlTfAm/YQ0oIoz5lZZ3wOW7Em/t7+fw3h
1SiVvpee8w9GFuDBsD41JCriqQ8XH6UbOOh+WT0yEyglvdNUTXVA6dMNWM+3RW88
IZHP8y01gQCj5LLVaG0nQoZZ48Ifohf4VAzpNsdkQA/QG0riXjDWq1Fv3ttCFgWw
zP+F5PpXvbSk7/GYBOiTIA2BORkznio9Sq4m6c4G1jv2ZkrHBczPRpzG9fD0dwDG
FVk+5fqtZVH3B/pLAGwBF5GdJgyWHi/uru2ZrE+mHcYqUADZ4aceL249nslKz1AF
N3butniFIR7fVqr6JITsh9gRGiRGi/gC0WG7xj9Nr4Z7WNa5vI1yzmRexDDmqeTi
Tza+BHP5b/eBcDobYxgMsEMK5Cw0ohpXVMC21nY2H+JUmiRe9nSNz4cuo4qDwKMh
QE7xkA/qdGT0CxxvDhGZgyBDnmf1tbI9/DNIQbqQbCiufN6APEiG/7oXouVseAn+
z7qnVqz615ejfw80SfR3BuNYvseR2s9FVk8w8Se1bk64FIZoZRLMEeY79jc87ZXo
9Bkz0LIoWSmu7SiPHeP4cwRGPYE+4SQg2EFdt13+9fub5LnRYQFjlQSwC4ZKdpnD
XnkiQ9nwnarVzOZUIuRtZqNXS8XHl0s4O81j3PWY1b+AXGSjx13IK546I0GRYCH7
QYeTGnqrbD31AgGzdKYi4yRLTqU1iK+fo5TO/Gxhtf4RcYGP6GawYmSyyf/c2PTL
r3MROX94MhHsDp+m8fbdFly5qQeWKDr4XOc6KXxgpFvjqE48pmiDdh2hG8MZYBOx
w/fAGx9344vOlaHDNA3rY20vYhkPq6Mb/3a/TpFaxU9xnem0LrZrPcTwA9UlrjYc
fhLbYJA8dlUfd+SQiyPvgfmNOlq6sVM/Mud/wO8Hbh8dwGpdwk5Mpkg0w7o13BEK
6jA4GGGGh207VrsyisWlZaOlApIj3dcI2BW7v1xUZu3PkX5YpUFIu8DaI2OpXAen
SNwxuuqcZqzKPNWQIOco05L19cA7b0q2HPNG4M+XNzXRQPAGEAEtQTE3lGBoAtGR
+RbpAOJtm/uzeNNzKo7p56q+BgksDg1uJjvsP2/riW1U1+mQ0Y/hEJTEbLjXr6n3
NHVtNdx8FFvxDxzlGsffVv8ExMYTqBfySmRuMnHPmzWvFnBQQrnW2TmAj5osTRHF
oTAN31skuI3d3jJymdcUkXkr3zBGno3NGHwssN1e9znYIbmM8xMXsIxsNiK69gNw
mRi1jLpdAYsoy3r0YMdOyelVJTjCiK55OtzFaj49L95XgYnpZnFmmc+lrOKblLyZ
rKzH4Fx+s6P6lcRUOsjcOer3nNCa/Oi4CK88iJRTkFugojScK6fmXdrbRGWFv49H
V6H68EyVzuvZ0MTI8Ev+qv5TULksY9yuOmmvAXfNTonGREBTgjR+oz+wnbTCnUaY
NN0oM/Lxk+W5p+uPM1X/0+s3UFS76cDJ8eWNNl2+1h2F9HQokM/7qr786c6HmQ6h
A/usJeAOqSxq/k7QCeHPnaBsfFsBeD9pIKUZTjS+RNiWR8w+VtnkXjSS0hkGcy5p
i8S2KwqTDa668xDQrYO+B6uO3GDLLGSKr29JB52Kr2Hz89+CWvs3FL7sxcNzWHJH
7vQitt360ZpBJX2TUaLf1rZfD4w2S6GbXCrdCcjzzL/g/Fa1/XGuj5NVMwyFG4AP
/TkMASJhWxClsV2nzSa3lJGU+S2qmJ1qURib2abquTvdinNg6Bskqop86AVrmYsY
IRGSVlIjlQupqs6Zirhu0OgSwB9+0A36pcN5qjs3GeqM08ANxNaQgV/uMQcgCoLg
DINMDOWWIXOquo2x7D04BiDeB15bij+87lsHC2mu0HR9ftYQwNEx3PmTjgCTGT8E
qmP97v/ciGioVCDTH1RMS//n71qWYi5GUDXKEbhYJp3dgskQOGfnnoXAAUM6gQfi
on8kj55B453Oc5qFCQbj0Kn+PEnU5e2i37W3Joq9Ujf5fnXylbp7R2ve2bQcsZza
HNIqX99bTyUxDhUejb7ndwOt68/JpxDXYPCcO55cJZCh2vzSg2yiiFl3BvFAO4Bm
DMOAIoy+xGiUL5Axf/UhiFcFr02CXMJMoVqcADchq9FZROhkaDerh7YAPAy8k4xN
VGI7SYXiwsI2UZlxtKCTvu9s753TS7beCquBDVnlo3/W8890PIc00q8Lh7/p2jX9
rpd9iZZNRLIC1+NtfRuK0cBsTeZ1j4vyGCeXGR1TeKgdVQ4GZFF6NrdcYobV3Y2W
TS/uMYoAMnsh4ty4DLP49Qcg7ReU/sBiTRL03T12Vv6d2jxEw9lhkw7x171VqvW+
GxTdOkTqfJ24rPexQ2sZBAocBzWbWycLPfsMWzU9hHi3aBoudThZC1BDnZpAFwSJ
t5mbVSHPc99g03ttm7tK02ns5dAvbNQ9sb4LeIXmt0vLJQOy5742S2R3KlN0aKuR
Wj06k33AM1KwvQXVpiuF8hcrYdOn2510mAwV4cwxpjACklJBiU1Sbu9T4PVXTST4
SdbU0tsf58ZbO5aQIIXheJx+JjP41NcFy60YP0H9YJ8YNudHCjV8uHVO+noErKuu
CzC2GrKDEyVbJ/L8f2x9LbpoQrHzGgUU5kYl1IjLbMtpsSn1q6ubHjC0CjttuG13
o0nQGmjPCTc7M+Ntl7tgDUuP4Ze+eHNM945FbulkBevzA5PpP1j8G4ES1ZsUcKuH
4Rasu2X7rzpSfN9CW93jifhRrwa8sSnNhSLBWFxCRJg3PCh29W+8EP/Pf5KswN51
r2mREVbGQmGUIqDIZWktrTLTHzcE+p7R0i38Id8Opp8awNELP1+y+xqkY+B8UeAJ
I8qhPoPzK03qytHMhMG0bqAToFrhbJcsVF+DUoSjUGyQhgKu0hiw6pWZFJ2cI0L8
9yj+QI5h18gYxUNukCwWok8xPQniSIKO5sorl0qXS3BWMhp7ReNYceVrke826kXm
YCqTbfittMLcEqq7AwzclEdw73PKJvE3Du+agbAln4tAdKNA5mQoZVUSzApKw1cb
GOsvyAIdNmC23WBwvAy6QN3Hxt5YZTbpGDQTxS+pcqSUGg1N90473jHYq2RyicUp
pXhldIJHfNpyah8Qwza8iAWakj+qBNn7PjXiLjuK/MCdvJx6dBNeQW8akT3pXgNt
lb0kNy2sUv07PFHpw2IK0XJ8TX9X1AyllP9f3wSoyZu6BjOn7Hyqd5pFF9PZNCx0
MlIZQh4BhjMX/Gm3usaf0L5Z0gt9bq8zJfOqHby+S1yeUOvHl3sJ9ggOqtgIOAP/
A6xrOEQprS1llE6hG8hquAeamMsmfiLKpnx7nHwEF3JnMZW8z0Su77V0+mA1AdLv
vzAPHvFKG8DpbGKfAMvNzRCZtp1HArO0153P5uC3xVm117unAAYXiY0usoGSpvk2
9HKg2dqnoKraeOh2iPfsE9S39GwfCwNIt9v4cd3pfIhGQV1g5lnTRxCFMFCpypm2
2Y4kmXcyyfPmATxtDfFZZlv1eVmtBaxrW3IRtz9GwlFbVS0k4zNEwsdTFI/RTyga
bdPE0+0fTGE+ZeAwzZmfpC3f2h3IN5YsEfJxqqqJS4W/3Pb0gASx+bWCadMrRAte
GnBZqoqAWOF6oZPQD5Y7pF+j8GvypUOXjGOCdV3wTFx5ONcbV59eJy/ws7MH7yts
N21S6J6GhXT5EkiWltH9BysAFNCSMxR5OrZrQSBNdXpM4wQi5Mp8Qh8Wa8Ab6F5W
OVdi5ZeRAQq9d74cK/7wca0gBLQdxGcJR7+5NEbAxbGIiBaKLUE4GUjxQsikY6ll
9CNJgg1aY8S80mAWPHNtrn8I99vtNDNVjRWJMBbU5xHVIudegnJ0EVBWy/XPbo5F
bMvr+hbyyMtbVRW8rjP41oz4XY78IS+u0BcT+c1SNyEsKrHuWVAhuw+JfEc5H6BJ
EciZNOgSaNtAMROCh2XK/DmJWN+bYEtOQ2oC1lcqFY1xAHeLB9lX6vIY5eKrQzDP
XBM0ct/EUcf+IsBP+QCE0Z53+/RdnTf7hVuS+NxV/n0IRT4q840X2MacLL1wIYje
Yn+vemq3YgLq/3yL2dP8QcE+kk3c7ksso+U/BCZ6db2J4kNsgPCwsc6c+jJ3WMKY
XRt3drWN6zrgz8AkNIzoNjM7od0zluKPhzLCCTHvj9iV6mfq97cu5ttZ4Lz92QsS
Vsr/bVvTJ6wSwW5X+VohjKHAAz7WGiyFvrPTpc9cZXwOts+e8haAjp1soBneR9mA
7rv0APQysarVQ3wHn6C3TsJ9KOOrunmt047cFhmn5GFxdGXeMnZJZ8/8zTD6b9CJ
vY5KE8QXKywuOtaJlqdV0CKYQlLFjFnVySUnwBoqDWG0M306o9aknxF7uwHN2AOJ
nrQMQuyQZbJeIjq2PsNmWwzNrr4X6Mr2DJgf2GTZ8Ykk+l0PLFzCp+Jvgls51xiN
MPGzNkOPDRjL8ThYfzx0lPtajtGWVu/c31J08ujmOpT3kmM364QRPnuqL3jDq/Ur
i3BqYsuVWIrsyj80trGfc5RTkUCPdqYrnCI6x8IhdJp1K/WvANryjbyhZhAnSGlq
NWDcY6f3DAg/9n3nJ6lvtLJEdDEuxkJtMSvH9qwLhqNaVaD/SdabHpzAH+lQCiaL
Gngqa4sDcDA0GG9EonbBxR4jdDcsb3GnVaFaMUUp8ApXM2x12glJfxoU9pTToZMr
wprLULCGSWAxi8B0fhkXhZcMzPE2OhHPS81HcXMgeKjWibkiIe6UJLPt7vdoaPGO
sH3vjYqCqwLHJjPgMXCHF3tuOOnZtcOwA/1KvghLuYREYNIY9oQTymCRyqytUR6m
wm4djmMghcygTHGT7U9cyckWPttQR3SwXQEd1WdD/YP7UzhH9C3zPCaJIBafLaUl
ylQdCh1rS9RmUE5l94Swel50UrNmfLeHQkGo39QMSrXWXPxzXCMvao4OJNJn3iZ0
qDb1aDuxNyYYOGFHmxXfFkJmYOCkXme90QAe7IwgwawiPM/BafqhTtkp9P6dNEug
lowU4js+W9X1iK9PqZBCcdZ8rV/38dv9f/pBRJe93FqoLd9/5Eq6SQiCO4ZLfUdZ
cSgnakeeLZNvRNc1gP4Wd1xNR+LNpjf5O1GnT2OG18k6B/FYfd96EmcPXAlFK1b5
tLlkcDCnB5b7yMfQqMYc5bbrgFr2uEQq3t25z9YN90WnSdvLIe+a8nu9cpPgdaNQ
35NXDoz5sBfwdqT5/d95jr0jnk4ktVFn8FtyJyhHE4KWq/icEVKKjwc65N/g07GX
rJMxm5btgfWsdRTXIX2YoHOQUh1bJdsNVx4LWBIAFKy6Ab+KMVW3s1ux4o0NYSTq
exJgp5P8/e5wmzNmddvHXsxwBAO3AXUknuEFB12Kmy4CN6XUmrOyH4toPZh9E0Ee
sJhefQezQZHwwmiL+bfrdi2q08EOyRrE+HlwV4eikYyzhpPmGr1COxPCV3JBIiw3
PsPrdoNN2SUj46z4393xRCpvl7vAnYfF79sP6JvYSgU3XbOqFo0w4cSLW8zwT2U+
VNRwyEi7a2ahYt6s/DyfgsAXxcCsJJFj7GeZRreKnJnsHx6cX2f0aIEefQ/O2Fn4
kFpgPYnrMtX98sJpPnx9yP9X6fYshH/xjcIG8xgZDDcSiu+7XOVG3XZw2aq9oz/y
vzLw5t2XWmExrO4rZQdaxDZ8g+2Zk/sxOWzfRtweC5t8H8SkPdvXFLtIN9fQwEpU
kbBYeecCzwk1PpgHLsEkd4RXcXjHBOjAUH6L6XRi6umWTDyu5i4htIkhN4iAfCJJ
ru9X9hKMCwWpcDyWDtVfPb21dM6Zlfk6Cls3aWcjsEWjE2SfMiUTEO5vuYwU/TM5
UjIjSJzdjLbr1565r5JDazFpEUCvNnr2/8ENxWk5AW35eOQlZqeThUC+f0Shd1+Y
xsC4S6SufgzXvf3OyxE5p9FRC0V5zFjdjbGpxKboDsVqAIafbPtlb9fPgd9yqmni
C8fkPVXuxu6crYBkoSvlYPin4HVs0RM877Ll9KBPDuADrWoyT5t3cn13l3aM+A8l
2N3mJQQIdUtCxwGzhZnwTun7dlWNn/BKt9RDlsZS968A1z/d0zXO7nx0TDZWIdFu
xQ/KbMRKXzLSxUmpD9zLF0bY2BvDVeuiMuEV+vlp1CJsccFM3K+DEkapAaD20W+H
xPTWezDEek+wr2DRGVm/7nC1YxZd1p228K16ewF9v4jQEj4HO9HuYKPxpG7ZALDB
K/qdQqGfNuzezhJMyvtQc9AqOjPzlS7s/u2k88hanFZwuIs5noP3EiRxYgPeNq9U
aFXfpVDxnJIvR6l3S1ijm1uxse7s8nFRY8IStoL0oKItYOCpwvjA2LZuTNxu47bs
18CD/5pPmpJjjNMt3sT3wSKGP/fCdNE9byIKFlBLkmc38hXPk+bBcrEhS3r2i151
E35adQyhPVYBJy5dddIqfUNMFZskYrEjOVopR+U8eKTv8I06jqce+b0Q9NZfQcpa
LnpaoOkPIIStnGDqyST04N4lfdjfH1ip49h0RS39QvsiNruUVaX7aIey08ugGIei
svmp6rGK4s7KMlbm5F0yeUc2yIr9rhxBMFv9p3L4mu9TgO0fba5ryM5X41NliEd5
9A5RB3H5g/U0OJ5DEXdOQcHxwwmbr/3yKi0oxi/fTsmc3mE30tk3JH+BLAsI9iEn
cf/8iMsCbepNOXZ/o+eYnLd60sdbzi3Fce2mfhk1fs+sN7Xu39KKv/THCNi1P4zX
cWINtgcI0FQS+DopzZ+SPM3ipfzPZxGFk6fBhukQm40R/Jyg8Wo7DZ/vgyshboIR
hUTh/8JcFo3mRgAsaN2LLT5x1cxmePbHnpmpJxcYdWzNIXKswh5NGskPL8al38Bg
0R40p2/fphBPKg/28gOt/5eo+AM5A9rpl4p2sc+7+T8CoeZ6QppxlSOGWovcIuU8
vAy8tHV7nAIy0ZIGK/mRtdNjk/yZY8XoA2v4XEDTug3knDBFw9hAlLKmE7h0O/W9
KHm7Zr72OI1koH1KDaMNwTcUxsQ2nUu3191efkrCk3+mbp/IBLozp5gVJ3rIziIN
6Dza7Pfca9Dcptcvti+OMfR3SW0TvTNug2+jBY5JjXI/WZibvuXj3WCAjDoTjp08
rvWnSgY5CAovaOHdK/p4x2oBAnEmrdt0z5k1XO6RVTEv9SKrYSiwU7vxKfW3q+zz
kdMIMtVSMA/43eG/54GAVhCVvzUDXAWmUW2HuQYdR2cXu2p95o1ClPYBHGZisIt2
802p5b4JPNXbCULgGs7yOGCQO5s0FIr8zSlqLSyG1OfNO+tGD24rFow4lN7pxqpt
ED84Z+v3dFIvRKVn7u7iqV5+d5wpta9BosLWiDUflQ8HF7X+q3f2Gw1Zyl61Fw94
5qgsJWV/z6ZFpnpghxrhye62k+2z39G8v7NoRVBNiLjoEnVgid+Me4blXhUbBxBT
fLrgwxM9sgVy8UZoaDW0ZaxVY9UhiCIquGXNEeJ39A57AKOxsje4G0Cj2CECteFh
jjZ7JLzIB+IhwX92XP1jujLos5pSCDN2LfgFP8gD5/BL2IUOh+TLqJTqHl9WNjqe
OSySuLaV/DsLwPKFmuWqPb61ZGoiEKbTyTkjTaevH7DKFTb6TKmmcLvwv2UbiogO
fOiMMxXLe3N5kHBir7E0zk7cAXAWy3GL6aSpDjfFcN63306ljaMuk2Ci5pE1DfUL
IPnlbPL/cPy6qhbvRnDwpKldWg3+uzoh0xxaPs1zMO/ZT0JA/n9To/jfjJ2baaUf
jkqdKftwtTydBV9qu8nizvPCFoL4DVLUZKyNKCId0STRX1qOT5nTW9qKoAgDclV1
ce/TLwA3xYCoqj+6OEle9fvNMpUs07kS5ywRD+l/zwb5kvZULqQQQ1Y4GslUttoe
0tZ0+TiMLaEd/7psKbfeDEDyrWycSdHA+5eRaUWORGgt0JCd612ekgIPTsAYa46g
xPhJvGJKIXAzg5g3uQsFc64e23KxC80yiDU6bK7Q53uzxlVyK3Ht0YeLwsEzkPsU
TVGv9a+eaeCWbGW26pkvwAuSeIs8Gc4l0IeDRrlQC5FwjqRxSixHCWfhTxs2SJBu
m3UUDOWC6O/uyluyyRE1EUSmiQ3mulb6hZ7bjTCVk1s3LrOz/UHI6sYzXTZdinIE
Mxt50DVtN39HF5HxlJm6Sm0gQzw8w07s+LfCb6paETLbIMSMskuKcFDdoAqiKuz6
j4br+LijLdutU3sfclN8Uh1JD1j3nSuN6xc5faBUkQ2B0pg/xMtxuuKj/0sgr/kP
qt2V3ezVZMGkFrCLq1am8XVxn1Pj0Ki9lDRiWKno1kWtq6DD4WJpWJVg8q1diCQ0
OBk01hg78QdZM48GlXIH7mPpfJe+1x60Wno6IlWWn56sS38YRIwSW9bUwlj3t8FF
k5V3/J/CD6GQqpXWxAYx3tUOJOEn3jMGrCi6xIh+SLOxJdxq4aDIQH0mIArf6WHS
qojXwmqnXD2nZ9jSgMeymTUA2eGPG01eU7rOElBA+2Di4wvVCXsNKc/aUL5q3RaO
iVoZ4YB3dWBlxm9mx9JRkcI4dRXqhqR5boon95x493QXGRPx+eCzMzII85B0asXW
VMUP13FZUfzxp/p47cXNUkhv/LaSOK4n65FV5XX55160wKTMsddrtWjpvPRVI211
Ank0MpIsrMEh+57p4Y1g8MaP1RFWxY4DC0fJRMUQp0H1R2KcNG28Ts25i4/HeF0y
S49hm5KScDjlYtLbe+GaUZ/hIcevDM9pCo+MzG5sK98TCrfz7rGoJHUAS6k6eLCm
TJVMpVrZbJatlzA7bfvLRMX7Shw3nIAPZR1FjmlPlR6QmIw1EBpeGAmSBh7TmSOg
fUMI6luj9BI8JcW3l3M3sSv8QxdG1HOnJLRM9uVFTF8oxFSQ++e0ql1gpKlxvWc/
aPNqbwWEchqa2E474oy0ExhwN7OiGbAzKlv72FZ8oPgyq26n+tdeXQd768XYspF5
atBBZ1dE5UdPhu7JsZRDA8+VBUaVi+Uah6XWSYZuu9V9fIcianiMm9vE49UokNju
l4sTvyLsBuGFYTlGUYuD1HeUn7tNLDPjz6tUHD5FwSUz2/i5EStlftA9YIoBxt8H
nXQ078xJBqBjULK1kUJJOB8bWNg5VyvTevH38QHEKlGN59ecKZjetlvLAMtCGzKm
2NuE+rkbV6TErxlIHHfpe712xvVQZXkEerrDaPODxsAY+3ceQY9sJXEuIf+icoGp
g6GKmQUl2Jnxr2gSN9JhY6q396B1x/hU5IBRZOmXUjVv6riC6pNT17iB329zEk83
9SBtxUMuSmgEXzH3MHo0DSJYy0fa1Rgm7tgo6PM2CLsr/0YqCqbo+K5E4W1p0iX8
o5tIBFBu7ytHWD32RBn+HO+KkiNJmhG0yeVQNJAb/Qp8H9RFuE/rNgpW0TfG8NFN
9HQheNplgnuKkjNyuHGAtcYkHdJjMcaSOfp9+Axe0fziUdWuBiRdzqLGTLMv+yHI
jcHEgp//W7P56aKTKROcpuNH2p+USVI0K2aMQxQZyIbZcIviqK8uVIVH/DI1yWL/
bDJlR6rBsAesG6LIe8uNwp9TZ0fw8MPzUVz723y51OBiW/7QB1e3p7bmp5J4RULY
QtzM+oFAzioWeCBGYhF937N+1wBmmdRIwzaz3VXlXFZJ7+EiU0mGEsQGx40rxvSb
toPzPeD23Co3umKICkM+VBXmTZmlLqPG4enmnAdYFnnm7oxlRawC4JKBegWfo5Sw
DuYxBZAmvgl+xw20hIxdJggNTlOl9970XL6UpsVxuDm5h74Yakj35p7DGCUP4F5T
R/6ID7P2MxfQVSsDJSkM/KXuVPIIzeI7LiuRI9bcBBDuH08yrcYveOe2rGKUOOQk
qA+W2M6hUtquYbVEFFfgt4p9ZyoZkdXIpD55KotpABo2WvyyJPsFDEURvol+4ksj
5C+27c68o9Bszayi7YZ5jRA04DJ0VwkKVcWCj4cZVTWpZSOFlml1u48Y/htH3TSG
azLzTjJNpbbkLlV2uDGt4C5+BlQDNzkrSenYGlFhTYUR8YqVF5C1NUKx0vpZr99S
A7xNvnPk75jhZF8LyAVHWP14CbTjwyYB3PApdltd5yxn87SLoe/vVmfQC/nTIGI7
ODw5e3+8O4cJigtndj1hrjSxViakiQv7TSbw1yvmKQHsAuoXX23o8fkGqSusbFpP
aNWf/2W03H2hWwvZe4h+XWmQy9oTWVLoxpxJZnrIKbIF6m8rqQanBkv8mEifOPZa
mJSRq2tDK/Qhc+Np47OtLODFAKsMU2IKVJbXSnlazkITN5fb6l0M69KLY8Z/6vJF
XPjq0c7Eqa8cu5ypcOWKY+zqwz7dMo7ULx5CQ+X+YHb0dMOEOYIJRP+nBcYfkCw7
wDXBXsxqHLEhm9UjpX9jPLtQTzrnJoUFOtDneuDx1fOzmmoGj44eFWbnD2RSZOV2
wd8VKOHbW3b3MVPGHX3PIphUZHEDqDfFDXgYUNyh4+JLBrfjiqcyrnhsFVtXUEky
W8nrjlEBMrhXSoWDIYqjeJueow7x3imbRLzSW4ANJL6sDbw/spghFdKdk29Dokc+
nKmeQPVYEBCgK9y45z4GlFn5iBcNLMEZ95CGWTfMpOHDU6SCSx0qsh13oYEVGuZx
jwyqorso4NjWnaVT27woOni5h+f/3BOuxtghePR64rWfLpuCF8SebYWY9Cb8th+s
x/+PtAPsPZwPiYKusz3QADqBKlBgD73gllkDv+EF0xqGW7+l55OK4a+hnnboM3SI
ghz/sKLK33ih4yav++ZGt9vIrASzyQhNO3VVUe/VOo0pd/eZbnd1eVzH5URhidTF
0GUShNpkRlJBDa4XfZkPEVga1Rq0FbYVJzNUrYsaA3a03B/N1oM+tDdSLEGwrIlF
9oD2RmUO7VuLmlcYdpMSm6Gkfi5LyCroD+wXEfBQZYXw8o07qdVuUzgI3SD4UWU/
+/5uLruX1ql17VgE45TBnFYDkPq7NT44kVwpiViWTjmjPKINAT7uL9DSuALdkHFJ
+HPFQZuAP7c+LTYNTTt2M7RRGNtLrF6HQmhRzeWhA67plvEwv/nlWvjRaxlPWRhN
HsUaVdP8vrt6YYfVHmkKUSI+eXvnJ++D/6ZfQR11vkPCJOq+ENxb+JPd3e+t6hwS
UiYpLM14tJuzwL6wNWbf6wNSl66PPNVrezgaBTdcJnVzS4g1uHDXoskVHdjAlT68
0l3FIySI1/NX97B8XUBwVP/ZF/e8Sd4rwbKDNRV2QT2s+9lTtlNlSe7NNhsEk83j
YCE/ivbNPJfqtAo0TibPR4MrVpN+GNU05UES+qkg6ktBf9FUSnti/MhsptFqPKDE
Bohuu2+Gc28BgVGMvcY0DEPEpKVabcxqYazWe70XzgFBk/WPs9sOV43hf97UNNbG
96hw7v7tQJcTK5TmKv4G0u0+EDwKDkzyxu/GDCVUD+gdJPEAqVKndeYW7bshY3tT
FD5ytTOugVcvcsu7+zqPD3C7IsfGfqUyvi6W3LltVld1LIHV4MtAlwENQV47wwdU
1+KY0QrUo9Fd/pZQE3NXDkLwDX+NSDUtkYgX5mKgDsJ23Rk1H4+IRFgx1keaiDVc
XTThHokK0UfAAXoz4ws4lVYwi4LHrSAz68ECmK+PqKO1Z1OP4wtLXkQAtEyLHqP9
+EPVbUD04KVm1DltrzZV5pN3YLBHpIJ/QSfbq7QI/kzbzVM0PEWjBTJEjN0n3yxK
dw9aLE9UT/AGhfheMaxlCexQc27Q7+vRb4KzEDjYyB8MYIEVBhnnVZWB3QYu+Ize
DaZy/V2n9zF6IufGVLzmcGo/qERlu6eWrMilwBrVZ6b3n6WcMYTCJrQcs5e6McOx
94/EVPDZ2sEztrFiQiSW0xHE5OYotVbd4gWiPUlcSoFgjWvJztpeIBFByznytfOY
38V/aP37MJrCUxgxRzcv0ObKEM9RBsLT4fQu9gDH7/TPB2/qqMTRXtNHvvHpx8He
kWSfeLuncXEXBeBVjdkxZl3oTYhNwsNK1QLc7WxAC+YI7SHPsg5WtqqsXLhQe5gm
5QpiYADEy6VPbZKceQ5Os09YMN6GwaXuJmAmm4L2j6unHt+tauZEGAm3AFoac4Gf
UNIcKmmsMStIokQMOSSrqzl7+UF1ZOrAknifV8fjq/mpYVNB9dpt1RbTFSEOANBr
nD1w5SXEntjcDyK9KWd89HxoXuNRm8MBH5J1ERlmUylAm7DcUXOZivBzu6+J4XUC
o2765I8AWvpvcv9MRVh6n35uYVyxaN88MKMNiBfP82pWPPODTIsgYkEuvf/B+pWL
uy0zDKROE5dQ9zT3ayMrCU0Qy1z0uNJb8M70qIIL3P63biHB0E4Z1av+RSL+l7Kk
epEHM8K4XHoY5QGuqY/mc5sgAuZ/1fjp0yKD3Qpe1bf/BeePr3CYxrqrtxlZW9uT
YyULMdMlOATkNIHYWT7qDOX7d1g4xAY9gszmOvxnS2CAUv1sxnrLlS4P1wzkIAA7
y4VoqmD2CaWSkRSBq7uoe0bi+xVcDrn3Y0NA4A7Wbtpg7bPQC3ugnW44cSwlTauV
/gYRPzimnyebL6VYHOKfVfX0QeHtAfjD7xPZBw2jWsNxshPmVY/vITv52SjXXo+f
2HRzDcrc6dGj2aIGYLBLWUbIWeZHb+TafVagdiyTdpIB7Qbqte/YIZzm1kDG/rcL
l3h+V1E7sChtHnstFxwFv8zshburYpD4R78XUdaAgGSBRWZ+dtdF/qV5x9+tHfKg
AmcfMG7cYiPXGwNvaCODtVnFBPOcCXsG6MMugFEQHOlF6q39wah9uf18tbjp4SH7
OSxI7JKxqKY9QybPFkCcdisTTQGs+t3PT3cLXpJLjdlKaW7I8Esby7MNvLa8MoLk
hDwlpn+Vd1DRQagd/FRdjbiqFNzTdagGWY2PeyccI9pYsbTBeM4f1WcFqG2rhhDP
qKoO7fSFwHcSGdLCXYmg79BK2Y3DfCkffaBOfeVNWalA5ohGLeUA933rCDlkPlC9
eOsu5Q4SPVAPn+MZoZ270pG+ewGyqKO7oW1p08I2OcxCBHAncQ2DThM5yHF5eikn
JCuFZKW0Vozn6dPLxFllJELYCiC6x5Vx58cU+d64i2TmFHWLs9lAByVu3MpKmExA
rUCKrzkMhTceV0/sWssnL5hTmC/EPDwpA5JESaIFF5N2YHsR6xz/ucmaUsGau8Nw
lQRyMgd9SJG+ngH6QDaNZWYiyFEt61GHvaNEONb7TASD6kTwGRYKSw1UF0wka/tb
8gqyNP4mcja+H/1xGUOxNnzr+/YjjphkWHErU2BOdLgXiuRp6WYN+hzbJ+mhaKQ3
7P7af1sBnFIexyQWVqmHkY77Rh5OTSaPsnqgLf7LhZkUVKRo6R/mePuxoTJ1yy/J
C61I8l8eeUSzXfW9HIZlX30vSFAzVNcxEepdDJkl9tbvTEZzVgfAc+f7rcVtfJp+
V0ejiUu1G09Eoi7sE2R+JUQ+R2gbveMVPflQqSdSpPMmgjt3vQpuEznWQaHS0jXn
ZATu7oAsfOlPGOCXxrWbQ3gZuLDe/5kVVcYB8uwW8Y32cIRmkLJGgkD/qaRjY5SG
tybzJW0WyfJmbBWYQIVtlgFsGqUR18HnTJ+7lhHrxR+I0BqP0hBqifCS2AUEFjVx
9FX8GthJp96G9wkXGEx8dvnB6qNpUHoQ7mFwP0K9bAcN3auHC7IFjoWSLK+wukmb
1PEwi4BJ57+TSwSUC4DAH9JlxDsqv46QycUJzcDvtBXieEqica5j2KM91QxfK8Br
nzKFKdvVnMij++D7h62i0vTrFe3tSgNtiqJmj1zw3+CSiciiJRLVb6cHzZLJ0FTr
TLjY0rwOY+QexPzmqf2kUfSoJkYWgBn/2mh3oosU8atRqV64t2N5D2X3Dkyxf0fY
DwBZWgbo17a462pauTIFNWjUR+6UNaPFMhnplriBZHM3XBco+4YIh+H4CASKxYcP
mMNu5FfP1yQaj/ZEPDtnC8F51ym0MYYXthEl5eYLqwB85xlC7QlzuKUJheKH8Mc4
vj2btgB083AkESgP0sbGakcFuDlv3tUudoNYOr0bh+tzPRycW1Vza+ShO4p07b3o
FumCNUCC20bdJqAQfngEHQTVD9mwncXOVlMzs8Tm4ZDx2mFEBCkzaATSTS2lXiZQ
EJWjEbh2tfZclalcCAkKz6wwSGz8KhYkvegf+A7k+HkLZnemrtq9udOv/GwyMXgR
JcEDEaGqOShrAoF7CPPxAMh6b3+4FvFEAFcSztNlxVleGN//qkv88FSNIp8QpKZB
MwCAApLwinGaxWTxCS1mxYLdsO0CN79JtzpnSCIajfoGRMBYH72ccjEFX5muEufY
DePlu1Kunx7H4jxUxoS/uLY0XEcmoPsb3SSls2zY1gcAaRZfPnruYBp1i33xJ4NB
o1ts/1w2LBjbrN2gW3Ltc72Hk1h/9vjWJqAVns6PISuTD5atoLiKKm4E6DiozoSc
nagjMi6eYDhIIaJJlBniQaX9sSOybe76ioARepAGkcEbdEiRWeBCAAND9ZpdM3bO
W4OrTieeeFtAdgLz0Xvm7aQ7rxQKAv7nNjb0HE24eLAcxMhcv+d38/9Osts62r1a
JD3mlnw06od6I6KREm6UujqbRWtMDtVO44G0oX0BzDR3aqCVR5Y36lc7zXB7l9LY
xECbdNT7jFUBbTD4OFdiTPjy4/FN/jM40ZbPxCzunJ/GmpiRmgf1kzwX3x/0FKkr
ztpSGZS0y5skYgv2/GMF38prhrz06W9TR/A1M/bksx8SJRpAng4wgl6JTYB9J79h
9DHP4iXLJRiaRpsqUCOqms3nm83zR0aXUJ5Aa++aajyLXvhMZ1dDDCsZgQ+MCJOt
PCkGlLbR72iviedwD4iRA62t5PtnVur6f3tIL1zsau4j2SW2FJI5Bh6GUJ4z0ET8
gW0/kZKnPRwLEqku8yhFlVda1uTPL2M8iIYIxIPV2nfi5yCvnM8N//kX6KfWtYp9
M/5FtBL4KmVKQkqgurcXuQtwZY3+cC8u3E4rcLww0wccdkMg7If3eAfNyVqKT/C4
KFAoRwf299vk7pXUSWwQQz2/xpUwW3rET097+Uh4Bj8JnTy7yzYHw3YzFdsfClaO
6HTQjV/cImBJ3CZc6zmIO03pivhzFGkY5JOTfd5/zpd9vqxTG4feVHXsP4lSpD8W
HrVJ8LgWV8pm/YwxcNAmH7sZpvYNUtnI0DDIJmIN6e0Jpl4pjkwEsyQvd0a0PTvI
wTPCPvhESFujIaw+DFmIrXyl3270tXr7UyJO+hvGMnpkRov27uah8QI5kMPA6Tht
zoskQum3fcng+1/xnlyu9EuLHHXZL1lFyDqPIq/kQkQl1Nh6EF8zJiNumm4CUb8h
cNhkOBqVia7lCdNO+azyXkWLTIEq4JQysZqo6b9ml0N757OCO5flCs8cNIiT+1DU
aN8y7JPYcYrgP3/1BDszDGNCY4KV13SLG2sKZMP7N1ZNZSnqB/gDrdflo7KD5lMD
abNuC/ETk1ZCGl/cuQUpNDlHhm1Rz9mT/MKP6Yii/H8U5taZFDAMFld7sXt+tYdo
ozFd2z4Gw5cRpmZvRPgphyRzxyY7QTVfKZh2w70C02csNOhydoIt7ofOLdn7kfBU
2szTMfDbRQ8frmqw4/b2tkp9v7NJO0vp6xIfwoFbV+SC+M3Q4MM9E9w/NkOeV59d
ZE1F6E6zO77lh8m+AfGywJYK+SiMnO0ao+qAvPQ8humAzyHCb8o88MB9CPndtlda
HpLxopdtrR57pajDLmTvh/x10jXhPs51RUm11KRhLHgTTR1Bc2SagE6dM4ZXCjiN
3eKMsrQLfEAjIFtlZnXOD7nZGQ1U4DRNVyVDGfSXFZolcQHyDLbw240Xh6h9kTLN
FBg80RSDWX3UzIPZqAGTbJyrN06/fIWP6c92h0YexXfK60BhW8BaWYXEa2KJPw8L
+jkCN6I81t/lMYVf8aFpargSOWwrwMHKB1/evnUsiXBAL4XbgxQOQa/WOKKIXKYW
hmSnhz5MbHoPp1ebvMOVKZyKAQ8QdzwYaEbRzxjm2MPnF/0JiAgTN2Bb4ALKqQ9K
j3K1hzJQjsj6JTJzRIC93ysOkommdbnVkFKuLvXzb2JaGl80Sdy3/Oq6pix3Pr1y
zZqAo72eOJbyOQWi/l2zBlm9jzEGfoTOTNPOKEMZc/ZrEDGVob7LOUVGC1PpLQwe
CnSPHDKEMB5cZ4B695voarOdw5GTFf/K7RDiDPkC+kbF07qA0iMXOWPvDavN98aI
E7eKJb2s2py2+7/Y93445trK39RnsVTTL3a4QcMCK5fyjJOfHB7YrqgbnDukHJms
V/4NHMO+kOYTbA2HUchtfkl5v11k5wJ6PA63RAk1QFebkHbG87yzzzz5UOo82jRf
QIPC8H39rI/JzenrSHUnajPoZ9Y6jrwL8x7ZshYbwGSCfBBnopox6LWMNMCZQWbg
xk6AknQo+gRcGrVEC+KeWhucZlki/CNUrcTOE/6yvxWj0ssYRjs3vcC6l73NkUbN
euO7tlWkJHPBtPaBzOaMlVxQmYHBi88rikfSTfG76Bajd8Wkhb8G4B+bWp+EwGg0
ixRWZLUfxQr5Xmq6eF9xZdQbmVM50KoK83TuBUo9QYChu8dJZ4n/HX+rnweUsOFE
WMztvuqaPMZb+Hg/XPBVe0wMo68xxclrkZU+tr4i4+LtqIhEi1azqI4CSJ1RbZXY
OsJsLHK3Ixu3C+0SDCSERHheiWq0cMt9IgV7Pv+HOjF13tEhpObcTEXps/eYwGiV
/vprH5fImOTGMcDPxs3G2bFR9ZDk6ma7KuDiy+wkdkjSHHAxgVmhsQnOWVG7IVRs
izuClLoI2S1o2f0dZsYw3ZYcNqdYpJ2MpHz+YE89HX7wVpCC4lPp/gkvwx+qw74f
toMFSZDhvA/hvLDC8arwMr1MN0A261exyJAAIeLCtsZvbUk2eFSjGVt0sThQrjru
b3rOUY+gjqtMrlfhISZ+Zlov/xqPjTK7Y/BQFoY6ukCNVAPWww5WXzoBumyQvKUx
g6Z1Hz1HJlUPEoZ0WKh54Ke6m8zKoGZ3tV5NE+YqCTRsb3o4ZRafKR0BodZEhYYd
1o2HmKkmJOAVeHLF/n6D8iWwb81UEO2hVT8WCIn2z+mtcnEqsVpYA2iq+7HP6teY
WkPLYIHs/H4vB6oVk0Ysj6X0oF7I1XNbGSdotHEZaqavDRS7AamRXeQ1yjlwafhD
fljAsoBkPKdBVNN6jv3RNIBQu/bDJwnsoCGC6dvkscTRp4AE1mKTzx0xXRjHsa57
VS74WHEDy1vQ+aR4Z2mpKbZjY5nwSJlED6JjxM+ORr6s+P9upmf4Rl7a8raouoRU
ZKx3Wb4IPjb7VHkHAfmrMUxqurQAjnrcYZY8MHTlIXuXkPtM8Bz9N7BMKEq3IKZz
LEUTawlo0RJMT7xtzZQJNo0wijq1ckhm3lJz1BMy/CVhab1cUMcLJcAmanN24dm3
XEL/OnPWzs0V1hgYs9TlnXI9XQCYMAeQAv9ZfOjFGZVF7wQ3VTFv0Ih2gQpa6IMR
TRr9ou8xuREQukeRsuIBMhG7kDcNQaNOVJPAfKlC46PGnaMpsE37aUC2U8eZykyD
6bvJNhwGiv2g2LtvPj3jZMIDnuzqUl2FdrHlruZmg2Kx7mzxoxBZg4KhdP+V3zhr
jFrdgGTBL/5wcBqzo7hF/eh/f7ruiXY2kI7tsC0DnLheMB9PlGX91Lpr7T0Lfh2m
pfPt9FycC21eoo32pHjZKu1RC11DXW0yxuXXVfEHlBgq59G8UGY8N2i9AnpG5lLA
09S8qIt7QMrnRwkIjCOnComH/vzPjHijRmzZGdj6VO8r3E4aTz00hBs/uW/cjUvl
IMcegX40lFpwqCbnSLjb+V4roWVNswBkLX6DpXh2ajT426mhQMkInQaVlHaG3TTG
pK2oA0N+fZg8BVgFWIMY1PLNNSrcQEJI6mOC0P7cupuv2q8hlBncJzMEbU5KWTt6
e8nHhl0msPaI1l4Rc8vI1I/OSuVnsQ8z3gGhB6bfO1PKVy4n1n5OyQb9EeFFir7G
ZrMqToXmotCTa0yUEvTlj/X72a79VxRaFabNS6z40DSVoa/t48Dfp0slUX/Vf5St
rL7bUBGrsF5pCHdWtefuucjmiuOz4ReFYqiErMTonK7NfaJUbnY0wTZC4zFrXS0/
tmnPsQlu22uzUj3AKwfOzCjgPLf//0xKVxbfHlUTe5r5Cgt4XpWq/My7lLNj3uX5
VjWIpZmKOb//Lnzh5xHv6Gabmz5Q5AR4ar/WJAB7tFVi1n+cWKHNTWW1XFBMVYzp
KyE8zfY0xNGqAtVpj2jteEfjzZqKyntPr0f/uTkd6Y4+D2FFJlK4/hGlq2QL+0ly
3iIOnp3U2q4agvCVUcl2/MyhZvPJfKAWjWdAkLIUVwIfYdjldak5qcybfaMDX7yL
GS3VnDZbx0Wi1vkzCQ7XHcT0FwUrPHuyKPVBTy386I+uZKIhiU0L/PdWoN6WFdlI
oMGbuv7DzU9NyDCNO5xW7pAeoANqEtmNsiyzY18p0ICcrUXl1mssJ4eodJT92YrE
32BVUnBcmBbPUF7IQBLTWLFCOcgLVYolXqF0wiS0JCzxoedQBXmMiyUODGQBksPd
ZTS3m1dqDMRBJa6Fwn/5S65+AfT8XD3K/1c36aEa5C/u0I6y7cY8Nsb5oje5smxr
jmpBLFhkHPETSn0cJsnXWqABsysyukoB16pif0Qq77idYlBI4d37dUQWqx9U1/C/
LUepxCAscizoIbpDpWo7IT2n/ICupVlwp7Rm5QDCaP8w0hrVHLU5cqE6MZSi8P7J
1qE16zFJnAmTGcgd1VA9gefJjRrW1NGEeuuwt8qE1YaRF7QONJ6veM+6uUbLFZYZ
h0AqlPszvwgfnL8xPQ49gqBJ58REvf5r2OljNFZ1FsMHd1Ronsve6iWzKfAFGknV
nfnI+gRGAdZ67E4YNzA/rLfLwTSDqXF/52oAL8YKb6HQUe4A7T0UuYBuDwpgmBxh
F+m6loSFULlTmdlf+/BgAB1Bvyk2g17aXmkEhS6caU9Ubpj0TI/cEmauMizf8sQP
eoI39xQmCmcfTRWOGe5dOBUxA2p59ih0fgbfIXQpdt0WkATXFmGbVaxFdI3xUV+V
eZUBgAChLFFGkAPpNHTbZPcoZJI54w/Q27STQZATTjy3zh60SBsG7L/Dah0P+8f5
xFXc1pqcU6KrT3FrLltUhGY3ZmDpoWP3wjl3INyoLcTZ8mxH/yFr0tZxTDAHHT0C
XuqWgZKYKWaQB6udVv0HEaH66AYOW9GsQ15+blPntNKM2kLA3IxG0EVYxuRom1q1
ZL+z/mudzAZ5exIWTIIYbDjq/SofW4SodU8bjoN2LuY1oXHHnfRFaCW+z0vJqnB7
dr4H9ni6tTsgh01WVzDG7fu/3j59UiJx9vNTPAGAuhyyNgeEHit+dhvjIOxPvNb6
QD9ReoCGJU7Zr3MSugzFPyVj5jr4pqW50YooQPbKXQyGD+usrcwPlJlUvfzcOj1u
FJcZj/oZHHXeyBFDwDWaZvWFBqfFB+abX1uj4jeJr92OyIcq1/m4IGYp0oz/Z8g8
Pazl8f+2BJfGZGf4arCB3Z0l00gCpwx0oWDwjMaShwA21Uw4n+TU+TNrw3U2CAEo
wcELc0mCVpnwDgRvt4Puk/9n1NlpwoTL2YRWDxkJGoE+4llRlTtinWN4FMNO4/NM
IeP0vMf6j9AINx7U8FawbH+G/mx2702DTsHexY6p4Z6OTL5XSZBnwLbNOulsV29Q
gJagRY1lP0SSF5gyukjjlxm/6nsDbPlNybaDnjN8J3cEE9zTzok9RRBvPdVbL8Pi
4KGhUzjp2ToM4k7eWy0NAVBY36XKvtSbf85rPcJ1hyvieK0oMytKphKPCOV81Pxw
M4053iNmkLFgKDgQ7YUgXXZzx/4drPWeD8tPavq/6sqqbgp6HvvwB/YmP8fMnFmx
1yeA90DnWcctpRh7eoe9C7TDPHJeOyKwQh5UzkGgti5IXJ8OJ1fh0E/i+9aTG1Uu
vqum1zuzFWhDtBtMY6dz3DffWkD5ShR4wFRaI2baHkfIoyWQzgH+vv5n5hHhRuSe
Vg8Wz1RtnJRftwOgl45vkBznVGxs58YirJh5OD2YgIEdncankY8+UjCREzReloX0
hp5TMluhARJnyPaX3DPLNV7mROojKV0L66/kknMNg24Fgt2Lpj3TLPP2QPOAe2H4
+xPx/6QvjSdAMmpH0xxKmL95nRlBSQAMVerebyuv5R+vaOkTzhaEDelURR01pryf
fu8hsyiwDAZdmN/BOGOg+HNVFVgTBpp2qZPM8BHry539KykSXTr/6VOtxOvdy1d6
ihXq4H/8gcq6FsIkrWwvYp5ebB81jBCdtQQxwxLGuMnadn4KoWxIe1JuYjqJ03ep
6PysNyWjS6x/0pejHU3slQh5ZqfJo56p6LYDaSbJ2WKQ9ZkUXWvhE0HmYHenWPkT
nHTBFcA1HPJ36VndBUL0gemhMG73iK+Wm3sN8l53PrSF0jZ5IKcUq1emkb8dX8Dg
BJJ/s7sFMmvboiUkm2KlzgSeM8l5HgTiA5BuOJclOjRjIgnugIOelTtZHV2JZED5
1DhkLRxTaQ7DmEYWF3kMCAoVoPxYjGgBhMPPiXldja0oMGrs6ItjFOHzKk2V1L6d
/srKI46npbs5po7pjbHrTMmhRm2Nf03Hqeu80LTaI1LMZMwGJeO0gu7+SqPOBZ/J
xMhum1RA0QrCB8cHBGAaNAwq4Ldu3kqKsOO2i3S9zWKqUotbUJa5R5v7X9OTxOdP
tn8yxJONLua7ubcZXr9LUO5D96YBUOCxyv27TfdR5XrqQ+bhj4YQk+4jntz70CVy
WY4Ff9Ii2m6UF2/DIJmlyYa7WAV08kT9ElCaEDjl9mDStRPs2QUIkFkf28LvlGFu
5koI+uTNIFsybPs+9lFV3l9828dVOG38d748G92Dg5Tso5D58lTdpRX+wD1i6ROM
18BZrow4tveyy3Eq3GRY+KnHniC/2k+m0cM4SgSKNAVBGU29rJx0/tf/kjJgmdI7
c8W/wBQMJGjbW2PyjKJoDybcE4IObaENMNwd3cVOXsQrbKsCv63UyVr3AWf5QaN6
gndXAW5trq2W+ud1YYQIU1zW9cFNo3uiUMbKrI1IOdCmI+ENgu+Y+EICahSnDsx+
wP82+VgP5GGe9HnlEyFxI1idUqVs3wBdN/Vv+3Fo40z3t2hcT7TsjtpgfG6sLQkG
iTWAWX2owQnQ/Uega1dBTd30V9IKZjqyiXL0pvJBwwmTA9N1Otvdw1CQK3xSKRUl
qD7hF+dvvXuj/GTzfRoRPwsQo6zUqfULNJVhwahwEQFDWgUmuMDcvdouDq4u8w2B
T6Fpwm0hsw4908xHU2AjSK24O6nPUsPOnim/RpQniHRqDyJcmNavxF0n9rXk6A+n
FCAOQ4k6APSJoKRpD7rxtEvP9QDvjzmUM2BWQyAa2y5fd2aUN/C/oVInPNremWbx
WFL9PADdxR3uGCB15ocCli0F+Jc9NMyKWez4vmv+n9LvNgGuI0HRY8jZasN7NHdX
v4n2dQluTq1IS09+hJyU7Ep9mCAy7mDDFGDlSTVbBDVjz2oq+/727sEmEUfh8XsY
3Tn6uWfB8SXePz4dUUm72Zt+pLlnh7m45qIfIFvpTDwbnnqhRr8NxQ3vosPv9BZx
HE4tQrm43FZouvkjJLxpeczIxQREQqfBC2Jef/M9WhJ9L2rSs7VBByWqEDZgOa+r
eJfqq1DIH4zLNtebZEdt9S3HpMVtGNTXYKHoXslVQVNWyJKU8GJBFmhmv5sU2ccT
g6qia/8dHaaq+QLy6bGtW7hapDpMSf3UGob2DtJToBKoyVRw/lOmXcGGA9Er3yKR
Rfg8qzDp7eTmRIzzPVy3Xunomk59L0SsJA++MiEV4ou7Gvc8+rcnBQwY2yXs9M9q
1oduvE4CGao2wPJQxARjGj1wsk1P5e5mwJttQaMDxWaWvXrPDUyU9XyP3CcP41qZ
EpzwE6OwoQrVVCZElN6RG4qgG1BeF4tdhaVPSegv/pL9ddhJSBYQsrsgkWCoanRf
x5vh4sGW0NKNUJ+LzpYj00d5rgVmt3gADsosdRA6+sBptJIyB6F8FqZ35jjatVo1
+wp3qQTMi8SZZswx9mLf0gsON2BzupHaKm8UWklmbvUG0PTJoSZTdvD6WBSqRKyQ
HuKr2emNlcc3kUNHeK5XQXRIQwy2duNp/Ls9e5i3V1Ws0ZJdadNqiTb1H2hszHP3
Qe+VNGv5qozY0D3ct2u2q8cFLIrnrb8VtHbdUYx42Q6kNkSKa3zU4XEZfhEoxjaa
Lt1eHRnOhzKZozYSkUtDRREfTUECyKmr72n+oXdIVu82Nr8gQirUEfqNEw53CnkE
w2QyHi8kgEUJaoMhe+eoQ831he2/pZQv+X774ZEJnIZejzXmflGtFJt/SJw0vsD2
lU5VK/a7VLpyDiJXMZciSifdjbIpG6Eu5g3o97OLYfMp2BpnJFf4T8WRHDzC0v3O
rZQzyJ7RyxIpJWqUMDNfgde2QAE8u19AUyJP4Y1YDGFzoXNpa0vB/sC0TQdrFRSt
3v+DI1nMqLkkZfAY7rkG1V+vP1dmaqblOWuAehjhobXA4w4iB74cQp1g49nD5T9H
4PftUWPMwYfZrINGn3Mz9BqnqqL7VMqR2Coajnxx+ndlk9C/qcuVsC1g1FnpEzRw
yq7w2GGify7d2mxYNtQEb1wD5PGmE5mzzvyJK+c7izqQR59OgYmmcrR3ZBs4xI0q
sId160f/+pa8+3nl+UsfItyzjdFLhiYzcYT26P6NWSyCpL5M1DwBzDaJm93xOvIK
vpihTxEJj3dYmxGJS2CnQebw31Ob9kh04OdaBH528tR1DFq5xxkd9WHz3yPZEc3v
5l0Iwj1CmhAXL5HtfYhr6w7XWCyZd7GCXMbBeG1siA7wzIlxxznsZR3lTEkmddQe
mJbXcQLrG+sNFB5Rn4U4tZ7zdGbbuKtuPEWZ8o+YC7Wtty0vCXW76u0hJqtOmBkQ
skY6p3AV2n1u+4Q2OQtIbWVgAo1Mf9kyP8tFdWRMMaic5d5cdTm305407SZ0B/9y
5GpX7TwDuqttHKbqEMw+BDZc70NVOiTa8Qp3GxGPKsP6S0ORs72XdC5jskBXk6KE
byJAj9bI8UpFgxZknaJDaZ0dBWOF0vGqJO4355Z+9RjKfrAEpW/xvs763eDUIian
IXm9w97WEYQcxbtnOUWGbnWS+mW8s7qupki9sgl48NXb1cvKQWoIjLKDDHMvSCZg
RYw2F7HM0GpyxFBWARrlQpf+StAs7xjOtbTMNWwQz5jY9ehBtxMzsdFkw/pUS3QG
Rd/pjVDBNxpNfvmQUd0SmTmP5PhdqBPZOLwTzas54U1v+Sdxh9GVL7TpFDTqlZ2m
2qrKFPk7ynGUVeDsKQLpAJQUUxw7U6H76h4tlFUoK29VbrEZTglvkkvvpcDEv7u+
fwujOKy46ehyNRZ6bBBi5Gucacd4lDx3d7m3m5XwKplz9uSZbgflwVEhywPZUtAF
d3lKyxrs8ooEUqIVOvyVn1uAWwpSnFZAd2J+Bg867wGRx8KjoEoLwuuyvJkYY+7s
pJixsko17bL1ME+zVxZfhN9/XyLbm4Va7mVu6rnazfJNQ7MbZYgoMOcCV2DYppsX
y+mGdGPOLrt/vvz0RwYfGsI1wEy3+Bx+W4+8kjMTRonr9JMNwOXy456K3IUzYsFg
FEz01B3Zyn89AtwJJnuJr/1w/4H9c/TgJzJi/+UbxWnUJV1x4CTHEL2ik4S+a9J9
STUec940HGwlibremI+Jsxl7SvrhHBV4qkkTGalJg8SOuOotI2bFPkigDPTSO8bX
IveYD62vy7IKIFEzpp/8BX6OKE5mL8P8WlNjqwvgIbeyvkynn/+uhz2ko2NVmyqG
FlLxtNkKJ9oyJA46FLSTYciNYc+VSJ9yj6Pv9nP3Yzv2W6D5x6+OrF6acfAmouw6
PsX79e6jouk+NCiYBBGfZN1MWawMq8bX0PNeax+RQV+MAB+V6NLs88uA3mkeWz76
mi+BONFnAkOotl8WFt2NOsSYDIUDPalB4luUcdN/1tLeAkw2BNQzZAXXaQEZiBDw
qfjWG67sRmsM5gi9HdS/D7ZwF8osXmsxL49/k46BszkeYwA08cU50VmxJLd7cMHX
go7sDohlfXB/o2cOLinpFDd69hvUYuRPjxEwC2HPMzlhLwJHKMlJJb0ocd/X6Zrm
yWbIc2Q5SuE/0H8A6w6IByj+77A7U7L1UPgn5VyiQmWhRIhKM7Jx6Wu219agG2nv
EAdfXc790LnUGD7qiddZNCOAOcD1GdMcR7DxTorEyihNBquyHWXlIWAD1TIyTCPF
ex7He/KkviRXnbZAKVZL/ipRkzTo4pquZWNzp49WoXd7EcZNyGd9qpl3KwWKzb84
tKBqU9ktjL9Gq4qKnFVO4DO1DuyxMsBDh4yCM0hrm0LCkO4cFORRzld7j9EzGYLU
w8RY75cz0GfY29FVWH9QyHrYGJoXGHODsPKGVV5C7iqNYUeTni7of27F3Pti+oYn
cHKimRsOY5uQOcuEIZcM6Ezh3oGy0aw2nBMzVumChXH2y553I7yd48UOC58dIpmp
AIGUgRu5fyualhjKp5RcNMqe69rZdj6zmezhNC6yHWPtvcfhSRN1X6qsLAJk9jL4
eSvXnUg5gxECQgaImxAi74kfBE1thuD5ktyfPBD4QTp8GYyYMdcY+s7p0tYnG1FO
7hIIVc1Kx2JHSB0NKR5tYVK+rDFbCiAQRNLSdLfVM4gJ+QypOc9KRlSu8jldv+Gj
X+8uzNHhAYF+V2+rJM4DMAvLw8MczKASWZf4msdAOTWDhJR6maWRC7VsNYlyvOe5
4Slgd2OqoCLe58tREFgq62ZeDzKoY+Er7i8a/ZprwiaQlB6Ssh59q3HlT1+lYrN1
MyaJ0l+akHhgs2wgTTPW83kENYIe7zCCkWlWjhnRSjPQblnNrJhsVZHoN00G9tSd
Rd92CMV2NcD2+dVfuxa/XUtVvQUtW5GAaICJMVyXD1h1KP9K9Ckg5heotO/MExWX
R438OU1wk8Y/M5CSDgBhTB4sykBkr9LPXS9ag6qC3Y/z/6rW/pUxeDkn0ErxpoUX
tQJYccukXZsYZLb19bG4mgqv/InozRi950TtbmgwFQMoMYZ4ZPgkv4AQT3N0vWkf
jyqhrrK2Pss21yimNw4DRbYBGHUO+RYTXsqwGINgFjvfCCT9HU62gNFPrDZYad4K
4bN1yyToLFLbPSqtnx7o4bOTsP6pxtTvprI5VVpL8WCsIyYnLrmnzB2/Frf++z3Z
VWpj00fFLIv7HGivtfrwRgVInVfKs0Ne/HVpjgz0JAFHcdpb4d6TLerK7f2v3ekF
mpFUxdujioYtf1WjAQz8Mam1gElyUlzIaRMm3CAfyE+SwYm1LW67/ahj6H/1mLbN
pDTtUBJFJr/WxXQd6yIwEsF4BI4vqQk5xv5Ngjp1Rv9TDwj5xlmj2QM2PDHkpSXE
rHs6jjLP7A725vtBDXcSE/D2QUZvgiEhBsrsPMQYEZBDqXv5QXITW615pXHmdkiO
PSogd80v7Yrfs9BjUTC7pgWBRBorS3ag7lo+L7ux3FUZ1zcchbQK3JdJbh6SC7v0
7KqPnQpKPfA71BU2xvBNZnfZBBftPNEyZ+KcASdoEtV/83NV1emfQr9+KUrt7xXl
gw/mpXN7FLTQBA4GMTzuPmcSoctuGOVxeDfF/lRMwO8g455iCRCZYP0auZClg1Ov
Ez6w/YZCx/ZTKTwB/XGrlYtUZi18eiNlJbOn4CYpdyo+jJTyWwj0UGQsW4NTbShx
MKo9803usi5B32xinPOPu+NqHbTxvfaYb5Ij97R00G6D+D9PksxCmLLp8dG7fyNd
7E9U/srFX7O2bPJytgnvNgqWCNWbRQG5emsrtJ890mN/zVG11+Fmn1byqSRMCpQK
8U+mCAkSY06aDFssHyRm/Qv0r3YkoaASUuJuhuLbCno+Qlflv9ml2ilDDEtD0V7v
K5+xPdKdM4bxtwFZSc9BRrno5TcKABs0gLlofUVdF2Nrfa1l0cNcUf4absoUa5F6
OI2NWzdCJ17HUBeemI/rNYRJ/INinweErjxCfZY1MZTyvxBbt8v/oRf75cU8cdxL
b50lj7WnEGYiHiikU0LnYyKiEVtCq3YfYWch8kXoCYemj/3FuXLD8JVwHImm6wxv
Ckglb8TufhcnJKUaiLOMeolAK2cO05SFxuOLHq1i2bvEX392uDHWWAICCM63b56w
Uv/67u8xNmo3rx7rXiCgyUHXaZioaL5Hrlmh8iecG4Q7Cj9j1uGrQDiBH2naFOe7
Os4byYpLLkVkEPs5RVK9sz5P3TxCr9aXH65alfq8CjrVL6/R/lbiIt8LAMZQy2mC
wp3tnZ0MpWtU2tEj9CLFgx5/WGZngbowPvJerDMgc+Gu1ft4cuDprIZrHqnlKq3R
SHbDPq6yWwqObckotR9sr6dQdBwvRkRJb/TSaUtUSNry0z8aAE9BlKU1c7OHEV66
CMscu5F3bm4xPmCdZgqvFgajYinL5xO17wnjKXtxgVib/t3LmV3bagL9d4tKKw7u
DVodBFiRS/DqH/l7gkatG6AKvPr45+CbdKohq3J8N6wahJHqDH6/HMV9i7uZdryI
aGW2y2BnlTu6QA537aEPGi0XvOl71+WDXKS4vdf3mER+3b6gAVVl02+G2ViFwUsa
PjayX0qI1ouVRjuvZfTSeoeKLt4EXhGkU2J090fiA2NzYPIpVNCawlbTdHLYjtWm
w2Z2lFQ7jhUpweIDyNXQ+hFocwr6ie8dLtAVchEL2lJgW4TP0pIQGqSD6QkitI1c
DTHewVyFkzFA3oUEn7rWi2rfYPTQfGdh7WfgDIYrWi2KyrqEW6fNMmzNqFd66lqB
k1+raZcyKTbTi94uGQ4GJQvBa03ktfU8m/OCocB1z28SbvlOJ/0Ph9fHQ6MpB1T8
QTkEgmR5iL3PQo3UlytuzCJu1IrBHmMs7L5OtLlV5EG7TsmfB7rj0Sm8ivrw9Dht
XaFfeu0lMuZHc+ASK0+m6Ts+yZO0hIR0sR16N7W40g10UzuqyVYm1UGswqPrazsR
Qlw6dnPaKJelNXE6f/HvJUn9ARqnthITod9f12qvKPIZ+N7mem2fe1TD733XXmP7
Y3KlBuSfxkc3v3PMOiz4eDIVpSLQUJIpNd2B7s2mgBRk0jpe36Yh7WPkf4ierSk5
npeiNHvmUjMlu1KIgD195gTvr0+FqtRiyM5zg6+FRQQZZqrx0R6qaO4UPI/E9VUV
2p7Af3VnoYDxlVHUN/noz15rk9+ZgYN4b6UC7kHvxBInApFmIJkoSwFA23Xm5jDD
EpKLL0cutbJ29XEXFsfmfkCk9O9nl4JkGadfGlDyPrfIjX2xlbakdiMFaA2QGpHZ
6QiKX5UiXFQICGApbLI2B4qBlfr7k5Dg9zfKQ5gmE1q9Ht7/eMSNVjwGfqqjYqn7
Tt1AnpKZ7bFL9RMDxz4CWmJtjkblfKs2EYp8inU0HnAo6GKMdtNDO/1a0PjkYJZ8
0AYWg0Xs4rnC8zWY5sxH45EyUfmXwhqiYpFKDWJFGjaYsmF+sSUGdQPz0llKr+Q3
lsYAAaG1uLD00A6mGsZPBBseqPcLWyxiSZY0To/5LE7ACJ0Ktk7K8mgEzbO/bUXL
MoNhzPqRom2rnwHnT62E9cmJknU0SAGaj4k85fFR7v2NPAmBkenLBo1P/5Ruffbz
0VAyXfq5gEKVA//36kL1G0RIgpX0kL5aNxGByvKrXbFAQAMGINtFfA2soHfBUQVD
I74G1wRVooUbjXrkvdF4ZKYCLB0+LQb4xjEYzst6+4LFwxo62Dp84r9n79Z72Bk5
ca46EoGOhgSg9aCDXaBstVGxWwQ4HChfc8740wnBAfC+QW6+EeC3NKUI2xLXE3ol
A1bQRStuYyf8h8Ej+LT6cb9UQfRmo+S64cdDP1N6ZOzFnRkRVQ4mXAMf5kFPnWN3
aFCtS+5H+qxk9AfzHAVoBofoI8bE8g4WhTIB41K9xRV3pIRVxpIGtgbgCbMeUj8n
jrhGKqbHssnGZB/TE79Ad6sa2pNuUuE1rbSuZGY/TRncUKBVV0pV30R6i8V3vpoS
5ehb0wS5ZkiGEcmR3wtPsG0JMn9KFbxRRpg8l0B/9wXJ84egYKcSMqJ8le67iakh
wTGzGXdt5Jr6URVmINll3WKbTTbJ/0WKmBIOSm0oznisZFbIhSWDghc4+KHez8rV
jCf6fUonIeY3p+alCRoH4xqDcECoMo5S7QD/jrGUjvfthiEuiiacOC+U1NpKSQCD
VY2hvV+o/4O4psenc8B/L0mt0DNu43SO1hgr1+fazQ7EJFsUQFrKBqxly9DT+5ko
XyAs7pwh2tR9oNN+nhJrzg0H0Z6mJNNb38i0v+3T8emGqwzz1XNZ/CAwuda5RW8h
Z5Fc8IkQTCL0MMfefgIx1DNNEYYfxTJbFM6KvlxafpPgUFI4LtqkrEP2Mq+Td8Nb
uBwJMiBnjtrVJH6EtFAq13NR/sNXm0F/zXqXv4vgqgwDJczP5PJ/G0WFXNxT/4r5
tkJL+GIObx1bK8CmZrhRv/zwvmKzQnJ79HA1nHkI+1N5G2/HeP0otWuMNTeXAOCL
rWZIjMqVES7RthuEuAF7Awj/TaYRK+gWrVrmxKONMBHDfwz9C+muRtpzzJt9ytYJ
7f2Kz5JwGROhugkQCY3h7Pj+93F1gXJTiAObqbVqZyW7PhzQ/BmJyyeEmVAA+/A1
wwbl5rX+GOlrbl2UP2Mr20NftrdQXcIzyxDkV3t3tLJB/chJ3lJ65tqIinh9TUIt
LYt8b1kJL/b5y9aqHgCmaU8Wy72emYWdP1Wz8rzxId69sQy2vAVpxl4boHx4PYUO
Wdt0C8of9naJ7zPPbKqBulj11gPZIwuSxO7193XWoTKmuqG8aQfFMcj6T+D/V+50
tsS5g/raLQXhiYiB6uLDIuWYuGzFMT+2v6/Ouos9ZDwXkkCkxA5YxiiNkUkty6ww
o7XrywsmRRzCX84soScnaaDRdNP+pDOforOgQwZ0E+zHvTh6+POM3QSXBVAMigM+
6anPIngxndfRuFifxB/Zlh4uFpr/iZsL9d6Aw7SLTz0gJYPye+Cd+tL+pPlZJLli
sKos6KCBrionPNdVWCdwkxgrxCyRu8V2im8hcmO/YkX0nYNoFXZlQVE4ym1Kq+4a
Uf3LZDxlHIuHyw4EdvnaJ7F9M0qLkFQb6asAtxLM532MOu9FquUhXFEehX3ypzC2
V+GbCneIFYvLGOBoB06kBFmirCK3opzV9AS7iVew8mlNQbOC8wCMhvQLljt0c1eP
aqRkXna9Z+8QLSkX0Z+a+oBZTfBtXLur27jC0qjsUVFJ3i9PDF60d8bRnkumpKwW
PIgRNA4ULiuwMj+l5l3dDb7rplTG79Vf4apvZp7d3zu4rvF3k9KTAY9qNqcUaCTQ
F5JhHgViGRH+fq/9lLamHJ+DLuwrgsatAD2qpxwtFQiagRqQRVUIKdMbflNvRP7g
ZItMkM/MUeCMpHB1V30UMkLVdSv5HMuAR+PdOsY4BzlMi1BQ8Uoo9y+VgLfsbreC
EBC+Mpu+4yOLok6g/Kg52DQaAdsfPcL607kB8fCOyuQpiYZEhu82kjO9HVDbkhYY
/6ndhSMDnxpcVXo5Oq/JYWnip9rnpmLGBe/LN9pf56QsNtFb60ptUO7b9ymYiwJf
+YpCJWp8pC6EcOls4BzD3nCaMtbKBSUYt8esmYuXd8dolf+KEKXY+f1+aoJA9Lfk
Fbzd6ublbdtXFK7vpgxdN3CjlgqQyjQSCVnM9QjWPFwj8cUTtoF1XAMdrHQaDRCJ
S9rTibCZAgyA+X8ZBGQ/Kmx89jVgUu3Yw1lEHWFA/xSx0gu5rvM1Y95k2b0Q8wPO
ezaQ796EpXp41mDE0+DpaQuLLgXKqBu0bF6RCHQYTaqg61jKT58l7bNjtE8Lq9pj
iQ45taBoT2zbtL0St7w2XIAiTF5daMrdzS3TFQ+dq497ZtNCwK48eAn/KQZ6fMxD
jZmQGGu7FrzgCwRlCmHIZk48tzzKjMoFgytjsJ6MITiEPjTXjIObnQmYnBCnn+LK
2Uy/OcJK8rifN/+E8OAcxas9NjjdW9y9SOhXn3ya/E23yiIXeBa09aFihJOfp9tl
idj3eTRXlX1W+SwUOpBCC6OUy1mvuE5iWh00oc2PEKVy4kIr/MRrBSCz//rKY2ji
Sg061J17MRk3NVb2QP8587NHlkoPo5OK8KtO4WBIaF10E4TwhECR4pyjRmzh0j8S
xiNwv1o9oxa3gfKBv/XYpFhV1Q+JpzptT4IP7jwXz7y0lZ9cGxO8JourxmDQMddu
8z++nk/sd1n5uzXLZxbD8hvvQtdfmIePO5dgd082D9muK2FQV8LHjh3AOez3hlaL
blDBmQjmUDIl9xTExUOCPEdU3opw6Z3jIDo2XFBwe21AxkL6XjKCuK9oOQnrEO+W
CBWkNGPDSHM0UvMaGuyIFedxOGl0KGTXIliKTM3R9xLoRDlmrza8s3nD+zyZj7yY
LkmlWUVV+r11HkXRMKi+CHVWxtWljEPcDA+E/16CGcy2H6omSBKu1v5edlhUl4kQ
Psghtr6tqkMxQSM40wmJ87Gjs7aLis+rnXEDex9bhVOu4326hWfoDQLraHc91vm+
UzCay2kb0CBhJtLhxgcrrlvMolhEGy1U9IfDadORBmVI57O5xYNzikSYQ4ec6N6U
Bo4zyYw1QsYo2coYgxjGqd2BIq9nywjULQzfAw8iP4dAD3+W3Aj2H/rumN32uTad
2zu7KG8CQJKyKlAkXK27zIGvjRyUPR6EK7hSarykWIRskWlkaI5Xt3dn5qLeW6yS
YznMP7RtSB7eqRocO309ikeT7xkTuEsYY5LZneVXIa3/5L0VGuYWc9lYCnTfvSa+
z2MC74aqHgyIZnsVjL0pIdfEmVBezJO7WUNkOuYXDSsWkp4VYpHz+A9dUBqxrhPa
g78BCXFwFllw0ObqOKKUmvlc/M3hR+x6wY5rT9tNvKwcn5i3ovub1MxgPr+jRg+v
dnz320LwkE4R3Xn2WMGkFEcet2dYJhmGcIK8GbWqEeEL3A78JVyvWtT+eVXbix0F
IjtZjf96AGRz57TF2zcU9cu3oZ1hj1ko1Yy/2KuESXufJ+e2njf+FjIsC9K7DwnP
ITPhJtVcF4Ns6QOYeMGihz/XDc7TWGSnDia1fd7Z+NICSEZvcbgyjZ4tvrlRlRGQ
vNNfBbuaAfG6ZyASN+RQwvcN6WkdHsZFAhTs5LKpfs75Ch1lZrJ7JU9BWuobSIi0
fDYocnJiZjW5RTwEZfs6Q+7TrtVk47sKGcb/7gp4m+OAp6ADX1xaN0EL6XIsaoDb
6zaUHPvrxHiSMWGWhd8cFromS5SSLjQwPuK3UFGV1l99kMosFRH5g/lbCOATrial
GscqCaUPgOt0DJJL2wSQwTNo6GWD16HSXW2LPnOT7qf4owQ/hYQlsxkkdkiKNh2a
lN4NyYTU4Hxswpdwvd1J5ZLdoyW9J6dpNgEzq9q0lgEox4fYV1mOIeZyEq5hqMkx
wa9c68RySKI1uVGdOUARI/Kq53ulzthkIOOp+UFg9gWTpSUVg4YD84k9pwUm52fD
U+E3usyBj4aDwwLRnCSscZfzH0VFUDBmu4+Vm66Rjhb0bKz1qxw0JAnxReb2MrUu
9trh4inhA+Z90lbPnAUMsDbRabxoELo2dorCiaqmsdh7ooX8QlRfmMfQYL9e9fRO
IyUe4/aSYengFSWd+Aom6lJHKQDOIpubCAuVwNijCty5VXKyt5mztmdaStOAMhy4
FlXUMu/1ikqfXBgZeydKhB+2HCYpHJFp+h4mXrGqn90QI6HhkgXPoud41GCJjnVg
Rv4MiMMTo2/TkP+1VPoAYakwUxYUEmfVG3ynOv2fggjEX85kIgjySEQ73T2msZ2N
tEFVqg8wd5bRMVCljYjPHxO3A/8tLRSDgqvPa6eu05LWGY9g4mj8TM8tOanhWB3S
CJlTcE80fkZzAFQca+HINvOrCoHxwLpKL5Q2rdGZgCAfGbDAB67sE3iQYyKRTLxR
wK614cQN6WEasEzsdGbZa1kpSNzeuSQ2trqBGK0RXknDlvh81AXKE2/20sAvIuH9
kmJYxlEXL2o6jDXMDV2wWJ27yIkKC5cZMBCapC3rZVIMJ5+iEojBZHUuIhZdRfHQ
/vZrJZzb2iQFfBiZM1M+64KVAsimJMNegxQFocor11HycvR6obhyWeB88EyB7lsn
2vcfuY4McfGHiMuMMz2L4NjmcjepMvRyH6OfMTgu9fjDMAkNzxrEtf0mR75EsQsA
cy0LRrF/k35WXFzC8a1NJHEKPIBsr6WgmVDjNFfcJ+cgOd8PseIiPwKtCrAlOVES
76fj9Yl4CMb6fM7mcR4/f6IDAMZuP8QyssOBB60X3Y1Mn9CK2qiYZ6GqMwfna06u
uhLTru3FMjh8523KEAoaSsZM+P3bZmlNv/X1BoVgKOirObcAqu/gpK6fquncIWL5
6SIQWaADLe1+YE/rbNhyy/Ddr01kXEjyar9NjnxG/WiO5cXYRJnv8dki4Gd9KO/z
jKi24eyqrvBK4DRUwRbZCO8oG5uD1sdIvPO8bb07iwsxwL2y2E9cpP0yPmum0HsE
Bb5om7hFTe2lx+rCdNSUsVE6UfgeFLgxy1BqUjuu68/Vao6gNPiDazB6C/6COqtU
NBXeYHcJ85lrMbirkuDYeYMjljIEl5tAM2XlI+kac3q3cStPEDUD+A+VYytBy8aJ
PaNNfvhlGC94QP52azNE/1Yr/STBjTrXlrFdf10RVRXLh3KnpIu1BMycwNv9zir/
9FMweJ3EwARa+qoNla/5ybQqjXeFGQcgCK5Oy8tF0XEHgF1Hdx+w/pKq6LeWBrLE
onGFxqf4/ubq5rCxHZOjsUNvF8ezQTE+m8EiHzlaxhNzrTUHQNkbRz4Bd3nJpNBD
4U3ApRJzagJGe9RLlCmgQAhW1koaAYFgBkXbebfmWc38jV3+xxW4KmlQIWwBXY9H
hxT/xGAOHkoWuRMmqTLEvVKsG0KjhBtBnQJ3/T2ZfKgm8c320BfPu2Q26WMlpDAi
4PHyG89N1byW+to3r3DIE2N9JhA62F5Or+d0HouDsoo4d1tgnh/j0uEogVlsVjyv
fQLsyPZ10nJJsNKCxYiRL6Sqqf2ajBpkgDDy96Kn4ME260XARA/iMHqEgCXj+aun
qgfMMHTZzpYzm8SrXTU5JjS2RjLGgKmJGV4W+vV1Pl6iFRi+/PC3KMq/qDMWjunb
MhgzgJplTGqK3kk/q8HXdOXJ4trrF3/kfV6i/kQNf8Kh0+fKSBtlTJJKPdT0BmIK
KR+Fw2jykltPlpHi/wpzgD7JQiJGthD92/A7+vMQXJmAlyfI1HxRDF+ggJ7S0YwW
YuCsQvAXEmo7zBlvjFGGZobp5hJP0gna9S+0GTteaGNhegqKF0kXtJI4PNBOT/CY
S9aN0OayIM1IWiqPOJzRP0a75DKmD1dDRT7LO7y3gxd2uo9nkMpfuQIiDqNdExIU
vbVPP7rx1dZ7Aift7y9r+pxQVpcJVOAFbqGxhbFlWB7qyTMhpSP2fouIe1qts58V
oetOTCkVz6qc8ouiUBXR7555kElt1btVDjzltMIW0rEOw6wFEyT2b1DVqWZt8fl6
c9Yyx3jnoKshHNHhz9BknvB1OdbX9QHzLuCGEXp9e3PGFAulsPDD+OeCaSMP3j2w
uU8vjZr6zh+O7/nsEcajbplntndGKVIxbs009iJQRQoDpsij1c74h09e5jO1/kzI
fYEVJmxHnh/kwOZhLnBIrBlxEvHCkOw2QmD9+ouXwh/TT+LD1lCv+XfFcyFTCJ3c
5WSYMs4Neez2pl6+e/eXyUT9naYc/zO3oCcL0pf1guzDSOLUe+wWYAg486Ah3Y9J
Nai+UZJoPdmVfUnOUYAMJ+S9zdhgH1m8h7minfRbJO7TPB0RuvWrFLRrJmI8XhI3
vT9o9OPlCg4tGi4fLHLnA2zOEY2SLvNnX+t8ZEo+Ct729E/H/3ti2WEChtOVe59r
SyfhPqDhYn63Eht3xVYZaFQM3IzlE/H8whRoZa9Auzkd0ZfPlmFHkEaVnnWIQjtf
k8dtNSagma6IPMNGT+WGPSD3yxiPOQKuKoQNAJSJ/t9KKTYC2ZTW+ubyqDaimf4r
FJg1qly4T0jhAdG13bMYmyQrRAqEnPuP7uTyJGNqasE/UuLTPdqZd8HfWAzGnpsc
myTGc3jbPBB3/dsViSiUCJbnRfNqNJu4wiEs0wMdGR1a5Le1GdMtB4hHyejZToxk
8BYSlIGiJuXMj8fK5Qs4VzH3sM48/Q28cY6fviARR4nVFZgImvAlSJcDePNQWvbV
d044kmpecgsWZdFOfzFpbQVPz/4LLpRrVu9qpsYVl52Z/r6DpoPXQEC0rCuV0pSQ
Q1m7d4rePTKKuxCn6GRbXpRiHNCYUcZsHkzGECfSv9dXahuCr09x48Yv79VkV09V
UISYosIV1XkOWl2BkxQw0RwoK66BFE5sFUEKn5NgKasJhEZauNOwbCfloI4doQjW
IdRjQ9G5o3G21jWh+wc0AJxLlwkeU1JJ0tEibBIlvbi21VyWOsbOuacNzH4GtIHK
lTe3gf/sEn42vVGQqh8LqAhsrhCQvGxRK7E3tZSJ0h+Rs9MLGliJO+1gdeD4C/p4
Eyva4reKL7ldq8UKosCQTzcyYeWawec5ZCTFfFF6ypJ7DC5sn6crBl8Zq26eWxua
OL0HowN6Rey4UDFk7JFyN9oClfuU973VS5vgdjlZ9EU4I01tfsv36sMYTgs9Vrci
xz1+zLnWmS38hRLH78YFi1lt+fjQ3Axs4uDl/+7lzXd8KqblVTf6CBlpu5mT68vW
7A67fX4GiNVDOvjJ04Fg7eg5n0Ny4vM08cEwaG+yNh/amYjlRYVmVouEYJnhVTQ3
2cpK7B/02kJ92Q2y5Krdpl8LDp4ku0k2hCtluw6foUBDlTpiPZkFxNNK0Y1M0vJK
rKXwDYiHpZ5X3l0NMIhEnjiFRL8k+xLFWeJ/mkHNcDn2zCmXLARmwjMIa8eoEsV+
U7AojTKYm2+KmwX0SZc5g4wshORJqkzdTQ7vLZ5TOVVoCTYyYTdwiluY4DDvGZ3u
N2FCHlqaHPtuAEb3BK9tleVvNUVOoHf9HTzlGD9SmPTe3i5wO1mIUiWO3fmHDO41
9N7YRiStaJTwyu60PHkOWZtnkrw35ooSMm0AHSZ0gcP/M1W5+DSYDxlghotRPwcD
7OW6hLKeorblKcEAV40quqrZSXirR/1eTSJko8zRCjgkX3pcubbEz3/TZTtKrDCf
W7b8w5ZNJbZRWE6QClpX+/rpkcMirWJLdWUa82ICP4xpULpAZD6qlMh9NRGsCVBT
yEmmcrNYjHmIkv1ys+y7RnuKBGm1xjlc3Tm2q9CS4jWp/CSXLUkXXwuRZ4FobLUN
vCCQ+N9yPGDQOBwkt8fgbBEw1ay7TXXCrlvKsMAwOOkWjWFDG7j2EHjXzv/G7XAQ
JBrvc+KAeIs9SPIc8pwo3eBvpnEQYEZz3YFTh4v2H4g1K5uE6wDiTxOq6BGJPrUr
4UekLBqFT+1F0aYp3yp3g6X/XY8gzStVOTkkCN+pxQB/xU+tjs1QvRO8FawzRGcv
T++Z+lAln/lHYDbrYRbZYBJGWO3Oqjvzw5xDDom+YFLLroJyFVPuec4+rSl0j29C
I+aDBIlEMHmdL7kI8QtxOX1mfYHX+Tn+zql+u7LLbv6aDE5ugmoOTk9jRZPqJBhY
Lo6LEUFgfv0Zj7iCf+9r46oxIz++AlJPA1fdUbHykeqATTHL1VQSGai0FTwP3JKR
wu+NSA/9CCaP0PgTOoJ04Pj6t48hhEEdk6tZAK0al8KtgQlw4PQayALbUBIi4GHN
WvnI7qrs3Y4W1j6Ifz6mTEWYJsx2qh7AP2lOHawwXYmk+CVG3ekl583RtlYVo4zS
QFZWfjY9PlvXeDGUk/x5Tb+F4HbZ3esYz5EEOWiNId8T7DzxzX2HcB1sYmU1heCF
92b2imnGk3HOGqUSyVK95jFD/zD+QH95UX9QrI785INJaGNeCnDP7JPp78n3iv+6
/CJ0IlrjI2SAVbGel+wsl7sCtKx7QpA0qEyywJ/HL875e1oexPOMY1EFzA401Fd8
kG6PoNmLuC8U/AKYHTwF+di3MV685d3DJVrm+8Yt8W/hZS4MVhEi+KsZoSsJvkdm
UHOiJop7bmoNc+8hyErJimKgXppRAa0DvbE24yVjQQVw/QDBMrBY/MDhSLFw67SS
z38Ty60Q6v2Sjsew4eBiYbH/u49fNRHrIMPHkAivFQQDd6Ks+gzK3zgM6oQ8125G
xI7IwOznj0znmWGE9YlF3Zk6fw0hMCKisINuCwtR4EKdtS62iyOZvY2jmXzQYhun
zdM6/GblIonQje5YJlH6518xG75NeQwMbjs2X3vXrTiJMsm5mDDk7ncBeW4/rAuO
Qvs1zAYsvg5SrsigiDagL14etyxNWzWMFjN82G+xGYAwmhFECf/wb9ISWLacQUyZ
YgNtBEdVKZ1+oK1es8aVK1PplvgUSZNhuICPMiRiujLeKxXkLTRCEteHGHMwYnvC
iAVjoH9X1768xuivSVMgKa+ly/IubhhcZE9pUYEu7w/4Rpaw2zj2h78mbdSMBIjy
NO3ZuMDmiLDlMpN6L4t30HPOGOyZ7zEh47g7Lml+W3dHtNl2lk6VuZhYRlK/Bkus
RxxL+01UjHC7IL9glC0AjG3L6Z4GNxCFUjtvA4JBWe/zc7+uLx6ztYnZLw6vj8NN
tLXT6TsTGVlSWCuNqsh9mcmmLvkqqQS7rOqUQZyK6AT/35uUx79qXQ6GptrJ8yae
j4kqG3JZ0aIJbLy7VPm0LILiGWbHOfVN55oMGtYcuNHZpC9rFoLmfKwAdybtHYdk
0+DPvKyayrxphjd0mBsox23tfMfOoM031aEeMyfR3JGs1ptA3xEjSYvzfZ9NYweM
rtmruTQtaXHkCI7LgYc3hr74Fe9QcAZhJ+M0Nt5vVvYWUjhw63j+h0SxJQ9eaxjV
h4PIo7Jh8nm/t+Xv+zAP2HZYOo/SbECf+3ktVAUb7i5BeWPJNJF9wS1yhrj4AjJ+
Kjp4IPSWbm5K6Sn8bWlZeAxalPuaTu7wSbccsD5uSGKu4sfW0FQgHa6Gyk7vMy0G
r22CQefSfSEDQOXz2ZWylQNgpefDygAPbAZB5RTQK7PXY3KpmiDh95f/kUEc+phT
rtLeT9MCJHDh0OMrX6RjWmHmPxbUcIiWMlaZjojD0dGoU84Mlf5fmlYW+p/6ArPE
Yr00MzZVFdlKvvvZNjmrnWXK3BdqFZ43C/X/BEiTeYF5VNBE2WIop9sBEvnE/4jw
E3FZ81JYX4CBGR1kOyGMwY8QOESRLlGDmlk9J29TO5uIWbCHJ0iIrRq5fMUOMl5O
gJ0/2bdKt52wg3K1B4WDi1LdDhHbbLNS8VGEWW2qbqgFax+Ug/koOifHQwHSOZEF
yv//7ukmjgge/5kNg4HThxY6j4/6BucYpv4abeBTiEQnzjgysPipgYhOLwgZ7H9v
Ln4f3vBP5AUnc6UFPzrQlks3wKeTNaeziFvO7olFavuI7nwo4fCJPzLEjp4B30UB
NlCWYhQVWPpU41hfDTZ5GbuSQ5VySEZCh5/D3ggpOhkX/vns8ra3/vJrBOto2WSs
oK8ZDDKciTVpnESbxF72mQH2GRRPoIjKilOmKRQzY13A28vU0JDA4fEbTPFoijb7
5TrxmNh65AKxaDbEa9F/WDmPCxEKpSnLqj8672BbOt3du4r/rpp8f6dXOncRmUzD
/JBMC0djRtbQz37CLC4BSfbEf88S7zVhUUOPKtWJSFjRluer8jYnZk7xitu9mZiX
6DzY5ObE+rTHVmk5LfO6iqnqP5bMbgpendkGMuzhIow4hkuSbjK0OwSaIGW6T8Gh
CplunxWhum6cJf6iSGKlJxAtFvtEHeivypQHP40MUTS//ziyHozzizDduCdTJM+P
0Nz9dapvDN0pjEgi3XlS9Wz/jGk3CX+8c+QYnfCDwyfYV/JCuRY+OFyWLdd2hHWq
3vNrMxOhk2WKPSzaRlbzgwMClqHseTYIeM7YxAiK+fCVBtyuG0HVUn9aXafeyv79
ahxtYyuciwEgVHN3Wvdmnf0qMUx2KO0t4vmkO09TYONOekegGY5KUNxDONcBC4qK
ZrkTIVeQVsPgUAizRhG1tPREONOeyscuMXsG0gotrfx0Sbbbhmgecir3a5TX+4mq
CP+heZdJv+ct9BP9p2ko41ekVqeO2qk/e0l0BlUGNMJQpa1aVnK/CR0QHRvgWM4V
dG1waCcG03zQZg/xkYvMPGFy8cf/meIGCP9ySoD3n1JBpxVKFI8DTY9bzrykOhrJ
sXoEs4NAw23uQe9LN7HqeUkSVEBPnMyDPgl2EZns4z/ZBm+BUpeg8JpTwpxiaWbn
IWecei5auHpIBShdA3VaVuJ/UexRDvpIxnBLqq2KdszQBJA7KU6LP1tiplz7Okj7
whpVwSfCPP3w1tAnAF4GREwrEIn247ZcG1HCo5a6jIDWl9TuLRl+1UogpipHbeZI
YSWX+8RHmi2l7zJ7v64yK2/sQI6qKHKgJUbW9mGLVBNx5gAIrnjHlQla85FSzPL7
dVAaES9nWCpnzmN+NL84qlGZlGRQhfzsxiR0OVUKVnun3FB83ONXzKgrtAJaiwMR
3mZSR9dVIOSpfHBAJ3WcsX0M4X2GdMixiZ31TI5PLnw0ID9gU/LnS5akHMCtsZTc
A70URBIXZASZXU5wL+2rDdehd5jaX/WUpQYP/IyeJbWD2Tq4hIJ+rizdD6wKLN06
fbCFnKWVECR4S70+DoDowZdvU8cn4tDxsEyKtRFPqPGvkfmnFxHKeYo22BtVm2kQ
qimiND2Iae9FSLqXNbr80z5zlop+q4N0MpgjkM8+I/QieqjwnRl/FzhdZAjQbfKn
8/+1avO07gbglMwfYTjnAT/5Kgcgta3dSRPZsc3QIj+bmTy89Valv22sir85dK+U
ahZS5abn61XhfdHKY4d5oRgmunJAmMVmtE4kkYawwvP+gvR/OdBl/sWu4KwZ5lmT
e/FA/U7mjBLb1MFNo24j9/xduDOM/+zpF8ZRYxTWSQqU4bT1gwaIhlzaTW7HpTq+
5VaK5u+IASylYtrC7XH0IYuLYulHPn2N1OArVm7xxDMyd9TmbEoAUMLpJiS0NQD1
TBQPYUedV5De/QkvH+Bj/M6BOcyhhVrF2TCiIH9a9uSKOReVXHAdwJxBHCX4m4fH
mK49fbIZJQ2Q/iXxJUvovD6kvlz37RVHtFnahNq2/cJ5xMj9K35rCgAmSFj9YK6h
mCY3O7lxSA0pnPU83NMPyf+rzDuJez3gyb/gBCd7XDE8SjgyFKgZNawjw+9267T4
B5tsQ0EYrCjEcMO9pZbJn6NEu0TcXLSsS2HDJ/ILgr79Q82kO39h+m86vcnlsJM6
V1RngYkewyQQwDbQIA4pBy+8EM1IAWkjL17f13nJUhAziGZjac4HBQT3FoF8ieAD
9ZCDIRKCeRuSVtXdkByhstpjlQ9ZYVtXLHyoDXMIZlDkkwJyEeWIGs3iMENJs6KO
NTMIyqB7bp814F70I9Ma0sEcapUauofmwYrczf8wWjg4COuR5sP9Kbma59YBxjZI
/JJbt6EDjFsIqBAtk39zkLpaHhELlpclIwghbB8YQa4zo0SFiIV+NkbtePb1OpNV
004v0Wp59GWGZm2RhDmqJkJ0qVqXFMdqOFKs1GM/ujLw5AFSGC+UwtzOcsozuSwP
Pc2IozMPRrXv+L1Vq9p+3Iunf/C6FXhI+42Ha9YJGtuJibacqSY+t02raMt07p0t
VR1Ax5yvXKUgETHgjcdQaV/6RK8ogiKlYJWmAQRXxZKQRV8EwtNvBUptop+GfmM9
GzvlZGFNgXjwAF65sQQ8L3GvvZ2A4IVC7CHqopS73Z7ioiI7GWHx87Gs+TPgjhqb
skLC9+5LEjvZGZQelvVsaa2gmraNBVzJmtdhi+hdUWnFlFpLge2Rb/qRuTDjvifu
1pGnWKysdTmrtuj5uxgiBQZySaGy1dYCROzYS+LaaxwTNb4fiFlNlI2UVlp1NcMw
wMqkqbvQvqGXPNB36rQOEQwG1j716W+HYE02/CcPvqVUOJKP3Vf7NshiDoj8wxDN
zTQadpzwds5vcLH/3AGGA9mmCTs8efrclTvBc1pP0jjexA1k4SLR2X/NLz5MFUu7
Hvg/QAKgyuD4//6l99GzNhMKlkFVWFyDAixaHOJV8FgU+/CSQAbfx/z4fBz1LCSY
DcK2xcjg9jTna6ibd5tph3wDbdw8qqiM+WlFpLQWEVcR8k1rQmNd3lQPXfvZ34hS
k2RH+LhgKidkJc3IbbYVxFzNkZdD84iSLKbLQJrjDrasyaT+E3kfalEHTN5At7MA
eVaXd/hpnZGQPTe+J4luCvPip9u/9l1VU8x0aA/dZk48WAFdlD5cLtYFmlREZt01
aT6wLDfl3nHdrU+mKOk6VxGu10Qah79inqyuYYRK2ZReSMSgSXbZLHJZsZRlLtQk
dYdIoItfCp/VFQRedCN0ecfqSGpxK8hyw9FdURbxHg5Zw++YfQjPWk8Pc9ljoTb/
5nILtqqrlAl6GEJn8ZGp1nrRSdrTl1PKf9EZR3C35l5gX0Tewfeziqk9jXjMnTE5
PZrTl69JkkzIeuwQPwqZWKfidcTK+sts+gF2xB5JEnbxucTK60Bbt09eQus9PVYC
9Zef1K1jYqxAb8DHnBMZ6Ifj3NB4ol+nwsYkQZJJvEhd2MVK4S7CPyZcY+i3FYZD
u6XMwwIZBIU/VsNhCEio3ekd0hDRWRiidb0rBStQas5B58hTvS3UDK53uagb1Egl
oRSMAtWigcJw1d6BLz54PEUHsVB/fSdyeDS6XJK1i4wlzaweT4rU8j9PDX7D3LBq
yY05U0tXtkVMFvmI1BOWuSy2mlkcn/HYOlYgzfxZHzAe9v4T9lwI4mKdjV57qTIH
Jtq+GlMiL+eJkWDyZ1Osl/MTG+u2kAYl4lQVvTLRChkNUNYk6d43qTUgVtaI+Lan
KRpwvuAzjRnDPdZ5VAqrynLl/XvKC0Hv10cd2tXLSiB3geYrVPsXdX3gUtV8uoyB
hdaOzfq9A1HKZ7U7MfgYxiI15dIB53f2sCFUxzto0I6MjwywkLqJzm+8u3TLiR2O
+yFOT+uz1cxMMmC0GVto5yxvIzf/aMJpcVcBcaV6f3syG39gOhoEfST8RW/NmyP6
pslmAZkFuyT3wM8Bc6RO1XSwAxB5SkllXk/EKxPjrcVNivfYgp4/P2l1LI8LrTcT
ytbwJ0S04yaKeoRvoLxpdX65dQXReAmkK4V4oB2cnt9A6lGyETu6AYhnKYh9hiUC
h2WuaaZaGdFubE3Hz3GsyVR+Rm/owAPADIRJ3Iu/lsRbn6C98ETVJJUbsIef4R4n
LkoR1mGcFbN82zlFeUULjm2yFCjaHYyQI5iLVi+1x6ChFO2bjD2n9K2W0Ln4qjG1
+RfqMBeQTyM3LABNy6CGBw4bBupqqCztV7otirxBtbE1nt8i0rVayl83nGNY+6Or
cYVlOCPTCiKg176CtW328zZWuf6+bL6Mh2qBM9TG950oy7cECc8wTddM78lEzoLM
ceA9rdgXXPDbyX8hHWUER1vQpuQIrJhDO195sPsnwEFPXgVyM2FF5+3e49J6jren
6BnaVL5iPb1ndVXaLX6K0zotgbfc4PU3mngi9wbw0zEZSKGkt3OfkaUNhNpxZBnI
4EO8xCddOkK9b2euPeiCjKdYjXiUT9JcAWF3SCZJi2mbm9X5TFiFyAW9wBOrnLy8
n77ZsbAydQwJ7JBMQsWrQdW6Fp6u50qL565vgKUF1B9ehdCOOr9VYmibiFtuFnVa
PwJ6j9pmpQcfWMn4af6Qch63NcN0eg8rrz5c3n/Nes9MqeVXwxlK/FJB4PIJid7Q
8HdeioDVK7RG8puz2+1URKwrAZ2HnH/noJJRYJlV4O9E1vSVAaZwmrp4qAwVr4Mz
yAykbaU5nmtcpc0u1rmbew==
`pragma protect end_protected
