// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
KpxU5cro1m3mzGn8oI6gtMjaiMc9igeeqUYKWGBiKlXWFXROvGmfbQluBgur8sAwyLyb1Rf87vAB
BUuzmF3rxvtv/R52DBBjqh9o1v78vSFiJnpNI6iupNHwGZOsgI1x42I+/j7Z2cP3Ril+JiyBAeKg
jWuwrhhxyz6D7SY97f7i84PblSyiVgEOhmTqFpSb9E/tZ1nFn/MfszuUiZCywVAnHQJyKvyrmTSo
euPtQHbqyugcidj2y6HVOmvWZQtFa8Wc9oS2dz/kxYo42LWOWplqwZVOF5ygu7cvSobheqeHta48
nqHp9w12RIRqMg8hcL0dtRpIErKUXtnidFamAg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 214448)
GB0+dvEqGs9fm/VwPlkAGTzPDurY9k+VqUEHPDypoYWX2oJqDubkZDRUtKMskjokfNkWm9qRX6Jm
ygW8zJkLR6lhC4AClM/7NfkoaPeeLPtV72+0yny/Lhh0moaWI9f72DxCZ7njJTjFBIIttp13JqxB
2ifyJ80dFgQf4UFQsh+lyhwH9jZCP2gTmY4cu+xsR/MKCiqaaltOR7JJgEPMprXkW5Xiyr+pZro/
y9vVZla065J9MENO9ESvdT07taLYe+t0PJ6SKsFONCyHHmVzdT+Cqf7Cb9XtNVYisoricej4yISu
S7Jc/pe0MWjJjZ2YGYHypFwCYIB6qpDHYo5i1o8/prVzOk5/msSZSmo830xqkpNabgp+L1ZBNAeO
XoSDNir/f9sREy1KBHqmjlV7XPa9ooljTovDcdTkYQnZIeJ6yL4MvSR3ghefS9S4Dg9xfkUmBZ2P
RUzhXF26Feu5YMCGFm49/oVnd4xF9ex1PZA5pg793etZqtQ/sBsYwuqyVL5Kyq9492U00MOQI3AW
qd2rMVCz5hK8ZOmMYLP5OicBAxVGZvU5eqCY/+QGNm6RLv4i+idFmirmEltjRAtX6+Sx1Y/ci+H7
t+oZhJhCNkg4JjrxoHc/S+a7TLeXEfD4FbT68GFsxD91SMdLnp+aP55cA93Xvygd5TVDEAZEn5Yb
aZn2R68BdZSNhztP2nyvGWzBY47GbtkDpPDIlWzHWTP4xHsN72JPI6+ckt0s8H9beRiouI1A75GN
/IWCo7Cj1HRURZRnAkpf1PCTbXnuzqdVrUAfm3aeGIbHJYI6M7VZA6u86GuOr8TtrrCo8OIVbqTs
deXs6wx7bHTz5I/ZAixCXtJqhMr0NTaN7uE50KPfeYepk1PHQ7YOahTyeaL1UO+65K0FbRUtCOsn
Ww0/KZoyv62g48TDZGwics0z1KaYRP41v0vANyUOru77NqCvxApCCYoNpCm4fFUSpGZVRkpaiU3N
DY1tcTVnQUQW16G0csQCHbjwQc2fSL/lB1uT/sl/ymA+qaxNuvBAu6/MwBO17l8dkghgGGd6IfLQ
4mDgp835culR2qjYP37prL6cpAG3Bb+4t6X4lxS5I9zDpGvqsq9aOycWC6isoTwAkhMMBF5Sm9xa
c96YA9Bp7+rhJIsTZ6GCQ1I9WS9GBzUMy3muF7AvRJsH8P9TB51P2qR/2nQ8XYeChOFjSaPgJ9Qy
s8fvGC77JZTlVrjEL0CHQ3xG3eVVZXoOpSdrhOCXjnujit3WMDyn4PoFzCMqQ4FuG+XqRebxKPGB
GJahKbrwRiN+d+CdsiZOZDcyiTDhfAcVX57BnD0Dq3FgJAbCqWvU7OJK4Bzxj000pD5JWhy1V0Mv
iHD0nE68otTP2tgoR3BcoRiFVQXfUw9Vq2T3FGRkp7vVNmpFqsBnVvdp8t6zVYXyqqCMHREK3yjj
jyfNsiOYN9hAqdGlM09+JuLB1oy6Dr2hLD10RZVHSS9qu3fjEGjMs2urDpDsV5QIdPqOGIg50GRd
KchmjzKch4NvcYppPLJ+79teHCeu/sGqIGHt6Jlnr6cgBZJsl+y5Z0m1hj9IR/MxsDajbJcO96so
IqVlCB1dlCsKWVt8xvT/B6LC/xbDud+sgce8DF+BJw8O1bfdGXaLc5pTiDAnDwsYTPGqdfh7P54q
QQwjkDSYfdcCdZvSw2bFOu6dmKqeZ4PIQhLtk5Gwy+HEGv/+oEe7oxbWYCp6u8olHvIL9W9j8UMP
Qou5qqivsn+RwRvPs+Mxbbky9V2wzDm9XedHAxcC1cqef/GzfjZMF/rkWiZP+e96MbzjgODDH+0T
PhDBkGcbKMjFzTXC4UUdP3ki+k5waW+z+q/vXdunvgRo9Ntne/INKXmxthGarVRVg42glqbRe2Wm
qBEc2KH9rVcyNzGHW8Zc1TNOVHH1BzhhOTPMUxINnjzmv3gGblJVf4VFY17iirD7IirT69SlkrUr
5ZwaPIqR6wu215Dsy0659XyfPeMPU13lvipv8/3f5WeDejCTXXBZrZfqWdg1LQ1+53X5AnJBdyWB
4Iyo7yJrpY3993xT08XN0nYOSrDrSmvUqaWSOion0tpo+X/fmGxQNS1O6RBunzmCo19/znX8TXK8
fANrACZbzB42d921D9IG+FKIhor7N/LjXKPnLbZFZHaqgiYtJnZ8dG+PNKjBibHw3FYi3r5+GnXc
xAHL5rGBctYBV8/lC182EplRAc7L0KZjrh3Sm6OYCvyyATIwwSfMUD3aGMbKgC+monMHpZBij0Qd
T7ClU3urIlkjJ82eEt9SDW14sVYlqWomA7wdFKfVoflli480D9m1Vsa1ymvwif5u1qnbGib8uqWO
BTFeWUO9oBYZvhXaXyMS0EHFqgWyffs/tRRpbRTE3J+zQ+OFvgW+Aptt89ZiGL9JFCoSqXSl07Gm
GpqCPxiaD/NPCVLg9sUh7cQNqcExjfMCvAmkeOJtQnC0cI3FqEHiBCG8VasKIh77Bsdt4HBdVfiP
ZImTmUmGLEpF/43iQr7BenLHh14hmw4F6YoUXPhtVSV/FQkalcjT44u2wZ6VyJt0n4UzvWunAWv7
9P98Y5a37WzeYMBgCWTJgcKJIgiFHkZKei9VbJtHZlBvlgXc/nYSB9Dy2D2UZSdgRH1MK1J0lNTQ
A6j3WmNCIK3o4psDRguM/ka8X2wV4SAR4gCb8DVmTmXURYqA9bg6qhSSVpqkETVunKpIA/FXk0kn
m1FxijPi3GIbg6zaHeIVIFA/1JI9RmLlL40fBF/Xchu9Yfl+jBohvqccMQsACmQxwoOC7wzdFkoH
UgNNYZbUHDi89LN08Hy/Z8Os3wwPn8Eyp+8GGIfqA6H55jaXr9Ib+P12unTgGaimhYPq6MTiU7SZ
LOl7tLSMoEEMbdJknsKazy7+t2U62pRlcuN3AK6/yVisTxyRE+lEcRaKFaW095G1/BpWuvosWrzI
gJXQapnoYS7pzqECjIhk6BSVkI4oxvXvrbg+irP+iSjE0FBpfVhZoaeOZDrn2adVLErinNEerpPX
mZ2EGTgKTwvkvYaVzAz0rpWtXxlcVX26/42VyG8pLjfC+icE918Zt9IKNXszHAfMGD0vc0JDV2uN
iTtuLYWXXQWTxWY5C8GINx0c/JboxQTdtRM3zIA2E3HfZMuorhf7uHbcLiN3+zzpAVB4gGxe/esx
co76gnaO0k6yNSU4CFEIfSoRyhyvES7O4vF2BEAX4/Lr8V3tpK46fq62nQPEM95Ib0E793tgaZ5k
ND5OY9jzV2gW5GzqH7SrJzfTGfNKs9BHpbYpbMm3goY55OXk1rC3ZnboZW95nwOvbdQDK2Gg/0m3
vfxnloUc+CtQIkejuY+4Dl/8Kv465tsEMZ52LjP8hGeu2WtreSCuvT2IZRgXJBHnT16xkR5dvQ9Y
JJBvONbCqgXwQEPV4SUg450wqm+Z+wKQB9qWbwtYL6ni2PzYebob0IGLH0XwkReRHWy/jzv0FD1k
uqMeSGI+fi41CI7UGGPm9VkzCqpqlBnLkTtP97b6UcdqC42+1c5X5GXFWHhkjITVwOvY84Z9qJby
Zsrnggh0UlK9vrw3q0rABmafT11cgF/zLB8tzMk/f+1S8uSAfSyK4zei4RAe2GoouksUAvksPVTc
HrSFvW1rsIuu1FNCa1OOd0Ob6JeCT1oMAiJgQDFUNpu59MeP4zerremjzgiX6NsfcUjJ4tvKIWkj
o1y22rTnVSlk6nU/wfCNe+By1ZuUcApATFYrgz2LToG8nUtI3ik90BmmVXBgYUXKsVM2Wp6WW68d
iEIFSgN3g93QWS+XAD/w6JC7igZ6slbbReb6fQ2bpiS0AibPDcU1GdpntImL0qmFVk4kQh7gs6ak
J88Uo1vrybNhbSUqpcX1GejcSPi4hA+08pvIgsze5MqjkPJvsy6yGhd1Kw5bxh+Ev87ghR8C+gvw
BSPcH70OJRTImEbF8GUoK/l1w4AcloRaTwOXRdmMNN32x5/S1lqt8UuBdwUtjp66szE9OVKBjJNl
EK5PHopd8y6wZBTHJayFb5tRR9J/1gbEua+lzgSP6RFJrOgsjxcJRQ22d9eJqqmXMY6Ul8m7iAiM
C8xo0n2YGz8DJExR4RF9KqRUnGv11+/vzf0MIqI/6Hu+o+MGNhC8hQuB2EF25PW0jPEyf32ZpimV
oaRXx+ip8lwtRAdLTJ3PAU8KcTFxSkIhQD2HX3+OmzswsJxFnyuD1l+jBSoIvDp0s+B7iYQIXI7x
WAvk6xNdli/FthYADaeQ9Yscw6bSIBY+zCth4paYfJ3MFjw/iMe8L/sdxleQ1jWsJQ7lt74oEeuB
sAvHsK3MxuUmw4oJdCPp9YK8aV4RfmCeUImAZAknN5ZaW2SPUP5gweTwXJVGdS4ftxUrQBD7k0F6
+xFxvX/Xfo09McQAvNItNBJ4O9Whz89SX46aIvfHpWM0Qw2++a8Du+Y53K4AhSIkzOq1KyCdfYFN
PhdmRLLnX5mbBCXyV+QQ0Gn+upI80jm+QYakZkGdylorMiG+vf+h6X4Fchfj6QbcZpt6WiMr2nya
zaPw59zXDfSaFePvlMsYrQXvyTS8ExyPK9NOZixWlnk0JOghjKDcbgyqzee+Xhq81WfRfNoupJzv
4l2rB/8sWF1F5S9qrlssIBMpROrQn/bOfU8osKFxHtbPBwbQJ9pLFIS+x2pGZ3g+4YK+oop8cBoI
U1ju9IGSLXgAkXZ5p8Diz2z371mRwUDlzKDI+Sg39Ai5ZLUfslhWqzaE/iKBpkbdX5OCtzDmwjmP
Yr3Xd68+QbAT1cH5Spbf9kS+RmxirTxjUD8i0gSTTdcuV+GWgutyNRi/Q+n3R/F75PGFj0UlkRND
zcbA1hXsrP9skWdmvFNOPjHDC1i0oU0876oVRhr7v6T9BZfHyVZrQXVCfYf1/1Y8gfXUbsK0LeP6
4xioeiS8K5x5mqZAXohqxQrsK1YoOBGUd3Ln6G/MDGsBvZ7Ukz0nBh90aGCe1oZJ/HVX7MQah5dQ
UWLNYzJwc3oV6UKHtgFnQ0m1CbPgSQ4cyTltoTh+W7/u1j+UgxIRezH/mU6UMjCdAr5T3tpTcRHj
rzO3Z5RNXh8y3gHbkRlfLc5cepsTHhHZbWJv4dJSs53V5TEPr5JvjfF9tcobztwH2Q+CdCP6H04u
/ro/NdZoqDe+yUHqS4jNWLuGLhswxexnIq5qCTxUvCX4P52ZF25T494oxdjJdxdc0UMedmQTEicb
LlAY5n+4QsckFpHz/zGqIfZtR4th+Ug4oLGDBuSxl2fBXYIA6yBRfOgoNxqajZMPW6KZBeCD0fF7
VqCrj/LKyYgWeACa40AQCqJdLtz792EW7ud51NtZpbyeoVvtGaJ8Us/v9T/0ysq5tYH0ZZN+bQum
yuaLfEXT79EAh4KngBJu5fgngTgPGG2VEJQi+Yx9KYMGg5E3W0WnQaZv3+YQKBNv1rcbB2iJrtsK
qSW11yWD9HJ0v9KF6sAqxlJ8NBDByv+Ic6K6n43lFU5Ktc4J98dihhET1Fm5BLwynNVsNB/XjEfF
IujUMpvNRtohkDQ5a10rAmGvvz1DBOdw+kOFNnPg6ytXjOZ/bWVw+x2x4DolpWnzaYBeeJZltjf1
PPGyyVOVTZen+1dmEE6zprsb264BV8M1L91g9lmJkkxrHEfKvnDMO56lYMV+mOpmtO9WV5yllA9Q
Q3iOMA1269IPsAIxPv0JvbvBtJ+Q7Zef06OG0Qlm8/0TttpAogXgYngIVHXrDK6G7qbOZfCCzh3n
rx43gc0PhRWwLPjw4A6HwIkFHWMc9PRJfyzEdoA0uJF9+kU3NA2628f4pyzaHCzwfkHcyE5F5unV
MHsrRfRcDNvBbXdALRtCvHfEA2Y5Ex9P5VjbU1jvRFKbxnmFvy1+6J3ukPIEv3tmfVIaYPl+38sy
uPjTwTc15FhULnd3x6nx0M4bM3IZnemlf5H7edjR1KGfuofWtKAyistIPIIsHnPFWG1ZvmfLacSp
GtyaPPA3vSaDqmTfHuNZsCtjB7F5M8hZexETcyzi7j6gjM2wSca4EB+vP6Z2QzFr7EoeqPkMg92r
p3c/iEI4vAQS9LWd/FYGq5Wncl2RMAtXCqY7ATv39yXQvrDyzI1e6wLYnybY+Yr7kl/ml/3/Zmwd
PwD0hOp51I0Pr879dujaDTuNLN6x8S/+xw+OwGsb3j/8Ob4wt6fGRpk1IqdQg5fcCcyydwsLF4s9
XRvsQUbjyaTI7n6zl/QN57ggTOzcnIhUE0f5J7h2Cw5oIpbw2WJXPp6hsyCryOF3V4KRSs/A7drF
uF2KUxIuiOhF/fF5UO7K3Qwu2XZXAisbHptcV5WV0NNX9xmwwJP1gmCBlX+5cU0jrppfZLg/QY3V
esXLqPEpXp3zBhj4+rrQ4dJE51yJh8WLlpu6o6al93rsWSI1WG+VNRyzjESMxEj8Pr5p2vwExNgY
8qr8bHY3CK6iCA3VIlQcDTeGdnLiFvsGMjn9AX1UlN8soC1d264xXeMikNKNX8kdUTOO7Me9wtVa
xw3mDVNKDRVotnRSrYzsrMLU3Ie6DjCjUQKGVvk2BwtVsntUFuUFS5/nRfqnQFoW32a2gFMrVb/Y
H2WFbRfz8wbBD6/jqnavcpv3ZyNp9WWNfetbCta/E3bHb4NX9QKc5y7qQcYievvOzCJRDbIYENVu
JgnJ5YeeefRGZN94v5mSraH3rs/2cJ1heJalG2LUZgx3jUqtEOPr2hvbgGGAkA1KPSxzhoaBOK42
SReQ80H3R5f4poR6TSfRoQVHC66rAZOH9ZD26OlOjt2G9E+qwmhHaM0BfcYkhuGbEPSfocjQFLrM
MBYZfgHFYqiKbOG0sV2aBEv+0Nt/4x0CSBfmH81BNA1wABrZywbK366dswhJhiXhtCettyuPF+iQ
zGN3UVCfRq/DuLQTSqxqveW2+AG1wd+1mF4FxKC493VQ4Axqtr+p582IFe+QtsJSda+47I1oCOQ2
jpdoOJXfNqdw1esHxCeky85ESO9OeCVUAn+ZBW69p8TPxmtLRXo/xWbiZ6jMcMhLWOTjYlAUz86b
m7DG55TjFVJe0pQKcYFhpDmDaP0ACrHfofmL8HbyWA9nEqyyrvuE82I8XIL/+U0n0b6GvWyOd/rE
PmP1ZN8UPK4j/bl1MQYyKStqE+JoHv0lmJuW+avErD8WSmcDGaMSpylKmF+yz2OiUBA3Jt3JcRbs
GK8/0bP3Shi4cE+hnvE9iLToq6pXc4H3aZ+OHiCv7DGg4wIeVKAL/MbFEUJ7uG5XUB6+tFtZcVd/
g8VCYgnl5EtUtk2AFVk84PEGnWtIhzBK3/efG/4dKjETCNFH8JiRbUZxO4HBcLuzj/ZYG34pdBK8
n1nUYBatzSXEhoG2aQ6pfr35aNnVAzE8OVXpoN90TF6qbEq3TqColSNTsDMBqr5bR+Z5H2fctDB9
52SdNqINeMRu+wd1mWEfUqUtpMlvBpY/mqEI3sEMo+GFcuSh/hIJtcoUFhvlMFsi25Y1PQr08ydp
PcteakHCr4FKm/E6eHvz57p7gzbQKYeuISWi8uip8hvCMywJP2fNCfScOr2eOW9tOuD5VcbQ2cs0
Zdrnk+L7HUdUy73OwBb5Xf28y/fXACyhUoe5g9jmOOX6DH+zJMsDQrMqPSkVzJ4yugVF0zy6DBDr
QC4DjwcORBCMid+dx8MQPtBMDMv/WkrNG5ENHU/vXDMmgKe34UQA2ac/GxEYa3bFCtEt68XQElG+
dA7lQSQmYzK4EmtDOPlXc+gIMYGKk33Y3CERtJzQ27HAXpqmoFiSegVxeHdJkqYmjSXrgsGOPmJy
jY/7utbt+wDG96Q6K6RsZ5smDLOqqXzPt9y/D+pAkq9wdZ3Op4SmgSKbsq6x+3mJOBTqN7y8AYX/
eGXqXezdcK96wFsEgFdXgGRFmPzPRuGxjQ1/D+zGpM0e17HvXxV39BDgePRvZsKzh4FIXv59maKk
hhn5UFdKcLSOQjG5d6bG33z8zM3X9Um6IeNBEnuyRXfY0whl2GCbLhQ8251rc9Oa9nmXo6VtJfpS
kXNiVYTWy37lBV62zdvj87m0FvjLnDgkH3AFDMi2kwp5LXYli8nYcP39NhMpMKe+znhFfHRjl+ac
e659MMYRNv6y3s1MpkxazoKESBk03rRtjR/jl9bU3+U3iPgW0rSMLaP7PL/phfcTU9bPCFG0g/Pd
vslHXuzkDmi/gk+ScEGDyXV86SuipF4J1MzQY5HR+3CFGpk0FC/gQ3/nJ03oeRBQ+8pDcmria9wr
ay80I+1Klft1pw2qV9+Swy2BrsaI9UuOdSPeqxOGUMVnBcWwuOcO5yWmW8qCP8Oe8Xmiqo4EfW/r
GCheW9ApoK1fqZpbD1WkHqWOBCJmN7tMYIV0u12DFwUDM7+GHwaL63KvSx//xMN2odWDCQGSd4m4
TdQveb0n5a1BcX6YMIi496E1vvEEIXuUCj5vAWc3IHEaW3B3mNqs5kmY0eUqplUth6IsAE7LMw17
XI0nwgVAPajEeelunE6XZqf0Y2lnnljk0A2ewhOexfihCzsetFQlh/TU6p/u47JgOsC3rQCdHf9b
2O8gvtFQTH2jfT4Hh+oIX6IJBBb8rq35Gj4LJsXdGWcOVl8BtKNnIznEqkqSzEaueVN3wIn3G1yX
Uzq91dCa7JH3G5Gr0RXAbyMUj1i1XyH9F8ckRj/8Hl9+AsYK1pLIuv+4OoJNQk15rykufg2WT1uW
rmP+ELHokFvB4O+aZitEGEvGQPNa15ax+Q062zpF3FMXv8LRueyEkzBJRJD65kU1kacTQRW1vo2n
mivMR3+TDTC4LxrZrb7E9jgpfzle/JkwigIqlrMhDXrfadQ2fa7Z0rvA5RyvVBuAuSxYVuFQdTqD
q3UzdWGSlBhuOd7P9yc4YQDia7CHWo0jJ/wLH/xBky2tpA4qS53XWsIOn7FBjJ4H/DafmP/MYfVs
VyN+obVNfkMc/nhtGT7TRHZccoFBEMe+gVtwg0O2vlnkpInpa8HcdKovflIyn4lRCzpJ7uGz+9li
E5n2cuJKKt3qOtdkpHqVSY3uY5lJsDUiP5Fi0/+qx3A2wn9iEjZnBgUrRTGo6yWXTIPFGoSmiCL2
g1gBkqQIWpO+OnECH9/6EU2lXHJDi9aQF/XzLNIhvTt9tAK+3qKp3rm4bJcK1LTxF9wXRdS+ajF7
45S/w2VpYY55nKyDVSiBX2kqYvKadXXrVFcjT4wNZtKx35nESsSIrnJO4iFh0YRBh1iQXv5MB8P2
DpxcuzdzHW5gA0BF2nAVcLWXRMpYfsNWYau4b5GVp6UDNJNmZ9HJbv+bd8I7Cz/ZtTCWz3tPEfx5
6yFfSYdVYX5/k60wCd77Tw7G+Agv2iK0mCkS+eEUAqz6Z1/LoXH78z/DqFvlc1xDWyDWXSZhaM+w
MZpKlkoKbxsBV8k6c3JqPqyocbmBYCXscem+yA99XDu3SFhNbwVvXPLfpFFBRt5Fdeyh28od0lgh
gQa6w0njLt81j/Ym2Y3GFRwtxg87MXao8EjSgFQVvJ0ODqdo2SgvQKzY4U59sv4DbhyqsAnNVzem
0yJf3eh3J8lHLmPTSCcJl698K7NWVc0IS9wiFhJgy2qod2mfvIXS6NkmE9qnkFgI1ynkKAQ4woJQ
cP1js5RKTMQHjHAdYMklHDe2eiKzHm0rvH45slfKmD37DG6ASZrg8c13eyR2iZViy4uZrMdNdBkp
GTWgZ0mkfeazwaYYhZ8/qUhMA3fnHmJXnsg+ECdZTpsQNK+E8E8WhJGLgRgDSOaWr+RzACnJ7ShR
YmDnFdpAJ2eBT1g1COOuUHjqkAcs1O5XnrXlJkmIF4vuGMpCjNATE+gOMbFvotE3Nox6KLHYMAtS
w2AXsKuxLVsgi3wSCIKLFFgC4K8bxCWcMhYFKg2vPlAOFViAJiyEQMSLYCs7ecyPAXbDF1glY9hW
sB84fG1VwMCtgMCg8LzRFL+mBsQ7hlFQhej0PVqwhGWmEmURFsf7CvySOmCcpt6PYhh98T4VO9RN
0CRm9oPUcmjYwb6GwgjefBTfrAtuBe1S4YEy4KL2hr4ft85yLoWVgIB8bZLNpkwrdC7jTgbCYxNa
Slia14MSgUvWMAC62NTt7VC6t7n9PnX1XNvaS8UTNvNiQeHGRZ1XZP/A3QbJpn4v2nX6iWplPlMA
POfrmQkXy4XxamJFCdVPNbhZoABqGkiKbJ50Et/uRasFNzEuSzfGUVWg0eF+Ggo0DwmV7KQZHqqF
vuQYdlg3scWSOxMltI+TcSL0TbbQ5CQeOyqAjMrwfl6QTYtcU3k0ROIRgj718oTnzWB/7Z+NQ7I1
aL/U7HgYukfOYIcyP0TY1eSxGroq+//VV0+eTVnG5cJwfCCtTySCFJnMKaw9PTQyAmNircs33rte
kU7g0LtObv3UBqL5wlJmLiQHxbaeFSgO3JEy/nOEDyqM4xvm5UZEnllbSKzzTOdSKKloC9F9vSlc
b54i+URW80Cr2qlUgDMacVNJSPEUrejXt7IzRlD57VWegYOWLG5TwGKe7YoMuR+DY3hIpU4K6E/A
cqTAUL5HiENhb6RPZs5QAknEYVCIEEvIJX3xXgiAJSKaeM20ZazFcfSQypg+FiLBiZG5Ssi48g1i
kHR7FpLdVPYmgL4MVZWjPrNsFn/ik6wiWs4hDd2i0t7u8/eEskXXs026UPsgQcqzKQiMQbfTRAfC
6GvCiiMXN9gSMaYjU9j/LTfRKaxT6Rnl98g1f7W5+6M88XYAkkzvHbrba9zCljhLc137AZDpMTpM
bO7klXxy4pDrZ+W9Xn/LdsBig2oqbyFcE94z+yX9rTVnNKJNJqJZcxWMxAD4QYaibyx5KH8PaieK
q8wihezm+G4s/COhwTUPhHCWK4LlcY0m+X84QMutx25RziVWT6bhLTfnZESzm+daGSsLCjcTtHSq
44DjQWCppQreBh65QU6UhM5P1uZFWdvH9Be2EmEx0jTq7t/rAOAc81cEoliYgtWVjgVHFXEm231D
QNLJprP3592BeHK+XpEILmLTWK6hxZYZr1vav2WTW7mUbVFtwsFaFaSLoqwZloQiD8qRBLSvIk+9
omThAu3eBnUu3cMgNSqF6VZPDTF4Qw40RGyCmZ8Qz++pVTeZH203s2QCjqnznnzoTCCwt4NbRgYd
XeyPhM9wxoFODWeozF0CH9k65ZSqEwyx99eD+0pBc0P1W51ajRulsZGNuYFwRDQYXq3cbsLurq1s
no2wYiLU/Bch4/gmYKibGFwf+3YwQdne+daGFls3JMjxKnacT4OVB3dxVL7kOZZw+eyrT7KCp1cA
GKfjY/wGv7D/LFqgapYHUI/532n4kzxLsVuQksYglN8hKzqjYF13J5Su2WtMFXSqZAAS389lqNmg
cmlWtDwGu7DGpc0U7NMvGtmG+rsJ4Cn7X2lDizp0UZKiH0/w7JXQExRfNKcOvbQEWRt3F7+BcGj+
CTWm2RiSusN7t1y0frd4b6DurStFwgNvJFovU/H9fFutzEi4nMqKCaUdY69Xb0JlIb/biCehKs13
euZ068Z1k5nLapeEe5eLzyxiiqIbIPZrk6ysXuBA78KUc5ltBbTUfUXfkZd2ML+FFnScoeBCXhpr
xgrDKugkKHXJOpVWblmUFOoOrDsp4ID3kXl8VFB1O6BWASowmNYqUQerlzxhaSY5cFlgRSKRPcn1
wnedmiq/6Ue9MK4IncBjfrY0p6NSbDYnmqI82TC2nu5ZQBky/+b5cc1xAUTsfZeLAWOvseqHIfMj
0v35w2W++5XHRnxkfhMsEMhRGat622Rya/55ZCSFDJvH5LqHF1sftmS4dZQoYRINiEtCfQqzCJ4c
Fq5uzAMcJtixtwLx4AnZ7MBTiVM82eVIGQx9vlAxNRA4JDTiObqqs6AAm9U6Ib4L3Zn9fUd5pxkg
aXX3iMKfrSxZ+nJqJzctGyrvmAKhNymboEiRAUkw83xLHhZhwdzeFiBYegiYr31RAgyUS6j4Prjy
3pYxiCUoy9BKCtJMsbhxpuVoa+o8ajFX7c7dGsXCYmHNn7rv+oWm4SV3fTwRVnkqOtJRmzVdxv/B
Zmk9uAN90ZrGvoXpMU0+/ZzLRd+6dTk+XdhAuLfSSA4crlsjGhy08wbrSJN3boquUjKwT612jhPH
qr1eCPsnQyUTIxLWUmmH8MIO3hzPUctKeFtyq31/8eIBC2uslVvdBpQEQFPoHbvDcDKefO8yPMiY
kfvC0OSlaqHBXzmEX4bRC9bUkpPNZLnX3uwQ/52JH3I9ShT0s/ngOO1bS3WkcPfNeeSON4BfNCgM
kg1PfBEqZbCCF229zIirVaEGLqa5NgGrZxFeaHqRTWqpOBA3VBAXDl1stUXnYOxCJ4fj3kG6sLyO
/f8XshAZ4sppL1+tU6qQUKCt2xazcalFbHh3BZ68johzTTaoGfYhcIJwmGYW9Xqb79a/gWUxyihe
TVyM669CIQOiQ60RDdr/c/i4O9BO8bsm6d4H9p/wf+X4mPRNIB3wtD1Re4EOapzuOJKNd4DglQbA
qKLCwxZVdd5/dsCcNmG5hN7tWb61gJLjHp7fEK1xXjQL/RDmdRzg103f77lDfrtWR3s8B3C3tiE0
ps2w7ZeeaVdn3u5yag7K3MiW6TpI0wk/Olm7XLawyRygdMGRU6PLG8DJAIUe/yPLPMTnmaCZKCME
Jcx8Amm4d5+CarMDcpBG3vn+U10RFhvZ8U0jujsAqKMgsBkFGFfW3aZZep1gjY2i3YQBCtE8GG3W
uDFqXUVmJtyXik6RnKLC++mCbSUyGcXMMhuutkUo+Bw5+poShhuvjf1hp2qEO8Pbey2m7YhGDKVZ
qtbvCDPig3rVhXRcIasBp8fTO6Lgq73OLJO15OEV3sFLOjuK5czcb9j9JdjajAJl1VS9W+VNCcPa
f3ABCtGuJxpLEBxWzbYNkdWcm7U7uYY1TviOFpsr2f2DLi7XUYSgoiNT8zqkxmHnamglBPuM8dKR
UtxuFsC//yHv3TspyRa/lB2eHGT6nAqe1sBC+KgKgr4RvmYS/2RXuhfWaxPb2ujSNvpRpSYN1GLe
wbHVHCg822PrQP2VIlJzA3EDQC0bprMwmYa2Mjga/9WzD4W8qL9Nfo5V18iqPxpHX/kNe4JOQPcN
RMTM2TH7IceHmP4XGBZa7aRUNwuxFEY4cnP/umxwfwnT1+8LTnRQNtQ+da7wFCkKmC0/liJID35R
VbWc5TOYxIkOuaEo1tKTO7eqnh7uKgCg7QlpIinhQo42n4K3wfeuhFtiQsikydVo5Uam4rpeXRHU
Rv3/uNMIwM80zrPdbIVSlVYrxgshbYUFcQPOO57kq+ZU1yUn6kHv6jnV7V99ru+ig8gqXi34FdH3
jLLnynY23NmGpbKcGRw0ooVr1Q2qi5NiOg+15tgEfWxZU/MCcxMiaN9kTQFz0brSzDEcCmW2eD8s
EoMFWNLWF9gKriE/4TtHvFJ660F1HLHHP5mCTMoi2bo4v03VTY4G8J+8s73jMk7TDQ8j/dRF/3gH
BuuQMRSfM/odCYUIbe/DP4hGRjNhsIPx2YUx0Ox0lK4YnNJGRSDLQryU2SYEtd60IATvy8iZVzd+
VmnQuP0CSY0Wgw/Ac+J68+RbsR0pwcz6t8Q6BQDMS/PiBGKKH7Ml0oXPqzhb0jBWGfpR6dgg3Gn6
4Wg9fNyyWagl4jpBvtNrzk11afZUX6zHQB04/5r8ke4dZPq94rPdgtAIsAeOUjpjW5O/Q4vrw65/
qxlcAh6bGFsx3peq/YFgRO1u5/Xz2tr1xwyJ1OHqX3mjaUAH7GAod2iQOkexUNSZTMus9owRTovi
DQrahM2CkH3Iwx9e4badTF8vgD5Ogn44bTUhPhtzBo9jVBuJOyDEwRerDO7US4IRJeJWvNqGOtzV
++qrQwYFfiJ5Gtv6JFn2f/hiL67fsl3i+vwupRlYq2dzZ/olQeWzJmPmgfYqJuTDvcEEJ02ADkjF
pFYZIawgevIhmLNhE8mGIvabjV/YVPfkll799zjytyl3pBoJcwv9FhRwuzETtlCmHq7DDIDlGhy4
UASUe5czH7eGDxPgU/f/KWKvWDXewkxROYbQywa0VEMrU0nM0NqiupJhZUoWTXuEk0x/NaJ2QZNi
z+J61mZrMmnGkx31/RNFUQPfSh9OmPrpco5m1+5cSZ9wrA8DA9wdbGJmGSuba9Yaa2b9th9fqqYP
OCWJGYQccoFEqJQD1YyJx3x6e/6S/ho/Ahr3GK2uyOPUWqT11GDav7pMDyPCnvTeuqCNl5aTWFCu
BLi9Nsns2jd4z3hvarU+Zxix5FoHhiKPeq++fO5SB81ySNKGet0sR/Qt3yYIekvn1wi9OsDKKp+Y
Bhp2K1Dkw6wVqNHt6NCW+VTVTCeerxhTQnzVIKR6XaU6OI7PgnDe5oTK4Ejz/xyYVT/gt8B+BGJN
amLRrGzSRTrLjweBPvRoN5D2E9UpACNNcMLHhHd3kSBDrY7VKAi+YqFIniV8T+hOTAP7N6ttFSQd
/PZ1ffDOzFsp7H1UuXkJMHjAUf/54H4rQWHp+lD79rb/37NS6ImMUhbM0WvsdJNUXA+AFy3UjpfY
3gA84ebjobmUzbq4efttQ27uvDACCcyok0dzDxO6dsfaxa1izY/gKCawQrSXEhhj2CJM2+KlW4V3
kWpNqgdjTr1W9FW4lzOLK9j91CWnAeCtHFqIYJ3PyKx6rrRHFIb+hrmnSkpg3A9ki54HiL5vwB+p
jRg1yerh5FkiC5SSU7X+XQBHnuiZnmIrEmD0XhUrVbASudf3oXu4mS2JTEZ/WUbaKvbTvdlaDIwM
2yJ9Sg9+dIXAlA2JIjZ58zd0092Butn4M55WfftAcLDb6aTIKV3xmQz0Ni3NhP+RCITUhvYoN6q5
FqYN8mJcinTixcQYfaMRwJGdbhGpuoPBeYaiTo4DHVJb+rfQnBLSCPiapGKNFsnDmh0K0IwkUmZn
zl1sCIIQxAzgut038uqtFDwaRbGuhdoiJRBrZTtNn1/3T6FHQgTCHEsx++EDA2iw9ab2eTQtwJpx
VtLmv4EpyGk2XruVVuJfnrWyz/fNFWd5dPAjdDxEsTZ9op8nq2fvCbCROovi/DtdTn7mlKkf0+br
vZZZ8p0qybuqlGrbRZAOddxalDhqs4ViQi6ckrRS+7w7xivM+DRSceQFzZL9de8Ch64B00EgGRI/
YhIYzSlXpcMINHvSNh2dxA4MjzOdjCojm5MyhvfYri88DCStmewS0vbGUPErVCs7ETySc1q+qNuI
MkxisRjb0rrXDsQo8ZmO6hxLqGISgJf6mKBgcy693pyMm19DUptMRe9nGOmZkraopiCUXIoF6UIE
U1fWOFWdjTMMBZTY3ePBX3+qFiq14mfAr+kprak8TO9axomCZUeiHmlrbFfS9/0JmrnIqLoqFFjS
Ub2rUCaOEBbz1/c2Zk30jPB8V1xUvXOerw/8P2IwjRGoHJc5OVFXxpP4pt7vgKsEUPiQINujAYgD
V6OtX9ri/u1eJ/d3cqK/SJ6OclF8jI8mhS3E4Cp/ZiSvd0BnL9Tv1sgsV65tHzmjKfOnNKMVlTV1
+/9nGcpmmQUOs3pHfvcSDl1mXu0/XDyuKTFfUcVZ8xE0HmS1eHzBcT065Sxr1FheQqyMV8qH8usJ
wF67dYRDzYtMCfZhg2DLCyQMcv0iiAfXTLpXCb429qCWkWNGZsYrNbpGC9c7K3lPYzaR3EDi/TPd
zAU0/tRE9JtLdNzO4oL8YDUOwscy4LoN0cdiwf95WkWrda3WtIR9Na1xx5Kwyfnn6xbj+pavZvM1
JcO8Qv7Y5AI1t//B1LZ0IVtxeEsLjD5q/7SptYcBsO2pBq5SFtpIGMv96jg7BWHCOtIyxyfil8Pj
UuJ2N4KSsDXvPO/vC7Pq4YbDv6ZVvNDm6Z/tkNUgzUyW+vk7pfGmV+WTLwrioz+hniYu6FM7v+Yo
nFrAXDnlIRhEr4iZ9EWqvAc4qF84327BrtnceFGMnKB8k+vjgOdjEfPxcpO9C0vFMqc1vxAAVupd
cCDOxyF5FrJnWFWmVTwMIC+l3W+BP7ZdMal3DEqF6/Ey9uEI0hOK8jFupXZ1TBWggLUeTeDirD1h
4sFnWW32YTKOAKuMWWcZ8InjJCvNWA7jnK7qEpTy8QTnbloc2OyftpcumF7CKIXLDk+yyIzMKyNo
uaSv/qjVrGB4W3yupXZ1vkhHBifIsAahlzy9jrG5P8xdXs0WjLaelis2bVr3fZSultwn9TvTsSKr
nISV6Ddzbk2vKkpuFQeJ2EG4ndCxvUNQq35+sTBTRYH3KfDIstVGpkqoQnl3403x6l63EWRPRWv6
HohWbmxtInldpsllKs8XPQgW9vObKn1U7TQHY81NA2k4VC0AZWPSxlZHfi2uFiv8jva4FPovrvOI
ZaijM2zxTa4+Ivuvj/gBFkzVz5/l8YadQEOFtuXpXKukQPnt5xpMspw2UeTxA2YX0IJxGekwrpN2
/XGk6uddXKMshmQxgDKOKKd/O2RHBKSOWShSsZRJiYXfsbC4CVKpze2BlBR8Ekh1omADqbIpomDo
lWYE+AzoGl5H6e2eG/uRd4OwxS6gre/mY3q92P30Bcns8S5u97k1t3mdb2vhCbgUJbCTFpJYRO1L
Jept2LoqSfEOeYYEMcs23vKoMPvzqTBshEmUvbDYFAhv6h3K7A9fvT4Or4IDBCVcRhJJhABTnoRz
3/CCQ4vhQ4xz7BaswqVyqwzP7XZAOJ7A5H54bREloaG4ELcF3m/IOKRVjd0UShrjAsX1K96FOBRG
uLwWpA554lAn6tY7Poee0JDLQp4xxAYxp6S2EP+VOu9OuF7Q2vYUEm1iTrpYJCfeh65jSG7VcebZ
IszuuYzRVrTjXFp3FHEijbrzf5VS24IgCdZRbHD7VJO/63fmHLc/+lmoMkaViHcGtiXiWexApik5
RkaS4THYoDUGyFTZhAJ9hEO6I18Lk7r0JNtNDbbKorBFSTys55Pea++0xIPzUuWKG54mhd+gTSOb
K+N3IK6lQtekrs94BmlQwBEuQybcRnd8dLu6NPaBjn3zf2k8m6LLjQ3hxEOUS/Dj/GT6iTYTML0a
VazK8YUqnfzoYfaUxyOZTnruePK/d8W1/LCG2Ve0UXWK3k7WNtt+c6tzn8BDdp2n1F61sEVTQurT
OKcBeWDB6Ap4sJK+5URHXv9WmVNAokKxPBGEsBEyUV5NNysFIZuPmbCrDHdT8MwSq05Mjp2wjVcs
ZiwriF5FhgkiphWsfd38siPfmfSFaGZfiS0+B4n32pvPOisKpD7v6hnPsr7lJMfSdPgkTMemw7bJ
RGRxo8uDwI0WqGI7GAeWjHly65b0zFO5TEiSy0OjLuwAtN0q4APumx22fMKlMYW+insYVbEXdoFK
Wd0rnnYk3er+Isc95YH6CmvQ2ujwQaSYy18P3q5VrmBomSgW96MZgrUrCKswh5XM/cTNFck8bg/F
SMops87F0rcXc2GtHfCHoXCTsl0cI4KfXJurokVp5bSlpQhwATh2PchdFbZH/dKzbQI/o/RbJK6R
UPmPP0pv6wo1EYc6CuHm3JRBqtg1WCwQBOFEXUJfnzWm+PuaGTnxFqZvqYmw2dOHyEn4FX4xTAaM
3UwsLy56kCRi4hM+s6bx/3LM2JlozT3/IV3RvglY/K3fuU2ddV3Yc/tzhQraRVnG0eXWoHQYTwBZ
VQm0737gPjG8ymMFtlXrnTpVBrdMO5reZwWTcVJOuNO/H4A3pX7rVycfpHE0/lOVZkXjGifsOlSn
c3/si8f41mFUp6h+8lJZsAWeIWdnVfxHvKUvszRs29SaQXvFtPPNw9BY5CYzSTMZuLZIpyi9osok
FeYEt5u/VS1Jvijm2EIToDVS8W4BeiXfiBWkPUv8oa3jS0QQNwdiNaLpfr8EFd33Kdyl8uXoj5Dp
ZohkZC85FTw+SsaVYI/xj/mkSJVTC1T3+zElctBu79SVHoAyIxckaJIAZW7TahSYllIcr4O7xCqC
PlpHhRippvcxOxk2PBmvzGI65Qx3akcYAXNX+s9xZ/d3Aezg5sqA5KZCg5tsO8QX2ixyU2w2T9aI
KI2Di8nfG/Fo3b2qdrgOrrJOrHDiJTNJDUvgZt4FQokCKCz9TlS56rxKxMasqd8oaaG8L0eLi3on
viNd2ho28mDFsOIVxzq5/rv8A8EA+L5n5ka3F2mCskBOoa1nPa+I7ScZCYhCdjknSp+zps9uHPF0
hwUtDYYNR4Gqk3C81AxvQQdtQa3GSuwbszuPgD0inOxsNR3ZSsfpUyGrOw1viW0fRQGAjSZX8HGZ
mXV9QNaKrnMA0ngXaBdXk5iinDiqDv+o9LZuFKlCYG9JZp6b3frjEPRGkJ37J3uHK6oYjC7OKae4
/JdYbuzSVHwfOFH0SWA/FHfWvF3mkr0LMW6nIeqIeoT8HrZqmRCvsf6MVB7mym9A1LP62WSqGlXQ
m2c5hJhlHlSZ8aKeJJj9/NRe7YGRFLLDRFL2Hd+l4hd1ENm2M4Esn7hOXrSdboWu0cC5jN/RONa6
0ahQM6iG4cS/u3j69759IK5KzpyTN+UpKcgKxd4JnybA/BrYX1fUVpjelh5hQexnkSnhpKBuDRJd
hTkduAFAS7R2xIKssNDuX+0xuShLd6epzUioT5sCFMvXuqsga9uzL88n2TuKeG7Fja9ptCCWFO4z
4r8rVNsO4JdrtnQwyEzl9nOCeFvJVY2KibCsY17m7z4NrB5XcSN26KC/YR70Hja7PedRRulsFDBN
zc04fssrHSvI27/7atiEcO2TJgsnY6o+6fJL40irmPGGqt7CuzqJ5DYjJDtSlKkvnN8dS/LG5a0S
MJwxNiTpuBk08KGrEcgGthL6beBWRRPzPmpvHedl4D3cesi5Dcx5Y/3JBznzqfFxr/tndi8T7lqK
wGhqONXb0KNTtOiPIjvfyM93HgrYtrcENvkgI/FUco/wOFrRyGT0qOGeIbGzydPz0yEPXeBnPDKi
pOiNI/jH3xgMsU/6TdF5UoM8KeodwOykf/b+jQbfGuHBde5SltCqJBlEZnaMgTv2uul/EHvoUJoe
LOXtz719cDgZDwUrKnFV5wbXMwYg4scCwtJT/q9Cgd8pmJgxpqJuzVzm4N6kc7sE8qT+ZX79jCuj
mLbTGAWffIolguA3eassQn/PDx8FStk1rieXfSqS6TFLOgXxvJczWe+nspV1KG3hbPBZw5JVGDIe
8A8B7aJxyeAGw8sLQeijnD6Chfnavqx9mpybORgqe4qFZPE8QzG+W1/SKc1hSq0R0p19GoMDluUX
PDd9+4Dumxo72o8qgaZ2i0oZoPdeIkX5eGm4h2YTb2i1dFg2l1/LogTUJSYWJ7oklhvQUtkaHgJl
ZEhD6LzILxx3rOG9ivVtWxt6lCCUq+l4aIX6QKCuObZcnMGYK5zGCpEcfes87WeZOXMci9GRvvsQ
08p+d+8LLdFE9vIXbP6/B6wU+SS+8rvpSbK6C5pI7YblWs4UerxV0YhkrG/3iL+3ZqnUKUxNbHLY
o7n+zhRHsqDrQ0pj7Wvk54n926TEJHaCizkuVw6r6EiPBRjEcXfdPOpSs+5zyziw96Fs8Hr56FER
efb7k2HF5gDLZh2m548N9Xh0Es1hNaW69umCx5IscyadtwY6gqD6UUjW33PkJ5z36UgYno0p9vCV
vyAOb+dc1KQ8nAtuGG65s8b73u39alGEek5IJ8J6TZVD59LFuoHJXCWy+eq5rp1+FwojvZold74+
7x4miEY1Z9lWliFjpoP9j6aNOrfgObdFXUyHELo+P21HveZoUlzowhIj0N/QMofmig7xKuV/iRIt
l1q439GGw88uVyuw1kH9bxnnMB6JsTj2WuiaHT8R2n7ycnOf25zdTdB3Ni0MR2NMxhww0vaRCtea
PwaIN7fjePRhWszdtmAM05q7EKm2RlJs1IY3gFrvgOEX8n3rtk3xdH4r0mXOjJ0FMPwLX5DvNd1g
hgFEW4AkYDDt8VpqRSVmcAWDCol3l1w3HcgN3vYiuHy3vs/Eh4y3vCQcSAx4zXWfNA0OGQSKOJYL
lDD96Dm0bmMgqj9pivYXnP67g+rzuxDVDwa99F9At3hHlaljj/XHx3awtPORb/cZlySlPMBMao0a
rKFrrdj/ZymcZJH4RkBOloAIpdioLB39ZXkQ8vC4bZbDt3m9bOpFHylVOLRgAgakhW2DKD5eEwk/
qeTuY9zj1Ark+a/Eiyy8rGImTEb6w0R0nGNIu0Q0ljW4kkpwr/ntzCSAvsxAeS1xJaiY/pHDoK26
fwKjuTkxzth5fvFeH5O6TsAEJDv11yA04Bbop5Saax9lfSL1BKySsRKWy5+FTzuhjhssICoAZYLb
EfdE9DN116PCRKyrhHltjrU5D9T8/vCCCMWs7x3WCj0f7XIBi5t1ycz01upNW+b/ZqkOJEwgH9PW
zB7rqsnTQCSQ+DCaDmWBq/Uc7xhX2lwfFpTjPha7Hz8MABll3FfO/XdX/pSUeMT8RNl07yUOrq6p
g9rfn8Z9JZabLWWrvn5U6BqcYZTRHKtlLnJD4ITSppKCWd7NCrzxKfQRpSRyyiREDebqDiMb+enY
A2XuU6Ky6hS/nXPsEKuCwX8bT/bF77gsI2izqQaKh00UzPZM/JuLAqI7lw+NDo4mrfeRnivFwZEj
z8t4FeCfhak3Fi36MIdssn61XinkbbXLyX3F1HCxJlFyrNtQ04n7h4ZmEwISr/qWjHX8Yz/eA1fL
skEkhLw+DFhNM6RWvI5glhV4FZphXbz2A1WUonOB2f0+N9sL5qPQ+253tE4xhqkPipMlLEt27vhD
92YKTuDRp9Yhmd0/tqo2aCqzEsz/6YdklsHTKjyoMyzHrcj5Pdv2Kza9n8efRT4HqLkaclQ8D1+O
xuyYJ1IV2ePhGQ5B5tlPITQhm32YWraXrS03KZsIppHbiM3adJWklpsk81NRqQmicdspd05zOXTo
FHNdDBuLd2IoCvFsaK4mTmv67/W1MWInc0E33N/iBjnd4z4YhzgN79esvH+ehgVuT58k0TweTiRJ
jis6+WFyZ6Xm8rQ1iECxrsDVSms7IJLNjbCRMhWxg/8JN+Mn62p+szRmhlWOlPWbZbKwW+guD+4b
rYLGTp1Wf/m4o7TQMj3BeNeVD4YA0GstQ6SRXItkBuae0nByIi2cMorQSmjXbiZ1wzXdRdxHV1xY
YKAbRV1lX6txNQ2zYRpsHtdrK15hv0Hls8d7/WzbDwraHIT3QVCHjo/sxm7HZEUT6bUQFc60JnFe
YpZmdGOXUIjft1mD+v4fBgPiNYr7n/lBGBzlALgLtGGJ/xG+V77N5yJcrICA2OQoNHQIpaHjO74o
ZtR1xDhCfXriM3IB/ed1drL7lagU7i4ePhiLkG6LfTQn0yDdCpv185xxne96d52YiO1kckp4Vk8z
Ct44yqqup2Tz2MIW3bHAdS7pJ1mc7r/S+sbXeQscJfeVI4mGAl8nw9mGs5di9+FM+xRgaIjU+j6B
iyToJuJHa9FAFxxaRuCYPbGsh8F8OjysEBfPwRzjZiU5IxfEIz+oEMfH7HHhbF/tssnke+Fpc9r6
w3pOoIeqT23lriB0lrWvp2wWRzB4KJ1SN5kIz8+FZUlPRr6fYbPHEJMGJl9QgJL0ySnunihGgW8G
gxKvHkPFOguISzG1E8eSOHAuNG5UO8ExDdDsWLxrUn0KBmfc2BbrbQRWxhXucQuTQViGhUjIuUnJ
A+WJMOOPoAJSMXur0ONw7MxiPyu3RddBS0soL7G6HGlB9cZBrpO0jJEbvi+Xa/kbeYhJsAxuAJBA
BRktEd1bATSHaY704mdklIPl5n1E41gA69sAzBLPaTt0ffo5w5PAzX6/gVVlUzPbK5gjJg4+aMbz
+pBHwlBFWMbeIQuZNfmqBWtU6ap6F11HDnjJMBJLCgIiM9U47TdzumqT6UdaFoa8aUUbvJd8zXyt
Xjp//O3D6+tihUKG8bZRfYs+nZwwWmiR7oDfB8smrwyMunsVlc1I4k8eOG9erHqnuIDVhWPHLGIh
rAQ5AXNGqHsLvneOhKniE0JIrU6FBLAtIrBKUbR8OBw4eOFi1YEdHyPKIA7ws24L/UUZgbO0eDJt
lrR0DKKwosWamKSlhtcV0K7XAlzhS7vrdEmQkxx1q9gdW29V0bgBfPHCdbQ6dnUH35uZ3xwKdiQ1
hrjkRDXp+fGdDwOKBwNOxAQuAMhGwTYtxwK+iiiol2cbefEglQyTFDQeJiLZliGc/di+/S2pjHvt
jX08GKcohzA9X+WG7QPdWm3tnuIlfDb5MaBjNXLcJo4bs0yi2951HtQSIVPu6zQ/dZcWQcCGpLLR
5OaJBHWoI3JmVjDrYhlAgy7VRiPIfnKuVW/VyVIMT0Ykvbo4dOgS3+SLghfZiyADagxMO+7jawKl
zaqGx2XS8yQU9fsa1YgBw++37kMmnKkfcwfaIGzN6E68KRyjlxJm2Ef/UZofv1RtxgPQ7Y3bLVl1
9o/vPrZ6QnMJDmuQrn2xaYJXPJsewwo5qVDf/J6GKU9UVab1KWkZ08ufpucOttXZ/qcp8eP7kBOG
jUsPEAEfd6F2UaqabrH+JDxVgkVgftbYsaX8EO723KrD7Xk8m4eohp5Fo0FBPDeg21/7oivuU5Wd
1fQxwEigx4ECLLBqxReJweepRuAhw7+rHw5zd5/em5rQ6mbFX0JLAo+X19BNoEfmo/di5PKKPTpa
lMK7y6imcvUuWm2eEAz8UltoLDOLsQqdjml9MXXZjHi1uizkIo2MIa2Z48yDW/EppuGIY5FCGSWB
wKJ2tu3GKNpBXxarWhQ7vtgL8E06vm9qglGkD9X8EpAam6+cpopHH7VXozbT7MENXAZNWwj1ev3C
h3l7/CN/hLCRfgr+kUNeFSGqh0/cJuJaFsicRedQMuk16OhWayNWCtHnWXGj7t8ma1Dv+O+rZUgw
HZUKlMHV/j36VTB71O1I1/n95SAyinA62tKm0iJAUQoFBlWlbJ2OOoLyV9QuS5wR5PflJ77nTfgp
RvnhmiwpbaH2OoLf5Bk2pfBuF5g/suZUsD339F/GMmRYNYQdsuB64MTNGBli+v8Fw8th8koA21RC
3plkhkeZ6dl1qF5qkjEY1ISQbruNGK7ox60b6VBbtwVNBeFGuWRs5/qFN03J0gBOpgHrL/KIc8Dj
L084aB3HLkjdoAPJJWZfKgNkY4wvGT/qaVCcoAbqdpKrSwML+BtMLgN6LQ5Y/DTwcep2xpPpS4an
TcVn3ozW+/nYmqCb8jQvZYk/ZOLWnstTUlPZnes9i8tO2nHpxBodL1lOmC74AOoXKOQsaaWoYWum
YF7I9ZoHTIAD8sI2zbQ/zBGrbDHtv6QDtBwRh1+ufXCfU6j5+qLstggyf938RJdx4DrRko2wTv7n
XoNkgDWJzvZTsSGr0rMi0eCvyw5+9bhaSYH4yxzLMqY2xGvp44O7tDkEC27bZWRDkbtQrKTCla0H
svuV1YxrIx9myXwzPebA3zTERc/9lsAZyjzbIh+tM30AinVZBsWbl7K85oMuyqQMlifo+vvpN5aU
d03zq4Xfw0Sv2DN+uvW0BS/L4f1Iy1esAwvv13eYZwXx7d/ab/YiTTfchKhBlzDFZV4yF62RFu3R
vH16gcijwS2QhVDA0Px9o4D0ggZCNZc1hz80GElDkiBkNcrhsd785pH2q6JABycixRwx1TfSbGHo
tIc6AmV1SsvFkditSumR6EVel1Dy643qMqd7B7xMz04Y4OF+QFBPThTO791p/8WBm76kej78M98z
XKxJrvUThq+6gwJFP0IdPhtRNVmtqUlPyeS1dCGYmLkjhjL15u04wvSIvMEnAEwGNQ9UDr5YVWRZ
jqSclDchsuMa6+qcwOFRAQjdkb+1X4pYStAbeaCbdw92YRqg20kjbWz3wBCa9ZW98/n1NSYi2u3e
hspcl8qF9Heu/58lrZBfGTNw0WFfQIIjF9g4D9e7UX0HTnV/uVSEaJ91yKCg34YRd9dD6r2iVk+z
bcH9B1sH8g8twiJf6DMTz38d6DAH5R/14oQlFUt4DpL2IqhGTaDF/gFY01vpKFtSriCBp2BdjBBS
3FFRINSSqIdU3keFpDiA4oW43lwZ88kmPERwtIm0Iatw4dSshI4O9a7HmSSg2iFcj3gkctVGB9Yw
x1+gb3eGwNE1s75159wOAqG3I+2y3v6hC6OcLcjeu61htDo++U7a3GKUnPCCqciujGT3UETdH41q
20gr57eBJTce2alzvOBFCYWuaWhmJ9Wm2Trx86vG2vapPekvBBKrg4X3acdInBo0IayIiiS280jw
WRoC8i1FYOu8nqdKckPJTJ1dx/sp8ea4P8z8znzz4fZZaQyeB42N1T2bZMSub1Jw+N8L+MYe76Yp
FCPiUkAN7k2p7c8ITU+Nj/6AbcUdU9BujrK+l/o8SRVTyUpghMAFY7mhz8K+TovxwYnXyqUv2oM8
sootvC5xjLSGzE3hNqnFooEGhMYOCxHwkCkqjkojyeeXbuLnXBc/JH1KihGvb+Z1rZh04BJGQDk8
eIUzXzOGoiaNIbDIXyT2i2fCnXF1AjY4ga6m6A7t9oNEDNJ7Tn8ctajsaftd1pXD1TFNJ/QmagFM
mV0ZcnOaZztrWqQZMhLe0A9YKk27jLazRZ+aZtXfv+mGUCakcN7URVSSwoEkJbAuwndXGGMCMeeJ
8CF64LSYociRhMAgXj055eYaFE3LvBtcckXx7oHqyeQyKFw0dg185ZuoB9V0p/QrIJ5yDnBESoZT
rC1Ajm9yx8ZUuJRoXgc1tnSkX05hT0Ws5BGZFgrabHicV9zbcn/jeVhtn+xjw5YCnS3ksoRIa5RL
+uBFNNxlDUFSCR9X+mZ5EvlPjn8Z+KNuBLo4Y7YLz4zhWG72rcwG6aiUYwPIeqp5cCahgejv44K7
ImW1zV7u9tkeWi3GuQ7mvR1pKVGPNg3BM4NC28R0jftgMzzP//natNNYghDT8qzHC5h61RUR+aLV
F1Jjqo2WFMMEZ1A70fN/qpE/9arltJJTqzpsDtETye1upfKkLGpW+ldYPuBQu3sCpjQ2BhRHU6F6
8LzqWsNZYJ6b40+t9MTaCWn0AwJ5ntwrdZE8c+NBPMhURIcHb6Uegz2pnkrC3RBeYeOazYEbqkdu
OvY0G010ZjRaBizvxOK8N+VDmB9iyffEPo3+8eMZQDdbE9zzzC7jps0dbBsvM2Ou/Xlz1M0+taZG
Qd8AC4rVu836MbdfxNVuIQ0FKX4Re/GbOmE8oJjqT42t+xeqsnAWRZqvb5XiqseurP1mITUwp3L8
WSfS2UJ++JVGbAHNk79ZFJtC/aTxE/2QYWO2M1uNyjKnYQAxq/r0cVXU+gzIuxRfXwaehYXozy/Z
O2Lll7aN//nz7yy/mFQ3GE9eorRtA4gGpY0PyjE/AURUekO4E+KGiF7NMOh6x22DzwRPtYRVuX3P
IzWmmsv2Sj0+C+RqKHNVGaKp6ATRPrIZqDMyLUAgY78BzelZuvvl4Txz17PvWuURt9jASxHwPdFs
99qOfDgN5xpq7cH2kQSUxgnmHxiNifA0+Dn8v8yxZ83MNlukdmj4m6HNk2dYKxCvjdpWoOXvjY9A
f02O18+VntONSf5G78naidQUmrSp9yCIZS419laZnFKt1Np++nX0uVvtbNa061nbJkrU8NYRAgv5
vyV+999WqqLN6Ybmm2Uxwb1Uth/U67BX/DIOqaltjfl1wZCsnWDHk5Zu5Y6s/kveg4/g6sPh6wGy
bkbzv9nU2O2O726hGYvLEHiUGpZs90VMAKYwZ8LvbwNttV86/arvRnd/eHLBIzw4ROIYZfqCNJMZ
d3/JRjvCl10J1g/kw39NAxUY+xoh7Ay/2TVezeo/LpXiszIOg3xxDe5duD1Ke5PwszLlEQb2LfMu
HqGoLYgNEqGZ6IbdqjILYQsjxtObOz9pfNawUwG6xAj5egSIP7ZsLK/OPXInUMRufJQEc65Kib/b
FKUk8mANKLol+828VakCrv/9zQiWSFppWBf1WF+B6LaRHoA0hEEC4JmEoZjIHa8ucwJN/NZvaSnq
E7cWjyE9577VmJEbzA9mJFX7c9A0RLLODXnZtxAzsZMqihwTnc0R9P6WgVbvRJNVF454eCwLe/fw
YzG2In2dN518GInf9kQil8+guhBu2s2KU9ny33GyWsSiBH46+HLCWgJAbhAAYTC7d4W5uE4Zex4n
4qRVUd9STeEb/T7roBClOvVXOi/P5xspAhN4dycG/mSz3SFpmkkLr2AkoQNGB0gN4mfQkjiauQ5z
tZJiLetK5a73Z3o920p5CvtyPfQ+S/BGHeai0b3bS9149rAxGHLP7cYW/A4KWSwXG1plmROJbALK
PMABlih3x0V2MUlpryqoQnd+7zR2ojGKXVx7+u2FFpz/zBwjQviAktSuwurkxEwleoI2TeMs1wjf
BTDf9/3QqtUf8Y9bPub5UytvGRkTJcjd+ToYBZT3pNdimX7EmAcSy1CnjZ937tckkb68UNjxfw7Z
ZcHcIWv1clQh13NrLJlmmL2SSSVTl/l8kL/EwUJxnAqPIB+kvgyGDBWv0PTrDCGT2lo45oVUsB0e
rTVdUMsfMfDCaoWjXKJWH4C0SCVB4lErTIeNPeCiH1QTAW1gZOdxJ4DghfY/+Wibt1Z13/U4NT0s
CR7d9kLhwURvmsn+rtN71zTJFP9rJsdCdQFhK4YdYmaRIle+/WlU/rFEET2ogOL6CS4PIsvu5YDw
nukxJZXzqi0pSLfM+9hsbvM01FuFppOimA5xncpv8ee2FI3P6Hw7fiENpJMf3+tKaSh/FuhB+Mu+
VHBxgTyYi75RiccLoL17zKopuiD/NEAFyeOSBFFh13G4aTQOR7Zzk73FO0GDbn/9JqOnNz4Ngjp8
f0pHBHHCxAxn4zgaIGI4ZPx1cPNnMM5VKs4j+JTVEdilVk1rkdLLuJ9f/7sYsbao5NHdAXGDF6aq
dnIUqGqEkt8+eKH1XIhyQeBpbcno8g1FRnMtlc/Wc4YuPP7zep9WwfgsLp5uvpIbnmlviDvHTUGc
lowEFlqQInR07xIDnhvZv0YvSkCNessZGSvkta6mfCLrWJ3tvY1FfYifX5Q9cfE5wvAU3dsS7/98
Hfp7baC8oMS44EYya3XerqoPypqHKKe+Dj5sPmztYeROF9zzUtS/ze4mGCGZX404vTQQblb38jvA
h4lA26Ei1t+ktI7FKd9wFq++1Sk+pn1gGn1Ce67Bzp62C+ls/veZTD0NYnD2dWVXqdStme/r1YBP
b3X479QUE5CC3rygdsNazvmsnerneszpZUdREuSSWunsYCqMeygFyNg7CipmfdpMxw99jhiVP/sU
1AvrpHVuIVm8yx1lJkB2jx+hiw3qYXkd/i0h/d2zXvGRDQa9StxFB3qEk863iVkh1lFvLnrs9NyQ
aWyEy2aCHIhWFC6cFZV2Ig4DG9MPgELfSv2j1qQoOGl+6TDL514Ow/20sUv1c9nFYVG0GoVXy2+r
sqz0TPjkDOfPqRIeEbVMu5U+npN3OcPS1cPhdl6ysjUzvM1bgwrlhBFBBdJIwW5KvOtTZQJ7Tdzp
WdLeCaP6z9lVwI7HiASA0KLGEtK67BdOEsFak7vmSh/dY3n7nu4owDEzrfWbePRMLrYhLYEUX8gW
GPDPLhzRCoZp7OlbsEDu05fbDqeWH5eYuBrfMSHmsMsbhHfwxedjb5mr2cNOLs5HwIy6ePNnD0/4
WSpCISFH8KK/KX7auuNBmoNs0RsAP0HzgstrKwmt6L9zQHqOKLAbEaAfRABGKk4N47NquTd0V1As
j+y5y0c8Cz7tntlb/57yCcOi1LxlpELH+7/jOvJynYFaoxyrfZ1b3MIzm9r4GdD4/aIWFGM9JzAy
yGtLgoiqV2/cUWpYihitbCU1sgR4bqykT5hiLmxy+TNTW9cBn5/xE5b+BDAWkIzwSRRAoBJLRxHq
1XfXeDWPFgxa4lV5D+ZvKgiq5EaYzAULsg2824oYwZGGmbHE8ypEvORwwO3v5H+RtlygHEg6rKL+
+/CZVLNE/NOXfGg33IfoGPtB71o1wjmBRJVTJs6FJc5Y2+nmUgNuGLlHhcZYQy/Z4Ec8f7zMnLLC
HL+fcUCOqO9LNL+2aAQ4BQzc1IjnhYtS6SPY4Vn+K+bi65grRA3RhVSf8iiJKmJTohEv5oBbpI5G
ZHQwxoccJC96nLRUZDUgAbwE638hGC8kBMaGnHVYsHkFsNISPRBm2t95PehjD+U/GJGs6j88kLoo
h33+uWsmbUxVJk17B6y3+1ls1zFZ6eyurxvYcKgCKnq5IGy0j9HNcVxg1L4NiqdTKh3R7x4fRh0M
8XhIau3w7TvWH497EjMhOWN8EMzQZxT8WtcqeJrsOgpT8v3t/07LluA18RbZwU+KmdGn07Zypjic
wUpS46uLbJVh0C4Jw3ckXGRJiwsE7MSOvatGG3O1exZIdoNbeUo3bgwWtAv7WW/NaSDAzldK9f4C
NzDTjg6kCFJ5UKH2pNpgH/UCuoQ/RYr8cC8qy+Y+bjGeK24faPgCzCM9wGK/bvHAFx+G6DBUCn74
9Gqw/ppiDkqPDTz21vT6A9YXjnLLqscUXq6ovbeG5s6exGPJxzonTrtp+/iLfDRKv0vYpsmJd/k/
29GIOkPMBQn6UaQpKg861ft5YR8+/r76S3ubLjGj97/oYqheJWSIFdKpT0/3C0tf8aZuvT2JiJwL
gkEjzGGI+FirmdmaG4P8MWTOWGnRFd+oIT2LFFMZuvgwyXxHV8MUG1s+7xWEy8M3axpQvRFoxpfG
84TsQVk0yAVGIBLPjdlnsoEkdfGS6DiQ5xvCI5WWsxeXvx8w6NMo1Lml6chQps+MY2PB+AxeHyTM
CouxNmhrrXV9dM8dp/sbANm1XzEM21rE0Ylt0TswNwBE5NM15o8/elvN2enrmK2K09xw9t95bLzD
RFQvyfEoHbHxKboHFclCcm38HoTXmnHY0mZS8f6waS2lNyzevp7hNbN0p2U9wSZWKmsBV0eXAt0q
t+ACAVUAWQc9453QmGVyO5i5qvSaMYGYAKKXFancC8Qb/epJUF9bfkZNptTJe5DlPqPXE2NCfY+s
BdzkTSUPKz3HocO//FlD+xBtprma1sygp81pkX9i+hVBG0chCJltSnyGAylFKn7x7WHbareWttUl
SCPuuy7IA8nqajIXXo2Mgr0JzyJPJztY5hQ9d8ywg/BDMHFe6B146aYVgYUk22DELULUQ2tzJtF7
R/eY+W8nVWggZ/Zorn2zAQ5nF+LgmXAcCaG6wkkGNqZbv2JXGfAgqEj/sOJ1OaAPnrBy1Moudmcv
cTlxd7ZfAg9D9rQP/mDiVWjgx5A6GbpOcWBNWi97GyQWrp/T+D6UjVaRoIJX7lcUWbra5NAIeJSw
bHbOsh3LHgyv9ajsQ3gQqiG1P5t5OfVf/Gm1IdZSp/1jWewCmWiUcfZFGHyYKw6EhenskdwgRmFA
MnwWraCt1WF8F2Z8AG312saD9RNkFQ8IVbg2XASixoTSzwvpOr9WjyUyquNRsjTpvcexHhDti1qR
tjDWYKE7wfKZeXFhDg1WUQynTf6Q5MOpzCQww5tQkRgPacZVh0WL/djVmqVFPYBKKRl3h5wn7z1V
/mhDVaUrq6pzxJqOPWf0yXDN5i9gSxQHSTqqOVdxWrltm/27/2WNj41DXDM3umO3TV5QyB8NKss8
hbJEJTJ6PSRDlrHbBg3xqGq8wMhni8nTIIUQrkghJKKzbhRbyI//3bbDQDJoDIBN/KkvljO6p6Yx
sWsmQQ2MakiCP8ulx1UqPLQRMiVWKIk5M58cKfAFSlFgIfU8Gi1GBniXrRxorkI2Uo5pq5sBYhr3
PBQZPXx5wTzNVu6LMqIQhXmu2EFY0IClorD9DB6woa8BK2oCC9JWHbRcXWOkn1GeEwUKA5hTF+it
9ZVdwEi1HObJKn1cuBKaE0VJKwNMBv9KJ936x43pJumZAPp36L5c6J1M7EBbnKLMTKTuFas2p1r4
OfKd9dyDOoo4k6as5r/QHr5d8eJnKf8qjy+L0ylr8CWZeXhqsAoUEfvgMCCBGU8yHTyQam+c85OH
sqCwJqBtquLxaJp/LlSTw0hERqeQnFgYAn8sRSNc2xaFM9OEVersf0hZYeeQXvntOkcQfJFobLQU
xYj8dHJzqT5pQH7nkkNKZRdZuLjWZy0x96JzJ/dGvR8eKUrdDJcdfhBviQvgKOmJ8x5NbEb7ojyy
5p2wpkHUFQ4qh3uTAiDQ/VQcU6s+6gF+DCZ4ROLjAXYaU1YUbsVxawG9TPENhZ6U2OuqHekVgxad
PC2Ko5jEe0fnNOz784ekXq16MNAwZF6EyNajH8i/djoWxOcpyVwWpg0AZfv7BVG0pL2IC7fSq1bz
bt7hJa8T0qfQ9t4Iz3NJfdcyjpW/ccYkGBLMTVwGQoMQqF3tS1UAlY8dePICcIZGPVPqzyGma7db
5r9Wh1fPuvOg7nsCX26AB24vE5rBS7v+5qWkIYu8PWKy/XBNdewoznpeLOeO+290QN7TAqIANe3J
i62sjST/HQX/MXWIi3OyF/JIydtH68mocPiLJ1/WJHYYVKkK+1nVzO1ZF5y2WqZHP+gTCdzTq4lL
MhR9mr0LvXmUktz8udTnktMRRJfZgZEHsEe2MCcNPzjtiJ0IRIlcBl1CAESEA1QWJJBvjMZnt1+K
cPbMdifYeBmY8ZAtDk/T8+/BZ3M6O8V7O24KlMWO4BHpTD+ffAKFwFRTODpdPLfyZuuhAE0HWTB4
b7uzz1s0qxPuT7g+ca3bYZd2e/rDf6THnOgTCp+tEEPJQ865df7nGV9c0SMYhf4g3ClOIRz4UGia
aTAwrruarOSCHBH82O0P6cTWxQ5hOSrWYuNJMEX2dvy/wHa8znZhu37nK+nar1JTylZJj5PCj8jC
SVvv7QUGhYwFsTj5GPpp3fs3CgGc2zNUa9OYZ7hdOOP9OVc89YGbPtBbdjdaQxRZTK09lZy7Ce/T
hN79ej6KMk17tS7nXo/Sv7HyJp6igK3gvguMaUJa9EOgLT+g/UjSTlqqyLuJT1sv2FrgBDfga3Yg
YoOBXKPAKi4Xt1NYvEckoB+1TzYzMb47cqdJNByJbsgLtDNTXa+QV3oY9RMceSSKd5yV5CYLnAdi
jj80wDyadcEVNKF/tYZbyMZ9wxY+aq/WSRz1oqqdH8ymotxm4wNCnc8mFQJxRv5tDsQpjPhM6xbm
hR0+PnNm8acpjxyPkW0+GDH4TVsuw4LMu1DOBgrdF9FlkeeDCkryOOl1iKDgKWjckyvCkkf4HDWD
D7xmtKx61DC9698lZLnnfyudCzhRzs+RRZL/99dCVhzh2O3eRIYNTfOivpBw1hvEnbsQmOR6Z9FP
JkdiN9127PvwO9rTc3GLmmFice2djE7NvYIJ4jZPsQAasYwdgWycDBJTdvxhRyhrEo7vDNpY8Mo2
3IPbaLz14gjyjs0LcHdzGRTgCBo59OWCFbXgUQKbBt/wH1ZUrmcTAGlIeoDzvhnI/hLeMv0XJbjF
RN7OPxGff4koUNp7BhJWJo585jiKhrLzyFq1h/ltBDRrhDzqYdj97LjKq3eQtR5/DpdYzNyNMefD
ziR6l9pJ1K8w5u0ZazrbyjKYFNjvHzPhgrnfccJzXvzF7eYS3dubF+ML61V19bP/wVWaWqIcGpoC
Bk1VPjY7QQsBs0IJjcKwdk1hDkKgwbcffd8L0eDQaHIfO5l0h1zIjuzdTgM+cEPUcuBhOHucSwRk
2O+kiMip6e4XCm+9KdeKKpEQ78PkP9jSLVmNIRk4DkvYg12+EQHjrUiR3VkeQv6fYLd5ztlK33Z2
iM+XrWfVXtrgQKb+FmkHDXgZw00kDCv94Z6HMOIy5XW2SnItC8Y9AwDYiveYRupgdAmsHGBANhQs
YlMl35WhmbK0XJke+2hP7zeQprQGx2LtAhto3/ZPEHfJbjqd+U3SwMQ29PJdIjAwhjjRBNC5/irA
EoSEO6zk2S3ShVD1mwBYKfqElFli5NJ7hyp33+gDzY5kX6lv8gEuHNYBuv6TJiD88RnKdIWwSv2y
TAOepJ/YeCRmivoo/2+sCB7gjMhiRU1HDWO9CO4mcACfq13IWoTVSe+xXjLRr4P526H2T9+nQnBz
Ys2u8TIpG8qbZ+tDn6YNkNQcTeJYrl4c3GswUssku9pUyNR3X2i7sG9PVYoBuSEg7Ivk1fd2mIwB
Z9gNLEbbU80LsA8xPiuG7T5jvwCE+u9cdeILU1kIJ9TW43bNjGOUoDnrP9HSQhzZrHR+viDoedvQ
l6AIa8lq0XZ/nAxsAbfoTkGHW1/WOCxfr1QhCWfal3y3v/ymXoKnnyfYA4NBAPwMjmgTcka4zcjL
HTc3nBJo1KbbYga3zp/sqpxZHd6pOTJO8i2M9Sw/FiIfsNXHxUi/FZR4/H67WafKbsN+DFCPACqM
nRKYuaDBvd10d3bPiOvxGMcDtxmWbuAWn7iCVrC4KhpvH1QSvKZQjtuBiM5ZVYIQG7v+cb4fGFI4
tNnOd8xOeSmL+gYikqZM75uQei+2jlDh9XXQw/aZ/0DLTJO+ZPCNSNwu904Ehq4Aa981CYadIN3P
nw2ozFY6ysmhBdecNbMxe8gvgPu3W/4PVYyKnqcxctmzKfpcdsIhtIk67AJceBBwHaY8u7tFRtko
k8gfGy/LBCUXGA+zI2b7MKG4j1sowIB2CFf3pklCubQNuCjoOZSWCFUV/9y56QDhNWCZUxak2Dtd
bgtciq+A5oFXc/jyfC4DHuUQSlKG6OiKH2Oi4VHAPV+xpIsqHkK+AvWUtSyIU5T5Po7zK/aa6lQB
8YFV95X5u3WdsvhDcNozyc446TxUyK5cH8v+zUGNiTGcMIyzux/NWY2RWGgVCHj0g7e1JYXePQun
I/X7ZOTyP1rGulCztKbDSKn8E9QXK8r7IHp9sK6KCZvtAidi/kLOaO8vMQ6irTjpZmIS8Px45RB2
RDHa9AGVHJ7voJrFcwCT3sU2m+yNGQSWbISfBuE1JIZFrq1hqo0u6tLS0UScXtAVDKEzxN+O9E9Y
caz8rF32L7hK00uolaxaYp4n6U6VMIWrtVxsfQQs0tuYX1iJjFr4ofR9nOZ/b4lTlLn3u16nHQLW
gua0GxGT5o1CH5tZqEF9FEwCWJ5ou0I41sfFkG59TPVVpwtx5/bunFdbEGulysFI2lwgTVJzlZ9a
DYrAqSE2CR2LDDUcuDbZwtUixzXqmIwQXSYSlYb/c0yNxoJttkQ3L6QiymfiBCeM8kNBxgb6YIUJ
edNpu7VXmHfl/GLR/4zF4YSB87IWgVlEtv1UupicxWxeYsLUUalw0RpVRMpv/iAfRjd/TWP16yVF
pND/P9h3pZno7zmQGgsxiHRX5uaP8CvNV6RmlDSv+NGEJ5lxf1g5FmbS0OHSJA2qUoTPH2cIBMSv
dXwDvTz4+f7ZLtOLehEXwhYQQx12QHygM3WaJiF00dW6Km3tYWbqji2AwYf0whKhmDw0qdLYScNm
HxG3TwMhAllRhpyCHW8QSwZP/wU03MWbDUZ0ABiNhe+CmtXw+zesj13fu3fr3BYS43yLvwQ7qBHf
IOWCo4IIC8i7AEGRN5SVIzL19Dc8uXwv+WPv2dOR1RgZP0m5PE/++Vs5VlF5xII+LzsLeUWEYXn9
iMmNFf5j/E1lSiBjR4+1aeBD6qQbQeej2teDj2RymR2pRFsbOGKkKd76Uk6dSMPuNOqwQCCcMUD/
mdkLWC8XEv1mJcaRQGrsTL5kSb/ybdyaVk3co+1rDg7cVnAYKYB9h05ePT3ipJHQomK4lYNAhH1t
wJbVxucxObfOCtOFujiSn0OzUteBdxgohFzGE27MZdjXPsOyCAkKk4QKLPYNFxG+XKr30AlMjUgo
lJBF1ZM6SknuQJFn4ow9EHMpMiR3Rc8k6nvQc0UpGBJ563oi7tPztfFcwupbolGJoRU0KtOKnuNd
VsFelGqFeOQc3viCJkTJezwbyUv4muTrHlQxm36a3ltZcMATjJ6VCkMIO/ekAd3StaZxfhIl1oi1
q7gDIcfbEDt6JIVP0S0rHQXzvfQs0P6fF9ErtPoNdKYtXNgW42ND84Vvfgjrx59LxpbyDTgw+5M+
GuQJ/qKgS8FmyfGtTGMUd55Tfy/mxj77BSmiUvnbSAe8Rd5oQfGnjOQFlGiDgTc9mwbBOE5qij68
G7UJaAzJwbOm9KRmDwoQu/2qwCFIJZqe7sDA5YoqHR521cEjuBjEFfp5U/xajzUCaICGsEQA6UNc
uTDJH+DdvrqVGDQRU9zbmOQAqmegZWNcKYhpsRUJ2cBoFz2NzWHlO/NWEykC32gxeVw0rGqW2pL1
tyVdm0Gq6YLBsqnvltR6h/bFO10U7Dz1hlBNlcjZKyTDseAJAXn3DGBgTUaZYrnIHXu+lNLvtlJC
FXCmxHt6Jdl2aiqwpH+V+c+flFbVv/wR2oClGQ0iEFqN/f2PCTA2zzxO1QCv35o3SEomEgiVwo6k
zg2e6uBlSX4MaOe6TqCidellE7rVjRAKdlvBDjzJQoceLjW2U3C9majt1Y3or972LzmY4ryEA2dt
Mm5Fip0t7UOYO3WxDZaqzxCD8NQSt7HV1fVc8qvRfve+AGMxyOTPCr4ie/rYGr8+dKbRNTqqy6kL
pYR9k+IQDKWYGwcn/y85g5zrwSMatmlTn16oOMI1DdkAAcaHH8CfieUAxXdX2s9mMINA5pTXiZWt
yuPALlHdirpn24gOxIeNpYK+hd7gOMAw6b5PNB+s/mve5JBCyJ4LUgYHLMjAdrQ33mWKurzVz8LE
w4XqPQyKN0gHI6JFZD507ae0O4piDnNnzgha37OcAGfr6FoW4j+lIOY2pPPiyn6KJ5KHVpMBurrt
9y6xgudZ2isfx9d43VS3TfspOZxMdYOjauNGniQ3gNLz7FZ5Uch5EWNkpdvyBsMWp1oXjHI72hGp
431zLwSC7GGvOPjgCCyKUYT8Ev+L9VMSbthd/PWOOkD0zjcOODv/rR72WuaWjK+d0+RU7a7CgtmA
Xd9Qm9+W6+29+oq5v5Y618grxTNroBheCe0e48LaFLwH4gAgR7++XDgs5YljgJcVqjsORyNeXqUI
Em1eDFyiZkFS+L7e6YW2v0Dm34h9du/Nnq67wWHbRLMCy9jtWa1RQh3dvS4e9/1qFcPamquh0Z7i
WcFfuEB2iv1b19yP9h2UXRBXSUqS1imEG8AveY7U1J8BFxa2gtpkBJ8Gzc3iYNhqMlz1cj5ciXQl
vUsTNbqK5xOpSsZ1SvEeKwfa6Pu5dzH7c6aSMqfkBRBNHzGc5u/OTgHy0rY2ygw7ovh6Qc7tsGCY
llwK4787LTeXldbpq4mePXdhRUqwrMzIlq71mi23TYezVGcB/fo92/aKnLbA3h0MkxN0mUJJ2dI+
3lMuvKmk3fsWeKVNXm23T5oNA+RG1q1l+BFj+EcF21YvK2Iqnj1OlyEuxh5MPK0FMWUOg2/eMijt
KlQJIHG22AFar1+IbIIaVWVxTpq/rH6rO6He/0Luj21dRALSsjdrvDrzOke4FIuBwASVfceQ3wIn
+myWcEmIQWMNmap312YJ0pkY0L5XOiZOH5jSCUl2jIxemrPw3pHXNuel71Ck7PVGZbH7IPl8V5uW
MLlgUX6zd459R+PyEJy0+cj29+4ccMwq/GN+X/sDANgOqz1KhiKY+UvwYnfxpCPrwRlQgOcyT713
pZPdMsLHrl3ifSRI17Ol22+AxocDOIcpiv+6po+iZ0dy0/FrbM/mggjjd7QEbJMTG+zt72RJjGxM
BSqDcrlrOpZiiXbQXmaFzrZ1pyGcS4U/jpl14tdJtThBusUU7uKQNQXgNXCZ32tl4SP4TpuHgTC5
ZfensXAaS3MnVkcb99O40Ql6+aFXYUSVmaAOau8nV9Aq6Vo2ykjg2H79TRnWC4rrUTSbT8TQzlKT
VJ6wqXGPRjKJMORiddKsNOhT6aPIGpZtbzpBCFlqOCnsKMUX74AQriTWzK94UHOLOxqTSylOsyFM
2bn0O0k2bQS0AuYlPhbrd1+TDAefn7JFTonSXDA6uGkOnlJt8sYwc48dORgWOPuZkcKQIFjht/Qi
aNdkuXQltJanG5rJ2Xt4LptBgASIv44I6ckveymgyG2QibmTeU+qHbc9rTy4WFyFeR6NDrYvvaYX
7OtZ6NhWm/B2bqI6LRF7vL4ri2Brp9fYl94Q/3Dx3nEJ8QU0RAbiJvqNc9pJSiiIfG1T9ASTev3y
VcbqdYTFcBgXyWTEW9n+sw17Tp3kJSkHWKPLSJ7jTGsXB9y1+bYH6d4nu8kWlL3rmM0snVtHKMKZ
YwVvUJfm+FqCOxCSleMPHpKecZ/HyQpROrkfiHXag5kudz2FiDo1LfySLQCZJObMwlCcemeeF/nR
QzsErq3ADRpIAghaddD9O18Ch8tTRCIi2UooDdvrA9zzFvWoZRuoBDLS7jqJDwbtyp6Hv8ksk89S
SKU1ASna+NKADsz+O8awIZu9UJ4VdEj/roR3WwV5E2OcoFTafNSfSc1Z3nOkaBkYAKfS/VJbiefI
3IHQzNitp3jnMvtyKPwgBz/VRhCUCG+dj+GCW5ZqHGbjd/L0cGdvzA5vV76DRtX1+YlbSZq3eU0F
+6uAy1wbpYh5Nj7V0Qd5y4ZbnlI4lSQDkw14+ScjG98YTdS/rAV4u7/R1EMK5YkSZskAY08bpDib
27QSEOGERAlPPfzbg5TalRnOO4Yevo04GNfEVFj4ujjU7XeJVOEvUlI0+AV0nCCGi+Lm4Umbrvua
pxfQRPP3MCpx81rnJxTx4Yu/wnXyDUVRXEsnB3KqjHcxr4DLMNesOG4gMmWmlyJTHDo7gtfde5yV
Wsraftk1pxOj5AdCagsJFIrTdjd0L1INBqx7pVtpI/2hNLdUalWaF6xDxD6jwazuPYkfNsGfsxAl
AEdEvG66LdMa1YqX6J9s9Qv8z55INY6TkW05FMBUbT8ANkmFdwo9waIMCA8TNcvdhk2y44btfK9N
Lko8UF50jJW+7SydmQwr4l9ZbPKRagfP+WxrW5HQEfrhoOnXxzUJ8TO1bG5iomtoSkTB4el1gHe9
uCux+3oAnc7H0rnoM5+avvY/OJPGthX2daI7UYqRAL385WKz94PmkBXz+bs/nMV3LfViXrh1cNsA
UcO8Qb1QEbN2XnPnqF5eLnbCgq5/foG869fpXQbAgTM+Rg1PPswS65wXNTQN+OE3Dyth0puBwDQY
Edg9kStWzR61vQ3y2RBxRevIYTam7MINarOYRSQmLouqEsmFXlVYjeH9MtxJQzQoec54bsNqdqYv
oiJlGvcz1h6KF9S5CmAGvKf0XrJPqU6p+1dKA927BxzrH5HjB8ExPCqDbFM5STc9//3Xeed/jnMw
1bQpp+ljNiAanaTALKeEAzJc/Xr+ugiPWAR8z2hc969EKsnQzeV+3GAKfSjLwTZuJtCfHyhhnQYV
TQhpfdw9C+e7R3gRzpIcfIli96/rdBdHqYgaCiCShM0r13epHIEXJqVz+tIyxOY1pk+0TYtXwq01
JUXF0mA0hPTMu4eH0r2fC0ZZTE9qbeSx5qosiW78l5wRdW2NZaqmSDmFnjaLLiWSsttHIhsLVeMe
KWJvrU3nzsRyjdi50R9WKFTxJhqnkI8qvzUL2JuAnn9j8gxApxES4yJ4CztMnYbrqyE5+SnHdR7a
CBwohOnmAzI81dESRSy6UVE7cLGfzU+XyWWeIHbFUALSkjSpf1GWQ2Sc/QXLPVgNf3F/WVMwN+bn
xxsLKl48WAqN7whyOY/sNYLwk0Vod6SDnHq+FjAm+Dyn3fRCsgbq4RBd/wGvNTqcRa6VQZuJmrxz
9OqUS1wY6Pn7qdv6QLwe90B8C7lw2WxTjntlYnQb2d1K9JVgnGPDioZAwyd7po3UjgHCdsdSeaBr
Xks4gF3VJcduOhupQvGgJtDBQ5m09R049Ohxass9krRILqfOJ6U+Jaz5dQGoZdawoHJapzdTdF34
sVJndcSj8TGs9c+SRP2yQntZghEgq73XExLRqxnODdTRgC4XA5NoVqvouG+Ri1sYTy6dENlTzJW4
f1PhLAPgjrprue0RLKFtDq8EoJWoMuEHUkQVYkgOleIODkA+y3j+tLD7+M/FZfw/9mjcyglzeVm+
CwdYvP/PFTOMCAn7wGkL8D/78Yb0+2iNnNCAH7c2826jRNAP4TW/3+bEetNB1G0yisM1dwj8cMwp
oXkORKv2IXNTFM0TxPhOo4tGnSTmvFSeaktaP1JXqv6trRAxhYvwIXKmtmEuMJY/5F194+2zy31E
ggjXwrYsowAzOgNvyngj828CA7sUgEitx6+o74ZwikfcSpz4zd2I46O3h9hv4l6uVTiTRBkIhy2k
rkzczTOxsrYCeAlAP4Q/v3GQIDJZ7aVBsMw4cqWdUXghotQEmxwWyL/ZqAAd/yO6rEert8HfwQw6
hp0WL6LgIO5+lTv6H+f2lMTe0vCmkSxI3Yv8sD6iUd48bQIVJCv7sTrpf54HkAuWI40z9g/09Ia0
fZ9BcMen4QKO5Gxpx0ym3oj8iZkjIukfWJjwyxrG73bart119D3zcHG+jatKdvUHO0kU6GDiwXJb
aCUnli/HEf5ZydM1IZoGUfLhAfRv182yf8AjLJrnXCg7k4os8xIKX8uUQf702xErY2Z89nYSk4ge
cZ7E546f1Dp9VmGF1r8PDwN0pPLhoyZkl5RPx/3xFEVhCELZAg8l1+F2ZUi3Qm8ZbUyGY+U7X6W8
vx7kbjNze8AvmjtAyDJ0LCUIpIwOCtAynYyoxrUQZ43N0hq2MWEXPvV/+Kis6qlEwGNf+yo49Fav
qQ2e14FCvM4DdD4yaLUvBeyRy3Mb/2zC2uD613uyVvM90BETAi2kx9bJhGosBI4ixCVfLYe9STYX
6XGmERSjmgFHTVApt1cfy0NAw6xO3IViri3HLnowmaMIVWwmf72dHrOTV6/PRNLGakvjCjKaRhty
aKKrQYbMUOkE5JrGCD8lJfxVy2pwzMyAeGRSRoYi25mmXGzhgURBzEc/F5NRhED8n8Iv45azTWqx
m1cRd16iNvZ0V8FirTdQXQsGNAgPs6E920BIVHhER+V7b4wURbi+FdLNfG4pTqI0tdBt7GXOITFE
g8Lg5GGyNe6Ui4Kd4YRteb7+BXdMjigxHjeE5vW/R6UaEzRXAPlrxw4Jjm7fF1kCQoqCiVDd/9nd
EQDDsUuuhlgoYUdpK3KdHEzLBLgV38boix5YyzyJnYHIzFqZXY1cl/cl0j3wrO/HyTdrgXo4L4G4
Gn+6/if5EwIaVoDshN8EU6jKazIBM6ar3Naq+jaQA0wmzxrxtOKtqCHMOu7Xm8Bupei6U+oU3uPM
Ta64mU1Ow/DYo9O1xei8m5PwYW8uYG8Mueut/RN31Lewt+106LkaicyWsJCWINt87ml7cO2EWxQ7
bhLNXijYzSmXKIBevq2NNcG3Tnrt9R9gH7Wke2UC7nWxPp4uSvFYyoGAxQMxFLmyGab9uVDQla/l
04Bp95kHlZoLfTuTCH9cAOkgmjCtic07ZsxCzTjxXub+j/VqXSwjgnmXlbLVIAnmVe/GzDVj4N4C
OWptqh05GCsRdmREUdIi9attuMkBhZEBeFbquAV1ndsow6nVh0RlII9GXuurujkTiDDNu7+ihLku
OL36qszmNzFjvyQPkRw3URNR7/rCxFopfojXW+zG+Lr9iHnzVNQ0/FuBPBMmkAeNwtJ9uRjihh1+
Tyun9TmQijq8GrsSlouD+D8veKQ8+BKfmz1iyr+T0KDQ8PfWUiCA6r2p7AvRzUMMP6yg7R3sA33V
BaztXxJXKRiU2PIlJ/Ix0Qh8AS5Kw3ykTph6oRSBGKCOyl2yUxaI5K2YuH4/Jtfymi1zzkmnZvkF
Ip3YzfeC0UyVmeYCnMy3onDqADnayEgJ29b1nu8XEIYHfPjwOIRifjmJ0I1ixJDee98BP+UVr9Y9
Or8KpPrLP8khlF9ZR0wdJWIhNalTERIG9ZokUkuCgLA3FS5zQkJJJeyXf5K3kZngQ02Md8Q45HyX
q7En1V1JkRWK7TLrNVCbroVzaQgiPpuEpXPp/Po51JJtbTrD3Dw6IVVMNwiq/dS303DXcRxwss1e
icxdeQFkZzWqDBvRqzxTkGWFoF2AzYhl8fmiPkwfvRnSP2zpqfHGPzEAoxKjnrfXdjlySeCNz7RB
1BzoX3wqtREwC/ISZctTTUq8bdaOpEVeETcX2hFxV1KJS2nj0blUKlfH+PCP9hxdyd102Md+ivmg
3z2eJMSms7Ud8wwFEM3bdSllcTmn0VTtkhgLig4DGRIaGqMCCRqr4RBgxD2B5jP9pJyNUSxdGJK+
kMoU5CHLCSpHjpBQeK+pi+HI+7YZzi9IptHxhLD8uoTQOgxjBLxV0mdNcUf9oRSAZpt6wU2MZ5D4
IlOODW+GMoeAydqyrro9GJvTz9OMGwNUCpLcKvs3nFvBznX1IwW1EMysj2Ch4bY0nusMvy45565r
wCd6ddctANs4LPBJW8wsahsoI/+7qrEZzM36CGUM3kF7pnRtnrAS7nRpfhl7sQmNQn+pcIPgxjIx
jMLeUgbUX8hrF+rfJPAV6+77W5LrDOfuhOk0L7wKQ+04gYeV9jqNL7z03MpqXxasfGccav3D3PCG
Hw8gPxqgn5lqhGYDC7RkiWvyfIqHV8zj48ntyD/iiStK9heEWd1/rfGP/Dv9uDWvzAK81Flpwdtp
Xn77OXQQOhSixBKK11ex4qoLN3vmue8laZCFLl9RsiMwCvEYi6atyUhLNWEFDxkgD/zXg2vVFXsV
Jqx9njV/zF3H0+ZaafB41qWmcvc6YxWpOr2Xzk69ULUtXx1E/dhcfus1fKvicuJfzJ9GM02pjtck
qjwZ6IL+m5fh1f4h6LpkTZU0V9Y1O0UamREqu94iIIGIbVzbgQnUJHMaU9yvdBvJ8lkDTNcKhJHw
Z2mDFHUUordksIsBElF57YeI/5rHrfMT+X0MeH+zfizrO5p4cfQo7NW0ED9hWP4xUJCCDEPW+i/L
l4m0SEL5lJFYq3KZc3GsbfPG5lG8HmlHn8YXG/44BCQi5dZBvKAz5Bo9k6PFObxFzzjv9m3/G97D
g9f2Nvb53Tg2lTwjYboMnqv+PBhB2eeMSbty9B6FZBW9zcpdrKguAyiejNSZIexUISgJh/1hY4mR
ZaHWg0SEWwbI1Ej0TxEfoP3uj/3YQRriepmYVbtX3QJrMgqovMvdtynvVHaEsPHRwoLfQySoLWx1
2ssoP6l4xO0W4MufUvWCzD/Hn3iJOny8p3/a7KkBcyiN1wfgPu+rlW8wRs2yH3rD+B57P0aSMD3F
5O1oWvXrLVTmnXlGjYi4VXiTasoiuihypiT9BveWnxaI4uwy8v5G0+v0eNPpBKoiZXExKIvZnmGy
kB8R/P52xNFu9eTDF8g5taqc5VBJSiB5e4D5KbGEAWt5Lz/xsbyOuZcK4hrvD88mikqsRegpN31r
u8feQed821rAP0/8hES/LtdVSGz8mm7REHh5gCV2zTFOp7p7Vd8F5DLYbCIfw0eJnqDu51sEpuZA
Q9P1X7sYxguyNQ3t/ZkN8X9n27bQ3LS67XSAP2tABM+E1D3rG0AAo523A5u5wgc7a0/yiUaGmMSa
qbyNEX80OkU8K3e1B9NLyfl328UC2zBqJz7Mg1CjXkvFA1oRness4e5yBs9LJSmDSB7Qs3dD+fED
dARsd9yn04gIZyEUdC7IylsGhx6sU10c6T8TEkueL40gyjWWsbysRffyFLRGitHdKMda1zD/lmSw
n02EcnpGkK/duOpHdV2S/YO00UbRxeHkAPYPHEfgnygI8veX1/USDcEKQ6yVAD8qWvtUyVads8Oh
eDNPI6vOAqYNI7QNsSj8BFftPgEERwthF5q661SyK4N5sw849X8t0J+Ck4iq8oynZVbxgP+aGOtZ
WbFWF1DKccOXcmGZP5iP2IhxQKXYaPtrAZ0acldyTnyB2oNq1fBiBkv2iQ75EIW36yF26QtOeRWj
J/MVUf3w1/Jt20e8I3qHhSYUMYeBhz1o7zmvKsvaUzkuWeWLpLHGXP7TEeaQo35xK9SnTsontwcj
DTnT8+MOTOa3nxxy5uuqoD00y1Lnx7tYe9VXPW5pbteBXUhauTpqKrwBJA8lyAD93nmtw9ZOaSER
B81ht4/P4OFHAJ6eUW0uA4UX4JytTWjSFPc4Wc8nt5kEaTTGrXJS1mY2piVfGcBK6pflvgi5/+Gz
yN0tkzYh5bCZSOFSSDqo3mQVtDMlQFiK5Ze9sA1bcL0axWd16Sh/RizA6YctzH6USE6jxRSN3Bte
fyO5aGAcpuh1k5ay2C1pNoKl1wPDGLu2ar8JYniehtnzOkxZjplkTLufokLZwEEXBGWbauqbaIso
tpnmqpk+SkUAtSJbzZsVaIseCn4X9gVa2La/oUSZdATkFdrp9q++Owc57FBQCFu8Bf4CU1NwV/0e
R+6Bk+CopEn7P/al47czaAw1r0pTQ3OPlPNCiF5Wu7tf2AQYoS2v7vssPtubKU52wFeTPn3FaeiD
7+ffq+surTHY5gZMIvm3P92bO8JSBC9p07FBpV1rJsllS+h5L+elva5us2Yk/Zdb820ZrqCXFw9z
8Xa9CV4Z4nzQ/Gh/LUB7DWNBJUN5Y+su7KzZUNbhh4FFFPwOkvoxShupF4cQhARANyP0rtvMQOih
OzMbyMOPNYHXhGRNxRez4LT3G5Guo1bU8bgyLmPmKk8aeGoA6rooPg0soB+pOk4sVDLMBs7roWpa
X4/4Dfk0NIUkXYgDEnsNz3jEOagvdW3smkwkxSseu8hM5vOTbEFhJQY/ciZO1YESiCKMaTvDnVz+
5LD3AEwIFBDNm8sEf7thzWinitr/bDWKBDUEvjefrBjCCFyjOesreDyeSrr+sR/QPKUadutE6ryX
nGdDJ5ezHxWTUJxWC2WTJ21gFBKds3MwhZo8nIQI5LR7SdUENpcMTFbALw8X6piT083vDzqDtQ3T
qTgb9MQIl141JYPEKLUz9J/521v5WYCdJiSeJO6s3uTohxklxFcouxuJhKUIgV9AZnZiXX7bOSU9
P73p5nWs5AUNIM0i2BoNxX3Ixt4SV0ZY5qNP7bJqseouYEY0zkBJUdS498zj5qyZ/75T/eXSRRtF
rUYU9/jTdhr1UHAneXipC1cR5K9JR42cqCVzumyZcEA1gds6Y8W4baFb/OMnT+enYdoHjNIbE1aT
nsDJIF1HPQx64potkUOqZ4219L3II6YPzpOz61VXQO81UVfm59aScUj6K6khhcgZfokut5tvryLK
xrtATZjymneTqk/0BKop6FrQ6JNin6RQFzWWfnezyNk0usjyeb6wqzkbxjSrxunkqe0Ho2JnxJmT
KhSeXj9QC9LdQ4tpbpqctYvkGYvWRG2OqFyb2Z3MkYO5qhGomaw8eNOSO8wZoHA4lwRuz+KI2AYb
4VMHm+unuQSki8/UZpIdOiRXru9qoqWXnS2Bb1VcJyFHKc3zG+n1IwItyNJTaaWJSjRgkOhhdSo5
HiPGxXkpNQB8hYIqRE3ZfFJqI1niJU4xAERGQpIl8vX4NL5PJUg5VXvYkhh+nGyrappZnwtkLE/F
PgX4IsfYO/q0I64DpPGwAKBMgyrMPQemwgn93Ds5nA1nA76gukHq/yRCTUKVKlKn5hQ13WqTysF0
iYFODMYsvaUl09S0q3+e2/KjiFj9hOiHniqYNIo8L7W+RKRXrJIwGx6aNYJNLdCumHGlGJ74GziC
/JnfM48eOMgTLhjael+Q+X2fVgRjNmD/OCejHqozbLcmHkK163NNQYYLwoVXb3C7QfMqRGWOLh2N
SfTg/TcIBgoawWimdCYFOOnWXbZmrh5DD/Z+WdZS78kb2DlkACMYqudH0zH5QQwri0IVWerP48gA
nEYWtc4OTyKSVWR0EGmwnpN4t9Dnw4xr1DA3kCra3/9uvictyicMlW8KcQ9+YUfJ+w0UkcmN7sq9
IAP3wWn5OPoV3F5+ZBexpw9sUDBBSzGV6nRNqNAhbevqvusqMjZgl7MBzELCdvXZbM7a9hxYx4tp
W6KRWT5RlqqEdxfal/C5x7xcobcg9zr0Q8E9ntoD2rBUjj6QK+gI3VwXNj536DNQNVYR5MFzmOmi
illN4HPKj3YEFDsvXGD8sBHK9h7oIUd/2KE1ECwy9cn18XIwmCohEmHIsJ68OeAshMuEQ9rYOCii
dob+1JVSg7aJ1blZlr0R6Su7Wl8YJ3xuRFfUkroyv8ovz/h2lBFKTMOiKXgd9CWv1DlP9qUn8WZA
aPirgrW3LA6+sSRZ2XCPsyCrpFCslDkZzaTWIC2UYOZ6qwxWeFkULpfF+d8NNBk8gsP4xdmdHwuK
RRFi5F1BIQdaMdUqTPLsr19bdsjY5w9qV5JV52ceE8b4rH+34AZz1ypcR5eCSTfEmrlDinQC4m9K
fKATT/+1mBEgk9LK4F9hP+VzMnB2NBvgbH9Qo+tQFWs8cFvVD+h3lrgHUO9KtLJMqGJQ6fKeVh6b
IIj/4GRLH07pvthh29Wx4lzXV7kOOZgbfMO1SSPam1KWZoLczy85Bm0kKYBpUA4kwKtmQcVa9kAo
KO9v3960IgF34JI+8A1GgUfrLnPe88gOcLucPqiIqSEph2IIivXZp1tMVrahOFwridPllbmeYLTW
Y/8ZKOjvZSfZA9KnEqPyUA28oPNspUwNUEIaYQbVPGfz8JAmCVBwXCoY5rTubiuPg9eQebVYj25P
wo+J9tnj6Nq66V2XEuiwtR1wPnQdlZNSt6OrLy5zBrnND9sJ9hk9pGq+TUCEvT4xi4yj6io6cpZe
nFjdwpjADHtQa9Bq64d/6ujwzswNqrtIiVmj035oxA9h6lQ8837u9wPMSm54sFEXB2Y56+PcC7gD
YhRwmXZUU1kUqlx+HDgf9rJmXdtUZ+GBo95wk+VqJuvC0F/OHMW1D19cqemTIHuSDdJbZGTl1WNv
FiS87ZoBwBnZQDViWmR6vzNz/BFrHtQ3Ev6jpIj0RUiDFEQDmv5KIkmMqzeYOhNtdWi5RVnNdOqa
/7p4SrbDvo8JGj+QgKMS2Wny43JWkaoMTeZiRQxJoX97GHjeoG2lQOV+P1h5PoEp37fK2BbdORuo
mzAevQRkuXt2ra6E/nXcIqKFtyK40733TY/PJp9bWD6CBVbjWMN+/pOAmJ/u+qmBlwzEI+Pn44yh
kPXlWEzhr57pf6iQhc2Exgu+HdeYKcHUi5/L7MBUO5VrdDvXuJPSCsVy7pMAGpuMD7TEG4SZG6CR
H8WQSghH+cSYPeQc9CugSz6bhNqKi7BGdLw77ofEpO/9Ban3raivtoliL1q5utW7RmYPAfcSe7EB
t1O1BskSipvE+mcDvr82l2d1tMVYCEg6injVesLRRbDrZ2wSPh5RFUUISU7YrpitewNMTt094WSZ
hOhq1Wr8zsPvYDYKCwszN5Xlqse/LVgoEF6FKgATaUnk0Ve7X4d1PjP8ntQMQiaWCFqjslUSuQF9
+OdMk9RtYWdEbuD21jW/Lq2dJeBpr8StcafykeQFaEH5iGbCJMEXG24kXvkTFIAblmwRd3lr8zIA
RfdneDSRpdjKQDHEaAPWmT14n9cMsAJYFRn3pcfCUaaox4E5ogqcYyV/Ng1zFw4i3JiS5VXEWH+v
gEcZRT9LyXWiFaOMj+TH3sOJ32H/UxcENsVOyS8y/E4rgX8d4D6muZrh+bSCzAH787ACAej67mRV
Rfjy/NKvpDCsjo9JU3e/VUWd419rL2bpRcsaSy0h8jc19t3TvndjQ+XBX4fLjVdRXqJeloB3kUXd
q2ugZWgncJ8XGO99xw8HhHvKLd1hOcjhE7yqgBPmCntzI6dEfu9b/wMFiX2APN8ALDw6Pn4E2jNV
1w5JuoNf/oiwGR5Vr2PGwxzJPs27yOVg2Eh3iupbt2LRutDUDX1NhDL3bHDL1kizOtGFkkNHV+4M
Soy3HbNJjh6XDO2/A5E/ilbOp9YqwD56gH7wkE3xTf0mnqmM43aC/0h4e1Q/e4us0s2E4XTpR1tv
1YZZ1hQgL8oCZu7lQrCvXT6L0lGTw6L3xdsMuvNtIiEvkz4/d2UaF16D3Aka6BDsUz0SIQnAZ9Eg
irXXauihv46pTMV+IGk8/Zo17vpCuu5vbHZ2y/CZX6t82CvJMt6Gnx2bvDUdYf3l45cw9xZXzenJ
qhoF/jeci8/IOcE+yw6yVurcdjnfso8CmIBrLxRIbtAyZTgNuJ3zBj4Ee6Z18z+lWefYNr8Fwg4I
AKwNL1sTglk1t/Lih1m/skMqVOR4RPAK6ZR3VpK/Sgi5FXCLygm0WCTN4ALKdeCVZKssh/x+etUc
rShFDTdW13BEjn0c0JQcfrC07I1TnM8w65HQYTL0Rv1cMwVuRrLJW9peNi6V8FpKn3cybNrbMnIa
P6x1n+2yCmnIy9wJS6lI7A3QsZknelNEX9RdRvJiGGOmaDPMVm5QfG5QoUV+zife+G4j0DtPf7lp
JVXIBR8NXyIbjy05bES+EDD96JS/qmL/BZUdfwPTdK+eUARPeb+f9qNrSXFZ1K4Vk3KTIp/IUWxl
94hPUklk5VGASdfUivKktKSqLN7CKi2sHJzCwIsxfXbtJU5q4dLPD5Q4VMN3zsEnHVUSQ+gwcYA5
XXzLyKMstUcWfTK9GYuDxKYunIMFE38D5BkjycNmnscbVq+c84yMOzCtrd9gFrujULEN6s39Mjox
/0m+N5coYB5JfOslgyik5+fqfAh1tzbWERhZAULZm6eQ1RcDLnG4BLjAfye0lPvR1KP4jwsF0Daf
QpEnbaH9fffaU5lLgp5Tzp2/chsdeAyhRUqazw0zD0tx2pP1g5OuZBIe5gpOeLe9Pooebd417QNO
5YqLCjzJ1epgWtR59NYsMXYZ7WZZu+FUKqgzEaUwAViLRuwnPR5+8aOgXZKuV4X5ElkeCDqeA8CB
OFGOL/QtFawZaJnACVKGt3MZsOjtWS77CcjB63omaH2JZwpMj1JmaVyU52a8Jn0BH4ddAYJ9QLCt
WCAq2f+EiZr0ZzSS7ykOZFFAJRk0bRPNg/G7LSXBID08gwmBn8NYFPhroU7arrDfwDVhWu7Wz3mz
q/NyIPT6MPEWeAIQQj5k4qPlzKzaD62POEO3OTrjwN/WXxA0dZW0PeTgse5I7y9NlhZxw+8QXPjk
Uf004RYL0E0ld45AuMToJAB7mh2gg8nzVAoVIfEyYMNqh220bCj+CmvwKcP6M9TDrAOy91Q7UQ5+
e2kLzd+m/ZCOGB3EP6DH2otAI0yvetYHU0U8Jg5ZVSmonyX5fM3id4to9Mc/1NMvn7r4ikTHnp5H
FCwz2Gx/sDu7T4mzXN7lOt+MbhIwzz5+GonMtYx9cHJLfxYAxm+d5EMmNW0CDJHQPGN8FfCS8WOq
1w9M9u6KxnagVTYcONrKgPm0Sf2UuKWMAV5dyQ0qF3gjg7n+v+H4ZRTWWcDqsjOkGV9Bt0doWNtY
QN8nt2ORAVwbxE6aYh4bcYpvmZ8ocmrgq8hB97RM9U9k26t/z2m3caWuxJqa1gaJjrLu3h3GKRTg
76z3FiInrK+wLOppuXDLeNVZfzmSnH4OzP+85Q0z3dUXg1w31tAo2htPKhQL6wBatcHkuLo9MpZS
33FBLirh/fUAArGnTR7o0toD91xbOg9uw2xW7v3Bu6GAXN/Mov9eGWRGf+zKBvZN5mdj0nqJu9U2
ujnxHJH8DyWU2aiZfxo6igZVeHxNon1m6fUQKoiwylawY61lRsB6sIkTHnXE1RCtgEfS0WwVIEeZ
wCEN3+WK3YvU3W70LqCV4aWRoE+9bOimdoa7+lwfGYZqhBGTlc/SEBrhsyrwakdMCl+e9RPlw4y7
b0s4Xjix8jojBDinGuza/FdqKpqhs22zAqt2T+pB1ghT6emTsvHdixwFNjhmmva0kUoeeJC4DtHO
PwkAfRmzRW9jKkWs8zTNRJHElHyTniodWYtlHjoZtdIpPcaLKcjWNT+r4qeboPENbYRwC7rWfuTE
/NEuyjQZl06N4oxWaoX8UNb7bjw4faWodut6qdBf8fyJLsz5PB18LjL4ppjB3tSQoaQO4oGjaH6q
66cRs8UVcZrf87mlNu9WWu3FsllfI//k8Ag8jCum+XXYadYFCm22PZTQxE0kL/c7XZyhMaeiB9Zp
Aen5T7MuhOvMja2VvNSdacX57Gl+pjSgFbVCXxsxDMfL1khy5ejNLdPsaN3EQhpPwsclngijJU5P
9yjwuOASsX4o2XfKSeIAroli1ElLDfv776S6rdcoQGCetFbghOQucmAcDT95UyD+EkLV682wCRBE
nyrCTzm4ZwqpEyTFU/kw1UMc6ghkN6snF0OsnkLHQbJqlc1tVT/k5VkQmqBrp3YFwkEC6+Tv4wca
ZJtcjDwNJQw3CnSaf5U7IdU0R+NYKk4olGfrO++Zqyh3wAx9Lt1dpsK2tW69vet/97/Z0W7NYi5W
/mq4McqX5bzuPxM0+63fylGTl5dHCx/Lu7ZD/CgGr1LmBTnAVSd4fBytgW7TKeld7X8ctfwiJzwe
Cw5yJISmUHBtWcEh3QQWaw+L2PDEP+QDPJdSVlnBU8YzU8TNUJKhartbqyKBnAQr99uG9k4EL+jH
GZrKaRpOhi6CFWNT+Oz+friOZuCUQrY7Lb65temLH5MdpbE1Y/DfJtyitjcXOEuL5NPoXrjlU6hA
4jo7p3HpeI7uGo1RekCfxaoRHaJ3S5mqRr9Uo5QaLsnITrz8MHEg7f1j8OcVL1IkyBLVhtdtS3Yf
5PRUd7VRbOhURzZSwZZHvolvi5/BlaLe3gml3XqczDlnzLjug4CDoq/8rg+3masHZh3KgP2zEulW
qae7GV0snPhFWkW0GxBIfVujD6yd/Wj7ccvT6pTjKB4Ew2G0pqguqOa9KlTC/9pMM511xECjJsyj
5ku50HjNzJpRVU78s9/3CMKzM/y0vtEzlNACvm3DH6hxrKQwjhgpziuG7p4a5VjMOklkZYt+cMo4
KR+Htt5zCZLR7MhSApEsKFHLEGg6N4Bn5B7gjyGXz6TwWjnjt+0s26/uNdXGu9x2/FmyZD4/B43v
kMyEYmeSjdsaIb4XZPq8GSeb4QJT9R8yJc3LCRhc+Wn/Gtz5tFiLOHVY/58zxo2bpGPWB5Gfgf4j
UoKyp7/lOxvoAT+dAZO1Vyq0yphnj0iew3uy8riXGVbGhaEQLY/dGwTeY7VoAcqYb7GZRelZzo1l
9e1XxM11SuEIqNlJ0aSUtVuX3bppBYUVAOTCfPwsGPzJISPfG2sGUszMCjpnKF6UUb3GfWyf5vJA
T9T3NhUycrr39ghkGTw9T8tMMUry54bWtuVS+4lA3qBx/K/bbMK7K9qpzNWTmegveimzUqtKXAbm
Hixdk2dhuYYJp327vOmxa6Ryue6eqyuS+kOu1fGNCuPPB9L2zZEp3GqT8cz+LYgS5WON7BiuoaRi
Om1af82QeNowyX4e2jKsEbRxgYuwl1znEW8G/Ho1xtGluVye/s0YAwpy2ZV+DQ2zIwRNDC6LQWOG
hfVGGmkRKRKmciO7zbBZoirC6q7KFZwHzE8zfo4o2EWJftCeE+awHVAaWvhYyQMYhX7m5xoN5Chs
YW2mo8xRuma67gXbSlqkcdYKc7yc1nfwVYBuW+/5xIq88YHZZ3bIvAuhcCpK9bRhbLxzW+kw+HAu
ej+lHPm3/JfsOKnGT8VVu+fnAdgsxqneghvka++tJzUa/GvM7hyFs01Vf2YUaMhMRI85gTvHRxHC
8YlFqBox4iUAp3IDnsXR5k1G3dYGblDPKPcFP4Q2dkR5KBKgOqQmMtBiWXMBSVL6laq8X5QQJ0he
aVQq2r6yE8hebTZap6fnbFiMCOwfMpNTrudvNVmknanIkNO/gAOISS8SGe96klXNgmocngcn61e1
7F9xYIddScd0k9g0pF6+VwigsmTXNaMgVzlNEpdaTSI4/20jAUtjKR9MPtrkOOeppUwCzc94Z8YC
4A7edHmlgnTM3puJTNRX6Nl6OHIVcnIWOGMng25a5pXt8KBsz0VQuDp7hWEvbkw9Mu+AMCQM5OGO
TcXNyibgYEBsT3ba6zzX9PYNuZjvothiN+17e3vu/+QheTSjeAPxHTBxQRh5YOCABd9FOaifrzfz
DgqtQ3X5DZ43YcDijd+HOtUD/xBeWI0Kk5XIuy2dli2n+ZYhijxYlOIezvqLWVN9LKZsYLQPLbP1
RDOBT/qAmD1VR9QNlEkz2c4PzL8o/LM6edL3Bx/6YqjT+nXAK7oWucIeHYL92MUfKENLrnQWXU5c
jqDZ3+naNC28J/LlVKOl78fqgSvJaZoeog6BBySzCHYR9dbqp2cmVYQmgsoKZ9/Fk9QwgStwxFlF
mWvWsMFu2s7xZosKG/9J3rswHNSaubxe45LiqFa4u9T5V6VXHyf+aj6hz/Jbjo3F2ijekaz4W9ZZ
UFMQoVNaO12chG7CTkf/7oH7cayaAsxFimRK24PmHbOYrIKoDwuJPGh/61lG6qjAsrbl9Ag/5tXy
b2eIGK5Oj2f+nCK409vW4kn+At5Kxj9Xjqbm8+5dN5sL2ZGV21OQE+AHmIQ3gyAq8KgaNQjdxCTe
Akch9wvSvlFUTHkG8YCrMwnqI0NP27aRJW9S4nICReWJRXHTojQ2zNnOl18/afbLA7UadeljPqCE
FxLdFJmDAo0gJMPH1orNzo0vuGlg/ic1wuaPkuZGH8rnRGcElNUJhsYRlfiobKe6P0TUBuxjw/wv
yb1n0cC7EhQWjsQnxboA0KiSgWmICNueCY4xa5498pnSuVymdb0rYcR6YJXXXs05MYcqfrdOR4Bk
Oa5wkwp4t5EKroDbdK6xd8HMPScV8bOmkAzqEMQfikv2rfrJdPLsjjIbocDhJvV9M1QRKR0ZzCom
vZcH0MpNE1HIul4x6WTlzW8QPJwZEkKEEEHUo8tw+uubXx6N2cXwwB8hLjU3Gayat+K3c7U2Mh1E
80ICnK9XXBSYvmUKsEhcj+mEYGNupwWV2aN8ok2J9yU//19k3io6ma/3IvQpHtC+14YVgIDexntK
CATMkUJdbSBwvTJYGTk3OoSLp1D3/7UWCaLvi9L6CqR6HHNwWvPwUMtL/Rk1q7D0/yPhOV3Is0yK
dkvBfCChJUcCB7OZ1TYeX+xtwzUtPZ1/9GkRes/hx/T+A5AW+s0WWy8YAa9R1TXLZ+3IOw9tBqZz
lb/ZMDSqWkCrAblxOyj7NYrMXClotwZYYd0cQe7NjttYYxkApGCFo2zvrRng4Ya9heeVc/e+KGsf
cPnrqDe/tVQ9q3UMvPmcyqOATPLhxUxt9+A2t9JRggpdlWyVEW0BF5z/YF63IKkAsDc6Zw7tz/us
hWA78+gl3/X/dS8BTopX0TzIpOFy8yprWtjdpPChzBOjl0BDvij6l3RnqTUyGKifWEx5HHKAsvhf
d9LVzOfl5UVw3G9Ngx3B3Wb9og0fgWkolu88JgrT7CxfAZAYsySl3eHKCRroQ6TdfhyLOGBc5WeK
buKZDLvKcZYxmUdHsSzrncQrz5BuQz+5GYZdA4FUImY9nEUr9hUf+V91szqKSu2ASTAvVMA5Pr2r
1erCil7/zKi9imcZGZcWnvvZFhLyypbLc3GLaU64CMitlVT0lSZNDZI/0sB7aOoe1kdDNOX3pbgl
Xe5wUU6qUvaXrIro/hyChM59IeGW957oHQd6FJhCSKzERV2FqmQg4p01LLOvRVC8xZqUcbXVERZN
l2rcBTfBOkYphK3ikkOdllLg+QoCJ6x6XMxSLAriklVTu4ZAd0rHVgwHGnjg4CiR91hx1G/6oaxL
rp70p4d0hghNwKt8+A2YUQSZqSF/RX9xrSz82SgfJxQ85uNV043GpPmHfuIgs2A5ydi1PJn+gHct
sn1eaOAvIadRTbbdtBwYcTEijsNMy5G/ss3poYLEW0XDNXbWlXCGejLHra3XQ+Nh/aGjSRzxNyDa
tImw3tnf5xqqnty/beLtM16ijQFby1t6eWzC+hNyUzNy2694LJNyNItA3b4Aor5+ivKccSB3WXRO
AIBxHShUJKDQZpjmfZvb6qrqIY1JaPfW1WIhDTYxjvIjQwRbJsqvCOgSCUJeAgkEeQg6FkvblmV7
5PLJo6cL0hgM7v4KOC3ZgJfPOuRkDMYwsC4NnyKon/L1IhrkvfDOE16q1n8XMGN7zyR/AyZe5e2C
BK7oQCpE6OMLdBEzXvikCZabwhJZImTZN2FceGmYZMOeP0rIft+N0RQ8Ceb0nIX8MFJ8NnrDtOo0
BgpJ0CZVM3vUqSxRSBjqlfFfmiY+cbAvQ8jinQSEzlXpW/jZCAHjtrBULeOfnx7dhczlV7B9+D6H
K/UtpoFKikhlSH2499ld18+b7VqYrhOiZ3fCg1uy1LGi+EZ1SkOR9GMlrs2+BP+5lEiZGypDyMxj
fF1JS3Aa+m/YBlV6N5Ol0ZXR+XC74MP27VfxhHFprVDmCrNLTS4sJ4+boDnkNXSZG2xZ79LJhKon
5C/HcW1Bp2eKq3P8QVJ7/ICfuCakI6Ldeqzt5Ima0Xz4RGonFtWRz+zm3XlDraUq3N79DsXDtzb8
9sNl0tmjsrQJjY5O/29oiA7q6Ya0Dyo3h/d4nXieGUT+k+aDBKBUGSNbXdRGSQMjdRRMaGmzBT8r
aRRWtXh0/YoxZlHEvNpijFcbFUgfYgqTZt25I1Vep8N/R+QPe/MJhPtcaMikg65zEif4PfTH5hY8
C/C3IiP/yS7m9BqzvByDtQ36+EQqU7aoAVxdq38qGDrDT8u1YbO9fEFyWZd+6sWQ7frto5bzY+Gv
dm/qernttzjlSaG+yt4BXTNxjF4nfhxExKzttq+a9mj2EVARE9aTwg+WzyRN+2PNJw2IinulY0cr
QOnLl+2Nf6G/I9ew9TA3iZ+n+zSFXPv20WhQ8Zm39lkOJzs9hY+0BoICert9KIeHDTOKMghrBILJ
79v3l8UZE2fu/MQW2JpOAhrM7xo5Y8L5SijU0Ub9fMUe8Qy91J39qLuhlonaD9u1Ke/hfsh0LIjA
ncfBpe9zCBsDbcZAZrWvRqGNnibe2Dz6SdOYOr4LoUfBvNiN8EQUpvwzjzdFhKcJXP0D/1Zq8G6d
8LsgUu0n/iofzS4YD+4CpjDqGHmDR1Jeu7X3wK20YD0srKXnnLYHousedp4f0TccE7r43CBcUTMl
vammV2Drpw0P3cfZhLiOIskY57AzpFSWLkNR+E3pE5dmH6r6qoOQfMRsCBBLp0bYBQDzpl6qFaGq
qdwSModeqID8+O30nn/lKpxSEtAn/+YMHk8byI3sUI0qB7PjayxwzSo/Hum0M1efL/KvbngvmKnB
rSEZCyckb40g9TbU3FcKkf7BFsDMP4wmEItnrQPDB2hNxJWIJC6rzWShxWnseKec0FVmVgzsXkxo
2jnn7zJUmY2LGJHttI0lJ2YVKKpDuByf9Nt7zOBYir7D1H7JqLnphUtVkpOPR6RDe97T1RcbZcn3
g29WVJwtzttLP2IN0Ip132AQsXWR/c+1lx3mgRLxb7M94QphO5Ja5+2BE1r6yT1+THNI5Iv0xwmT
Ru3JZbEOhUv0k4HNYH0zM+Y0u8i7RjVvjm93mmrTxUHG6RyA2HprH+gHLCc5rr+ergxc7InsAaif
INlbwzulYYbbftjP/1/VJ/9vlWtC76aUz/q9mKlz5RDKkTC/azhjT0hfZ7oysqcQQ+MlGh1AdOEE
McoABQNQHvaDZ/FIJH9UDYyBfV5Gn+fbTO5+BLTIPoB5jwsXWOoFqQt2lwvVahBSoT75OUeE5qBI
y1TgA2TXVPlfJEnl1zyfoCXktnMEnoI17ntS8c6QzykMZigHRrga4sXW8N/twQ8fyqBhMYvuymX2
HjzznMsISPo8VZxPRcMaXOjf7jKNXULJmn/rEbaqdIMNQXwShIPEernRLCuXPWPZDEPOYK8C2ul+
5dcVyiXurSqMeeKLNexcFr4Alg6aOLwiXTgGE8Xhr19t+4hNQq6p5uuXZ9PLB5jDZurHVPwVTjhO
tAdY2p4chhONCbLlTpjdIvLL4HL5fwb3q2YKqihxyoiAYzZL6/bNRAo9/ggceWOleulEjH/7oi0w
mF35PwqVEGpTpOPmVtGwV8ah+Sf/EmUMTyGQthcpgrsAESioj23/Dj4k22e5FO26iBB12dGLIHQk
JQLs+MRLrPDCsFp1YPu06LmVluGpPWF8+n8cl/Ap0VBAgI/L1z7n4XwD8GUIn5WjHkOR6BHJ9TKf
TMSGrP6APr0LEretgf+CHZBnoY3EuTVQUMbWhG5LTWhYUD931XC8nddebGgPf+9QAhT8Fi8m99C5
jfliHxEKwUpTEzpaQSlq8LQrbSBPkoCL/CeOCvcZpGtklEjodQygmDLfNOG1RhM3MLtMDfdz/L4L
kjJJPJLkCo5ASvGYnYe0zhCpvbh1Wy66uQblB4EIRT9B7oZQ9WOA2CCsC/ZstudZQ3FIxAi2mN4u
wkUQwXPIdgREkt2W5FLoC3Ibe0JbBptYBVCRe+UMVgBcM4oa9CncJ+2BTHoAVdCBH1qOGHV0S/eq
Y3s+GczIXP6INZJYYo5Ge2+IHUu5WFL6lLXFBB5jn0evGR9zhDw2CygBE+zfeZGjLxEszYJjAtWr
64GsQ26bscNHQytM43XcYq8mAJBYlvNqd6SLbrgcpUGajlTeNj62slQ9P/1FAPjyXDYnbncc4MN6
E5htcHnQDQg05+uJhaZrLvWmvKCuNb74rseiTEg1zPcWZ+cW3ibyq8qGoKOM1GNUhLTXIouPoNrt
ChslWFf9mFPCkz70d29HbDnivKTJu2nF1gmDARHUjdJBr7RU8vKtGlFMuTp1xM33z8FI7EuxYGsf
oKqPp+rNmR83o9wwIslDAq4vWS+qw0dpv6Sfh/LICeEoRlmhvUdQJt1J7Ldo3eyvp8jYhavQ0aUe
+5YTDe4cue+iXnrN0vXhjC/CFbMhG4DJJiMtC0U0RiYqMgeeRUPO6vMTDaU1oewfvAD5W801jsby
ee6Bw+A3zYOnlIXcIWtIq+DmnFEbMkv4Y9aHqPKxzo6QYtqtMo1r5FQelnGGdr1+iPbboD3JP1P4
24Lg3RwC+KEZYeYuKNYEM2fdf75bQRpxHsWDFSPAj+Ixzfvrz4kqm1bB6/haf2BV6v1Dv4uwWBtj
n50tNa13E+7yAZXN9hOW0JLlQyTSCo7pIFpoCamtRQOxs+b5Y4XeHBESv+We9hnE6uPc+xYRNVwD
Usen4HdzwfpJUAORsnkZuac7h1f9HCR43FnrzaCdz9t39tljQmLvGyi2TY1zx/YIRTej1M5NdMpn
8OlxBBlDhk5HQfPVFmCm6YGMf3p0BmdB5UuiqycUngpXiIEjAI8i57Vd9Gv31BfXZnsERRuv8/SI
KHy7HU62m+mfHveu/P7Z0oyB+Q++W32L+ZradTHCZDPExXThedUcQkU6rr96Cvy9NiRjA7v+vqMq
cnsrsx4kmYCkVzWtUDC6v3svEXXG7Izl1JDd4pJScA8sdU6lfBKWTjRgdRku1uMxDTxjD4lI33Pz
+KKdES/JJVJnH1Tu4c4ZMv4kmwOe8IlrUlg3SuIDltOEvX+UnQ69hzrm6hRxemhBYTLQWHubDFqZ
Rt1q3WiyMOGszYo3toyx8cwVl1oXU/WBh79Mj6Zo/P4wUCyMhLCdtUZJ5kLu3eZ6HJ8YYjqPoWHG
9cj/ya7PC95UC1k02oRzQb6a+u8wahCgGQ+CTY2TZjnDSrRXuoXUH7DsDndMGWI5smZ7puTFA/pA
FA7kUey0ZBeuJ8GO5aaYTxp9DgyB5yIY2kC6U9i2I6LLNvnMkLQkc+iSA6OHJXMpmdnnJjHJWivy
G/Ju+A9YV8itfcrXeTtjsMzF9C0O6nbMtVZWI8k7alYu6BbF19MOE9GOGP7vb30yRLTlm+kXczng
pgdSl+PFufPnceS/Fxlmt1hf+0ZO+TT3vGFtpGsbYwBTj38ZivZHHKJoCXiRf6rqWAtpvQFsfl8I
DZnF2+dAP+1Hq1lKv1V3kHovPiUlmTrZv9WXqCP46/Ynme5VFx0a1NoMgRpt3vmIDwP4/YhDULsk
iItFzTxbMGVcMCqFIJPuBOJAoIjL/KuIgdqdNfko0LYL3Ogqlw62T7V7ICpQay5bJaZugg9Fp8qS
mJmrVrtGKypCC87wPLV+jVCeHhVTreROiJl66/xnopfvFz/GZNdJlOVm3P0KaOh7WX2WX+OyBHTv
+fexKuKwf/Qrzj69xNWm72d1OoTaZ6EQcFQmumGF3w8AfWQradDmBearnBkCI5Nmz/Q7wrQOQ/bd
F3iueuQ29PK17W8R0fUHb13Nu2Np4+gd+sHuIaVfcKDJ6R4dYvil7SyvSh8dbzvPu1TdnqeKFnE6
abpJRRx69Djw/KA6HvKx6j+iQvPZN6JYrTbGXGQ1s7gVYYJ+9+pREsc9Mr0Pe1DVGSAIbbjioXp1
JOGVHLxV3Dq4OLeDU+n8C1nJRdpZ6BoSyOOJinQY+g70DudeVHnjjh7wusj7ym8q5/tYuZGZ7+w6
pdEwxvrVGRsl1q5V8DJ3BfAnaxaChc+7bg+uEjf2PT40dHJsRRa0MArApAFJMhRj4iGlNp4FgfRm
espBaJUH69iUNj8pul4DOH0aEZtl6oWnXK0beoapA/edxMM2Wpg7libyQ6X6AmDqn/rUXdTEdlNs
/chXaVRMA4/uUnaBNBOgVPyLXKRxic12guwUb6O8J0+0X8KkDmEhemITC37xhp9h0eu8ICrD3vhJ
vudSiMN+h7f0oyPwPKPF9DUrVfYckTdNCgo2vKaWTz2QOBJLaj8k5Xxk42U3LTWQA6cspGcUxJPp
N5/q+SlZ8k7vV7DhOW8XNv/N9xs2l6Yz8BN3tSMXHg2tINS62QwSpxDC7CccHRxjmA3JYB9YDiKU
7vBQ6QR8Hn5VNy/eI141WE8IAtMLo0mYNR/uxCn3H9BLpGNf0stbWNBqBCxdrNAbTULQbd3w3y0L
1CyrA5eYt6ndGngF+gxDh2SpTo5roWIx956cC6aemW3V1lhXiXjlZ37MErCqSKMBtglvI9XPCFPx
ec4KP3RfcmhjnhoFxiuc0rIwDgnZMuCZKH9LAxYDXHoCchJ100Z37Oo9vaYsuM9sTnYb10cHmXi3
Whr6eQRJE67l92S2ybVpxeq+zBDmprAyQb3p0bKp3NToSx07+r1hil3U2JT5D6/1pmzSiPC3Rh7O
pU8WVLchyTkLOkNtDD6aQW15EGSWUegTTOLvKJLCI10P0/Uvf5S8cN2Q9LpBsKA8TXK+NArNSzRq
P//tiT2G6Gg3uUxXcD+Rr6S1+onOYZx4pqiyfLCgOfF8Z21R+dRMf7u4WR/mI8A9R1TNzIO0OwPi
hbf/LxoGv3bHYsnw1hMKaxhipCrIgsqF4Uyxr2rE5V3QryJOTTQlMs3OIeshhSf4ON9dJOUmPA1s
TpERNyHIYCDrNQtFAgVe6KC7JrWpcqVlMv573KMwhcNowBhx95PwMYu84JhQEM12DDKP7C3s4NKB
0eSi9MnAQOFKpTBdXPkdJGwPprqSRr0QMBtbS3wsLV4GGGeBAw3rcsLQbyl5LuqYWmPAjsGKmivE
tcjaKzlFWesEgp63gVUOhJ1OmzolRmzlpDNKpvS0Rb4HzXsRmP+gFZ+eEomrzsGIt3fLiF3lw3D1
Q35LwkyFQcPH3YpszEcAeS1zZzdHwp8x0+kmGTTIGNqizrwisth5jJGylJVLlp54HOhtT1i3dSJk
2R8KaxR35JhFUnm3SReKBkpRU5YDurTGZaLjajQXl5c04erpMwxFngQ8EgX8iJ8YZVcp+xncaYwh
mR89YEgWsQm2E6V48zFZfDWVkkxvC7EI9uQLBvz6o7oF5KnGLi//rFguFgu+czytEGrmAtgEYw2B
mrVMAWLMQ3lZz8uJZT+1qdX0MFnPHkSQ8XcWoMg4LZoQBV3B7aD6lCKY4/tRnqX4c/asblbs+urv
w7hmDwJJktmYbKDLsaa+NF0fvinwPOmmHHxQjbXQpDEnUdeXZOlvH8sh+nl5qZe82li2UquO7nNT
xWv3md0+lMasEzqQeQC9BlLtWI+znu4FVYeYzD+ka8EGCBCHUTyS1vwY/R+NgaPqDx9uIqITqnvs
rr/E8XAF9QAjRrw61FR8Qd7cOWU0QN9jOuDM5QOxOf7HBa5iApAPumEJBWcDn8d3hb7unyyeroVL
1PGoD+arCgR7MS+tHXIBr37JV3VA5yILSxwurlOlqqkYHS1oFyF6g0pEhUtYGmcUaj6KXiq/dV3O
lSqdqxntfsJThBXzF33f+lK5WdH+z9uBl9m8udzsHOxIY3V+V23YEGX58LZLSL07IkJJzJ2wmhhj
FPF4q3N6g1W5PvBDewNRsluykJV9GYp4KsmebPR6cSkK1UUvybHZTHPvnkE6xf754y5D6epb0d4D
Oi7wSkpZMrCyCFHJOh7X2DmWzjONq/nY+UOdWA5B1qyp9scf7sYIgQMwMToEaoTCy8B2EXleklyU
bBdkoGyhiqPi+Y3wCBrErlL1iB+PgZ1YARtXjlQSgS4qmwkSJ54pvY6dO9zGwYVSDcWKPhnHzwgD
sYGc+IL3eSSnTw1Nhzx6WcCxAcxpCPlXE8faaE97z3H2ZGpsMb6r+JF/gevcFl1C8InZurZhv6RT
f0xin6UPR+OdXAifAykjKB/QmMYdjyLjghoH++qppaPY68c3UC+YF6bM4pDzW5OFSVmD6Q7XmJC2
hYA/b8eK8Atk6XvaUwDFvWKHTQ7aIJ5bMJ0WWkcUJqqcBt8r7oEvzU1AT+W6P06hRZpQoCqKqM7W
yaZpdRihc/PLx7qBgRuSd+NRgcbg4aSfqrlLj6m2DvKCSFWQuqdmNcekPxqNIuvfn9PR+xE9xtVa
xSCan34WQlCO/tvjbeT4FXpwMJe3s4Dhx+rS/K37RZx5n1NJGRNHJF2LV7HdHNmFhPQULQB28mTG
Gs5f5B1/R4GKic3ncRpmSZTuPTUPrk7kuT98KuCYDzsmybFXVAM+BLpZBbeghZO3lAKCQ5TP/dkd
dvQUFZ5ZVtShk0IjpGje9N6hr5kqBKFdbarU4sGYV4mbYsRSLoT3wQbrLA/2NXgXQDnME2nJAWpW
aUIjv5lxGKLx5r3LpwDzEzzZSo1QAw4bj7cXkM9+9aAXUEnGoygHE1GFZuuZUrHnVTR57qtjZ/oh
/j54qylrsBzL713bsQr81duMliYxt5gVX6MHqspN81VLOsR6HTnd7XP0YIBRjMkkylVPZm/NyXyr
5KGblaUgyGDvzg3lID6XRhqtYISfFdliBWe/pL1POlRHsbEZNDhDkMzaNFj/mDReabspyBjj5Q7b
9szHrSXs70uE1NSDGUtSMg/+NAcDOpkr10RAjoQ8Uye9QlliT3peu/YMgG49cwnhk7UbgvxyB9Xl
aQbJaRZutC8yHW1M8RTl/4UidvwTcD7WpGA9qz5hL4dF7VKjlz64GXu9MuKUjVJ/H6Sd7seyqPBY
+wpstoQO3v4TLkawm9xcYtmUkSbDOBrWMXJxb8tSIn6BqRIxtcjhV84DnT/yYaQa65PBKCg/yvD3
q7hGShFKJLSsISeaIh5Bc7rhOXim2saJaW08gG/Z6aHQqriDg5bbA/KKR7BDXfjXbVGso067fQzg
1p/mdSQfUpxrW3QutHevk4ZrFVFqMwPZDOT7OnvOTBieZIouZm7/oxnWMsmoymG4otpAAdcDticc
0djSd/o6/irOkP7vdUjRMEYYtWVJkRGbnhLVC7ddS2YiWVcaEPoRYx1ncQrh5nrPblKcWLu8uLA4
zd6enngQBNknh7xqoXKFmSVO6bfE2VTxscLKSI7nWhcDUdYEyFKnr3Gau5EkRf/0kduLID4KJjZF
fN//hbvl/0oPWY7LsYjPh9YKwA3grXv7VNgVOubnimtQDJRgIbHOSzWrsQlC0YC6LvVA7afOzCWH
cKUTOCaJm4py5FECMzvSntYgjM3o/MgOlJTsmyPR8cSWtwr3dleiSwYxSbDBk84TaWhMcrynYHh+
xNgZsZh6IkZrjugTw4qMyHTt2ZWZlk+ymD7oqKIKXSFnzsRORBtrWJyE26qmMEWF7kTQfQSBO9qD
Ia2WxUF6wtmqk+vIeunznstrz6S7YqlniiiGk7aJK371VYsMjdH7qZO053oa9c7jFcqJYJr7jN06
chHQB3obXJ4IwFvzKq7eYOzLaanXgnKJr738jZdpxwMTF7HqckKrcFJxdjnd6cnMjjPOF92GdeED
WBR6m2EgY5xHZx1Yei1XB3X4VVRvlj51DwMjZixglHHxZeYuwW82xkqdkGD96IFLsQ+VwqRCzw4o
EBg8xuNgdoFJQ4xUSkIbvxHMAZaRO2spd8XW8VGvBgD59poG/BS0feeUwoxWOdaGVqIE3QWggnlj
0bKuG65kBtFjeEYbHN+jO6ufvjxLH5Q4mW7jBLe5nGP91z9wkJTJ/Xyk2Vp+96UUJh0iH2ATyGJg
WVh+EeK0hiczmMbxAU7a3Y5oX77tbtVqOumfH4fceCln1UPLaNiCEeO3CGRUG0SAd2MKOc4RVXF8
vR1xIvSMnSDG0kjIPL6Bb53ZWJDPRrGtd8Pvu+S3vAP/pW3H2E57cr2R/ROS0zCsxybGzF7Juj6l
laq3q/35lZw/co9GD0zzeGi4v8lBA1u9XIzq9Z4he7HaYzfgTShVekG2veb2z/BMYI5yZHW9mTJ/
J+LP+BeXHLtwbk6O/enaegqI1XJ3A6IABHCSKZi/2Xvr4lc8bONR+70BgOSPia86kD3ov163YvYB
8XGqZfc/Msdw3Li+F2R/XpuojqBMZSQyvBloGKI+ORZm3nNJbKTooxsFDeUqWvrqymYy7LtDtlty
KrKE+qXLdzm2idpod2/wkO1GQWqnTLZgGjamFt8UE2kEaBB1+S1TKFc+uIKZXOWS/zaRATlYvCm9
eOfbJyaRRwNISzmXYa9uy6Wv9mOJAfxlfKfRYG8y6JHBrO73+Ov9Cl0wtemjWjGAElzftXaFin88
kfI0ijqtE4OKdcneg3Us8316LsdMbLn0wbqh38DC+SLQQx9RsBkUswWENTzkcFhQuEuBhFQR30pg
tqro2BgxAww1rSWBukCwg+3ujs1d0ywrhAxVago2mFQCvgNUA7OIG+X78DZVfaOPVraIU7ahArHF
QooI4bJ3ZDK597CMP8YDD76xjG3KygrzGQ2v2zxujye+T30DmC6XL04/IfITZ4DSphEWxkqaIA50
OkCrE3eZSQ1Kk1kUCU0sSMtFarABugWvWdHSiKgSY72s3HGOUqFLtH1YROs0DL/tVb+Z0LPhKXh4
fAAZSLxBwIVM/oaFVuP/i714hqTzYztKKLbDrAMe9QH2/0XCgCO9z+je8X7Mrzgcy7crwYkgBOOl
sA3ZJoi0vnVDlQg6+6WS64+6+2FxQRpLMS/KgEvf8u7bu2P4YMF1xpyrd1EoG/32TpmG8Hqgti5a
U5cpfwlfNVYXy+QJm88CwyJSV6Dw4K0frNXjZxdGeIU9EsSFiEL5Esi+3+XIzRHCdwmTvilRUPtZ
UOIzZ6gR8XMSUyxk2VOhNTDm3/uOmmgB8m2S7s2yJB1OVQdamROhLe9mc/EXMeFroMQKh1KhSsB7
j4vIIw7028F55tFxXq5KuHOEYC2bsoztj3/7yEGSwdivKDpwLhGextt2x6qYNUTYSQxD8wTe+gzc
yXlU4HDwX/cexR7y3FrSeE7CXL27raqonZvVUx0+0lDEjKfl9df+HABU3aDBcqh/5IDl3fbgWau0
VxBXYdxHWFff3biE9pDj59raMQtRNNcfaRhZpD/stjUeuD793Hhq4Q6M/aoM4xnNsNAKnd7suf11
JwHU3tU3TR5oC4OjA0h6bTaGjYuGsBZiO5Iczg+tNw9iRYT9lEwKp4mD8BX1CEuJbAoVDUBLnjlO
yjJmjeP5nLV3T/gwambLqOMCsYb/Fxmv0eFiBYyxEggmIAbpe/bEyzP0mTa+HaWt6kP9WwJ63U/b
bvxgbRn1BuS7J/KhN46s7axomurnu1oHa4xcGUU33TrB8s0TFzbXZajUVeEp06rm9wKn9Z3tzvQm
JHvdvQe7/bPkWPoUO0vOREAn2MGRB+LIvzqs+NKwTueYjONATzrAjJN2YrbTC9Az/Lq/j1TcRQrV
rZul+VbFw+OiqZypo7fwCxCmRfU3xP2w45WqZjol9uQ2ZOod5KATAtaWusjDV0c86OZQVlUKH5hx
EF/YsWWsDvByJXeEd+xyzzp2Lbj4s4M9KLWLUQ0QDcvIFmMzODFMdhFG4qM1Q3GQaY3/RmzbS+6m
HvdPl6B4mKBh/mevHchLaqN9RbHjaB9grtLHSJpiZIlfAc64Q4uwPb3tcdTRBDCOR/V2ELoJBPFa
1rrDeI2G4gaHQgAsRZ4wiILXcT016M+5wheXdV+obnvwcnf0gJMYYgDGQ0PKSumahMFRVzZhUAvD
0dXYodsnWWHP4VrCPn6xc8arIJUSsX2zyoQuaymxyRcJWIy1tUvqBKyJh3k1Jo/HgeAoXYJ8T3GA
NohBXRFTYdJeGBFEoiuo0gOHdjx/Bw5R6oGx6B+YgnD2JRo22HPa7M58eX418nnXPzR+NbDe2APH
H5GhMPi79Ch7W8Xqbf50DeO+SR6u/MS2s595Y0XCdeJiSEl38TjDIUTjWkeo4eX1c2nIXPcuml6A
XRTCyVc4GtncOGKotAYHg35h3fno8f7v1fVwaG+D+2/1+xSiJP++FvjbMkdJqumJyIeU4OFQ9ewM
hY3kP4tE8E41it+IbKauKNY6hMavkSQz+Ydunp1J2Y1Gqeq02APR/z92n1yNzTArF3A9VF0XvCLw
LAeYX42YvDYMbEF03CedhpLTRt0NnIsoiw8PNXsrIBP2dmsJTlO01weriwrXiipA7RAN2SbUA53r
nB073PTWspPz0e4BfKFuQBKKcNiw5Y0F7trC0TtBFJFhZXI89lVBHegmgPeYJLKFQpENzjork5vt
sQrDcg+hHo5OSVN47gXiBqE5T8nGexmGZZb0dMT0fgca944GQC/iOkxCC5/uK0MZMrussaBA+LiB
B1AF+2n75QCzT0ZgzZ391/NBCeSA/R9b6lKyYq0oLzbNpxl4igZoXPkbaDU14cHtQU6nnp9h32N2
dKQW/HSoQA0i+h9/IoX+FSfpP5aqY+Isfo+l0jZXlka66rm3zRLXDBjLrMRjHMVizfr6UN7GtBNd
6sq0iOOvRP8bc5t0SXSxQ0UKC69av8sQRJsjiopLtvMYQxTatZ/GqbhE7SBVTgStmMKb3/cGoehb
BBIcxaooG5Jp3j9uo/Rtii/B3Tonp2OvEchMrm1RH9ssUDD6+JeaprN5BO44x9R9kYqwRDNxgLPW
GqhRoEwprrcX2eYmrE/QC6unujMGHnUXqVy6c65b4Y9ewqrLJxj2D0XB64qAQVdwPmKDStvhhKmr
SelU4TM4+LVs/80yinbzjy/FgLcGtUa9Dorfe97g5uJi7tuyp4uawoaiTZu49vNlUMmLngNcpWuS
iQ7SDZ7mJykabc3JsEsVL470XZsZRDSgQRP7Fk55qowhzXT6D1FNaVwtQZEU3bRgnaGGXWhLcUua
rDcphTaMyI7T4fBqs/P1/IARXqvAlD/aQdL8LqyJL9YOhsoQX6ozqfEmFPcVGoIdoOJxQVz9mj/9
FfWxow8a/v9FiUuG/bBjBArZbRk3qbTZZqhqo8J+fo4C4exy0LEmJYgaQeFbhVUw5Etl13KH4ZJj
NzwHh8tNJUEUQvQLoBhADzxUfa2qyq5bQB7t8sk6l2DI2vtI0/moF4iL04eU8nityUU5vOVyitLo
D5Y1V2z3SITzALMIKyANXSt1/nONBhuS+S9StuVcFiWd3JqbmNN8HbBxQpjaXkkfAGtzG3osJ9zf
1aw5X+nGMF+mv1dX9KZ6kzsq3P1k9ksm89peHhRBhT7IqEM6E8rdEhZVDtkzgr8ZRSDk4lh8abAj
cHK7xFVf+e3QNtJE1o/7cuBbA4339gHlj1CvFpWMDd0xgcDxycycacYAuf6+P4b5antEEZ+KWdwT
3EvIAcG+fWe1fAh7gOYxA4DiJQC1SleqbtAlrCV+NcJX/WRANWFqLbUUtxgfyLCeDXLA6n0iXYcp
+8aWlLaPM7erVvE1NnWYnP356hMIshv1rDTu4BinYDNZI9b2r7Yf1holDfJsXTfIzwoE0S5oW281
q2OntmCt0pV20xhI+8NLItGL7QFraVYWtIS53yb9AIDnsHjfuprS4LQuZmENBPEf08e5/qLISqez
/IzgJ88HTmZYjhheWMbyA7fuVfR/CpVL+gmIPsd7k+3dRGo6nqF3uU1u9ZmBd+xHwGgG4Uh28y4f
JaGeIk2dtmWcMo1AvaUf/v7GtHDJDAQZhedFgAaV1w34tlRpDMX2MI97CvsPnbo+v3XG7HuE2qQX
9jE/pyuLKvqlBrBXb3UT3OExBEKuxrWoYsxTgRQkTJvqzuN66GSquEvpfq5Hlq1kQ14IYN80fIXq
V3ryRF0pbQSgtzTCXlfj8PyMZn3KNovX+hsqUiA2lsmSY+rVuyZC/4cTj9zwnbxyo6OtcqE66Y/a
wRfFZ4/DKTctGF+0zVSXjehiGoksRkrplVQddO8lbDkd6qHG1UpL9Ss3Tq5ntwfSTCK3KYd2j+sq
NhkI5ww9zAiCnZg2ncu1jWIm8ij6VufGXnhWThFnRfEkTQV3yb2pTFo1ldTgxpo9NW4g6Qa3TAGi
BA7cwtWAcgFB8nzyfQEqM8yty2LGOWScifebue4lTL6nz7+BfFURpW5UHmy0nUbIPqtg3oWzi3/l
KbgPoL3+K+fyJlL2nSUcAES0zv6MSdMVEW/DFrGc970mNvhPu55L71HdyHvjz4OOI3cktQHtYJDN
zg3cBZOLwTSqxEIAcMNW1aTM91pRx1I8Pkd0IETYdS4/57MLlhDet7G9UTowDKoGBvjrzqsWs60f
46ISjhC+fDXbF0TkZLdBmEleEUULmSHCLILzixQgafBLfd9gUZsuQNtglOnxJRjI33GHCNd33qNx
/HgaoELlPyizhh14Hpr9lfh4GCoxnhvvIvn8iXNA5w7yb9dlKVeid6O4/TV3ZctniGNh3LCVqskg
da+glluzN3+MjZxiqj8kLmT8jBEQAAP0Q+pdsVWPVf8meKgboPx4UsVdfpUj8OhcL6rT9001Os9k
E7/94PzVxB/9DJlWh7RuPSWa4D5VHjKE0F03JvfeE4ZufobHxDekgeDFgtL+6cbeSEIVMX/p4c8t
MTBx7pdgXhj6PNv0cYnQzA2R/1FgjUVJcpdfOS2PlaYu/+t66iVeEddFBHQFhdG3F1OrG3u6FNUe
Mqh8kWInlWb/PLxW+agDEQNNRG+oJ58Ed8fucCM9DKQ9ESHqgQGl7kDz6PXlWOZTk+fnJzCtEiDL
G0JCEu+pWIffNhnpAtxInUFrJUMV5HI8oAedgRa7H1emlvfv2TqR5BkFuGb781VcqysGYHuSfZil
v5LE7eoAhdUKNoB0se+2khXMsjY0U3dbXlJf/2qTV8P58h9C/GhWNiI5Uuscc+tO4t0rekTU2ntl
adqP/pD21sAiiZPWsfl9aX8j/+mJukxw8nUvBztkTeHYggM6eBV+4rXIBsXJnl3bX+UVmukfrMz5
j/Hw0es1gvF/CpLxfEFVCDhVR59K6rbVcyTf6n/sqSYSUtRc8sT/VMDGBvZrIhf281O0wl8q9AkM
1nbKU29AvJsEdtz6ldx/3B/5AvX9c7Io4DgrglaNZ7bx66G/UGjGK8j5R8HdxipyuZsZWsPMIaup
VQFDi8l6DLeTeGgozxDO65etIa4dVwx21iSUMfatvGUSsIjirr0nXBp3OySq6LEsWUc8wFd/YtN5
KY+OmrYW2Ad5NttnSMS4e0xh7P0Fu96YPX8tQWPr2unFpyfwRjEsdAtkxyWriqyaa7ppEwvBfT/z
QU0Po5OAI/S/Wr4qajzgqrKOmbmBuzqmPGHVamZpjiZdqlxHWh4eUj/Y6UVQ6Ktcm8vm9QQE3c9x
JjEXwJDR2UkRBPsZyGsg5nQqj0A271QXYc98fZ9NWAZE1Noz8h0JfgP2k95Z/ev397BNIA5ixW1y
/QhdsZ4BePuLLvcIMkKmUT57Wj6aJcIGKoSMt4c8WHnVjZh40PvN5G4qe0cZYHtuCA0LaZ+grmkQ
CWmeuy9UeSIr4ZNSZCsqD1USY1cKXwj0t51V5wdZl8tcBZyBVC2G5vWcCTJLlnEgZg63Yjs4B+2n
rpMIO1jrrY1Aq4drQNQIN9zUwL+z/4LE+kAmP6Pp6nU8Hv7l71ifNIKgAJICKsbmonpZYQFb7v70
JJGtyhYSeJEML/rXY3aBKuHVDSNR24ESNSYTy6L9BpdQ2VL9JYqTvW0X/yYVyIs1CNcwlH0PmMdD
tTx3e49HmA1UBVr4keLPcsu7kDPGQprsQld1Rq7kmiiNyZLcAuTminmZQlIcERk+z/9pKRyUWkxm
3XgiPAbvpZvjz79R07MqkSKnuezIoUvYN7CyZMKRSPh6qauFY6cq7noD7WoN83yNaRkr2g06oo7J
KAIle8PuSAIYtUhrAlxzCn4nAclUYLdA0ZF1uOOOV4sFXT3ChzMSC1DmWOBlVlNSoxiJ2SYpppaQ
muOzaSNkEFDX3TTVHN/mU8dKHCsUA0IACgqM6dspSt7hpip7h1ZwtA+MsMgwuf43Mw9KtChJqnqn
aqmCnkyumdzhWojN+WsBKk5Ed9fIwKUYQueLPFxQRx8UC8jiD0NWk4hyNKg2UfggPUOIbtxRnjIi
r41X3rGLUTa9ViJWT3RNk6HRYEvUp8wMYO1B7fu0PP9vo5kKVWV4dZSAsY1yF6o1kXXwHiaHSZrm
D8T76VW6c/HRswpZ4Ts48je/T1gnr8w8MtWecvjYd4NnmZUQ40axG9VIwtFAUOGDnwLTevpe2Qzj
DvO7V0jdOg/XGTrRdfXuLCNhoPQISVS2vbMVVOFx2GMQeu7tZYiSrVFm5Qb1wdkrO5Mj9A/Xhfn8
63Ney5ImlVBFv/0JdVsVtoCVz+K8zHxaAv26/4gRgMs4UrPLCwHH3PQllcZldmSXXor+uOGVa2wP
SbOI1IUrHIfEBYMC8ibzbDcXz4NF+kHy/5L0VWdf9l/g6x5xKlRgeVOmkfjXJ/drrtSrD4aNlNT0
hm7nMpbS8V6QI/m4CluYRFWlbX+GpDbQSlJ6Kpj51mDKla9cJQ1pcDq5/z52PAihsTuP2t8th5tx
ei4miC5tdlCKhiA4vR7AuWpI9UG6LqQKf9q4qc5MM7w6XOrZ94VFGxPg/E6yFbiVnquDoWd04fRM
3UFFAZKoIyoXSwegglYkCHFW78UxW4jdLMuS76vfqU+9oa7N4RCw+u79bdoV5vDtcaXsTW8U4QhU
KqozMoxMYWcxzkeKlwVKLRngjAIDd8BMNHEt9uqaYrMct5Y5PTckVpmW+qHoVy7xh1JLdoNa57kq
XTx/a07wuvm1AcFxnk9LHuta3i4BNBXJrJ7RkWO9+KKozuoePVnxB0e8/eLwinIZZU45ysr1132J
ozfWP8z2olAAWg+mw7/yXlur8lAtCa06O7dgOrzlQgVTBkQl+TcXC1SPYLvFIN9nr2sgAqKqnREW
ENywbd9zgulP3Am1ZQRERH8Wa0l4aBl001sOBBGqR8FQ+8Ke9oCX5q5QeFR0miCDbM4pDbcs5nMb
kgsH5Y5hx34um61IqJfcD5TuG51NZ2TzYQ+zaWjQsJQcg09H90aDV370K6GeYQqYKz3zaewWurG3
ubFMNfDMS30gf04QO28Pv3JBstuJ0Aqafbhkp4qPt6R/Yln+p33cU1zEu25CJ+o/+tqhUP7Zupbx
M7JbX1nSOwQoPiNsTUhz8NAVwqH3S5vfh0ZqQc3vEnW04UGzyO/Qp09P2sArsDeuyKC2PpQtKqi2
XAP9B+YfzQf+IR5mKKlIHt/PV0hbsBTCEltH93CJuULAA5F/B0fHdkn7cisNbZATIu5iEd4XSFsW
jYAbcZMLppgcsK4lGYeTBmDfZb11QTI3eO4K/DRkofbLstho/pw6cFoa8uGwEtjmJBFaL0M5EJBl
ZdHOL493+MBEfyFtrrMcrf1V84nQU0qapzd+T8wI7sCbuvLmkmMMScCRY7wn9eXROvrSUSkG7y1z
seazIapcRBm8br+bR4vKVURXx6mjzqlVrYhELs7HGi73MBXuLbxtT0kpMwznCTSjJWY8bBlsTycm
5NmgQHJds70wycDxO/X4k9eYXhIbrAk1MBIHA2jWhiSq5Uo+3w684gMCT/MszMBFuHVcaVgWhB57
/KdxLVI4xP8Ht2azu8IXTXFz0nCHU/4Fzfi2hBH/s9HIq3Uh4LUt0Q6v7kFr4vharXGePfge64h2
8MBxSEwEWHJXnHnqRJawfaUvFP+8bz6lp9hwzlkPS0hMgjPx69aATWXVoeKqHHGj9443HsuGawsk
VxDDOciBm3m2wVbd1ybe8kuTxIuos5QHtewDl9z03kZ45B+DL3GpEbZ8QRWc/JCUF6/Ug9pvbtkZ
q1n75+SY+iXj/Jw7iYfXApkDhTPv3NdiORXST4bapVCIuOkZblL9PiDF0zWQxtPd/3ZNTzltJSBM
EKWltfSn2q/MqXeZKLzyNteOq4t8C8K2X6ZOqdNFRVSnirtCOpmLA9epEiopD/tHqglfW2dHWWxY
k0sp9jQFXW1WuW6x+KtpJCS1Foy4+bCxJ+DEEtX8caxIWWaNdtyXITXyrEH415Dwc9uXlaA2ps2z
CXK2bZfbeOdI2yKERlB4AMnXFLa+XBfqzkljTYN+8usNh6PiQJa6RicueBfmMdJwjKZ1rF+SHYgC
1Xn4JhUpqTlY77fhGeS301qDsvMEM7vFY2479KW7sk6ZFtyaTqHRjtCCSxNznRDOrVIvKPckaBRT
5Nxb9rlEIZP7ruJ6Lu4ixABeX5UbzubD5VGePCxfuK1V9SFeIPqyvvivJrs6oCxDUxa4tKJ/qmKQ
YNf+trNLScLJo96lZ00yUu82Xb4nMQlaFP0NKFY6GjpvtRieWFyOVPXAYt4Xx9N2PEtbHXRx7Iv9
q0X0cpRZknhMgSVcuqUxvo45gJwDJpt3uUXzWybZtf2C3hZxof9Q2UKg19Hf75gpKwXsl0MNpEuE
A0zEMJjApqAxbruM1Iiq466IJqzmLwuSqsi7KCtIk2RlP/oTfXuErVxRedQYyTnWpLwqyRz5Nn63
1U9ltYLiLCUa+wlPpHvOsBBET7P4Ktjj0oCv8aINgCTLIT4YN593z3oRfZo+Ol1oKNx8JRm3IZ6o
/ZeIa3nadqlNOxuVdDoA6ATNvKnhzo/McggH6ATXYkE3EUvABOHLao4Kox8iaEOKNCZe21ffwswm
P1OQJyymSe+YTPbLj2LE4ImavYh4eJLY7AsQbIoyO34AOhh+EIFC0nYCkR3nOz6kxkijYPVoooF2
XQJlDQ1oFH6PAOCUT1JtQDZ2vkO0oyoU1EGcyjGzc1iweohinrFIPp2INLs1+1lF+kwBS1hCj2iP
2seVOKYKVFtxlr2ePuWZqlC5UUHu+0DnuSot5uJffugig6IrkeU1zTAao3gDKRvoxhMgpvNLe67w
zZy1LodFtzNAElOx4t+t4EQR3FdJjh9KRIXwG/WKQvxCWEj0yH2eWYPoGsFzkQ4Fihg5AbsmAhkS
roZBHwMgiK/uHiFtzasy10rp7yw5R1LrpEtVPJUi7NZ2ZS9ZF9qCtvfpJs3uTKSJ+ke3bY8yrMK5
tf5L8oWApu07VXIi6/eVQZphRUs2FNgQmjK0AReYcWoCMJocuZ4TSEiAwMBz2ZHgTSAteVaQM9KK
uKMyKppWj6wtliz1xxSsboyODFabhpjF1+C5qJ57gFrQ0YzTvZ7AEoCEsqYfAPK3QWWZg7LGiiZb
DJkAtYrmjHRJqA0c9x37XOfUwMysvspuBmgcOrORHBux3ZKhF46GrjV0edWwJYpxJLpHyuo9ZKVp
pkGtO9xl+05OV/PNN8LCwjBaLSGQ6l8RPCRPN5QtQ6khjRhdbASIMpWHn+ogfvGswBpyIs1LVK3q
GTmFz9wwO+FIH2HEjSI3dlc++9VOzT9pJt+ZY5+POM9E4zDl2Vjv2K1v1daLLkPKLEBssbi3aSPJ
kKHrtG8DoMhSZASSoNVzb7TuczLa2QdEDgzGY2ilVpVPW4MhXmAQ7D7VNcN5Mp3b9nQNqAcB0a3M
Z2X2bHegNgqudi2+zrZAWPb39Fwk6zzGOvTIz5RXWlN5KL2o7svJrzgI0Xnj8NIIs1ysUjWd9kaz
PgN9WcefgRG5UIiftiZ3pyqzTtLLeuUH///YtNE6OYvuc6h/jFL9ReeOLB3ssCEBDUUI9eU0LBl5
Z8++tKVUyIwdaSQpmABBfwkQP+dotoHjFY+8bx7X329STW0VTsQJnyfALuiWq2M4ANcrXrXaIa6J
VMr6cGHKofBPqIWPOm/WYPVdxeT8b1MRrsefE7eQh+gOLpMVZxgf7U7URH/KBmJODa4MuinOa2S5
1EzE7YCTMLAWrNi5bMGNcRBqUMa9RLyFpWjaBsppFvwA9LqBDpsQgqJQ2lO4RVva6je1T1aquYuk
Dnyyig+UFElAT22v1WwdadW0VCRObf2J9aKMw5QQw+X9gug8xTtpanhP0TR++tQA3gWw9CQKkkfS
7h9s7U9V32tYzt+eelzIujImUibMfPlzQJFHcQaU23xPSHQ3KGNiUg/rk3z61Fq3HVU++FIo0T+I
p2gCovdbNyeJXjOtFirTzym8b/hQM+IHgsWZBcigxwxRdKmafHCOofGN2qTXnI4bMZU0H2ARSS3w
+81NHT79GF7gcj5QB7rodbgwClAThIzxvdKoHEePOoxxbsSYVqMnRy7SytmJincOciSi6fMFLfoK
3jyYsfILuctXQQfNa6c2kWQU4KL+PIzzvbRVx4hCpnYlI01G5QcwgVCpp3iHWnDIiMUhowmdtuyg
mUczIhCb8hPX5uma5ZSZ4bifhK2ZJqlYnI64gCe3TQqDLgR0dY9e3SwKviO5BWgkK7iPZn7Hej03
qaGZk37/fNNlAy0QHbwfkUYy2jTz4ElgkLEqOSnmX4mjrSoVUIpXznr2jGoS7GeLUwv5FceAkUOX
eKK9Qeb+gzezt13XnnOYhRWSjVAOCywwrtTArCIvWgu0X7h83qHFV7YB9CNo5fG4COAftYDvS5I+
TKrdGAkG56quVgZThGCrY+hAdE9E57bZkGetk5SmrKa1ylfA8aB852WJp0D0b9WMJkUNfnWWtQBA
V/t2fTUdRhNn+LRLBD5WqbBPpawfdSjxdI2CA+X85cK7FUFd/AGQkFbVLMjGpfnxyIXShXw+ZH8l
3faDo9atA60+1Zccm2CzbzzMpL1XBIla+WJB4wnECVc3bPSMe4TZaUeibJqCzWrSyAHwLCQS/Kmc
jDC7i6uu0p4NS5rmx3hg6Wrrpd7TOy0c7D7+z0BHwIwI9l8rBu33HLSmUVnhwoIBBsKQqttV29+H
5L1qDwUxdVoAbCwBDSOBV4vnIxtJoUFYoUOZ/QEDp9dxnW4Fd1vVvnFSdjKV2EcBfTCVA4njz0R0
54mrhzP5mfc/LRw47jhJFZ/6eWDcUWdpVnfNClDv0HvIfQYZp8I6LGwPHZrh2mgkGkhkRYycGr6+
rAha7ZGNq7AVnZ9z7s+1UQc8EN66msITShvH8CBKVveIyM+K3gZN13kLNRY0DtzKyBrJCCdfKFEU
dZdN1Jh/UBZ+GoEiwlijSdovm6YsoG8jMBd+9s8LUOJIrGckLY2CiiUOmhk5gXFnoQwRg22HGlt2
HN8rzAWawJcOkrG51KpYcWPeTkXOGbQB/3srxuBCh9EVkNWF62gghL6/mbj07solE+K84qZhSHKO
qOc/wmDPNG6E4a1LnnM5eRFUv1WuAyvrtyVlo7ki1ClrrPtZgZM8O0cAPtkwc2b+hWbIoalQ79H9
32fSgaWftI+qFN2QHcrYSBb/TGIUBmWOjyjFmYBBiyj1Gn2V9hvr2n6Xu0pIt36RpaYKUucJXObV
GPRXfEKN3CrJvLnLaodpOImWnrqnWBo2FtGyDor05k4vP0W3aSPwsadhNS0G4epxp24QTlv8JU2E
eAd/5PlYH1y2oqmTThpj0fVZ5usSCK491Srx4T7MxIqbaDVU54c79aeWWKlQFGK75mRcvfXQSDCX
VbwkvXXTv5BKZtD3Dh4v7i0tO+7PtQfjd/HLWbN1mT7dbqTVf3jn0/tPZFyxK2g7GmcgMlyUOsox
bGeV8bDi1ldNEnbFNTz11dHnugiRzzwZ0pYWzXNycjGGCoy7VsamGgEcZuTpJ4Vrr03bZURZR7Zu
bNAbUutMkH5Koj6gpPhH8rG3dQECmNc8LXJlPVrc73qauVfAYLtacI5wOmfGBMxdrWfzYUBM0LTm
K4m9qMhKzYMOifEykj+tQQK2DzhKIa8uXT1f++eleBWRz6fa6e9oohqyiMYGk9yItr7lHiDkNd2P
jH9sYjhiWYKBlGobxnU9kWnZ3TQbcRTf+PfJ7uFzfifzFBf2XIB4SpmDm7fV5DH5pPpIPbEXM6hY
wfTkddB6qhwdQIaQcq0wvc3pL/DKyDT7b+bQlnab96RmVBLjYJTTqtLx8D8pv4miZfyhmcsDKcJy
vJw4GIfPtSHLFUeRR9kkb+CAzJmvjRfxWE37vHfhlhI+pBMl7unQBvg2Fiy36/rnQg9pH1lQFTd1
paqZSvKdb8B4rVdHy2l/U0yR/azYVGWUbG9siwMHR8DFF+/fpe12qFpt1AIRghTsSN8YFvjALNfP
Bl5eQxKXe9J9IMqRD1poc+1Zh8gVVsYGQYXqGrMBLwAaMlz1lE/DnYYYst68EtIc5DApRCXp7urL
vYGQpgDUM5mP4ehbehJpNxkdTPwlKm1tNyWgPwqBMS07bCdXsmh+R35JfqyJu+4+wCEo0Em5qMsY
3n5I+29fvUu4cjUBvhhdGlt9mWno5cbSXu7KSXWEnnWhTpVq0E+Csw19lYkGfznTl5/+TNTjx89o
3kPm4KBIheVUFUaFjAHcHvSuRPRAYnqlE9EGqoABL6+c+AxvoPRRAeSShSVtZ1suEdwSGaHpKFji
j0na4JunGumlU3d+hKWLwcMOd5CyetVxVrJQ6v4nTDpCN896DVrInewIAE3lHLqiEXRmx9GzEouh
/uR9JO7nomTlZRJp6V4XU4rpqqWCcxqBaFB3+ErQe5WEVch3SF06jkKlFXtrL62fLJrxDARnUDT4
p8uoPNvdZ79tAowIpZrK3qUo5JEBQX2vlW54ZeqOpSedZaB8r5X59mHrv5cnwPU68hk4QA8DwIwM
9U7IrmOkN4pKPqyY85ywYFf950THE1mwJh1XF1sl10rCl6bfagobx39UHOq7MlcnBMQnsYMO7daG
fJsp3vS8ztbx1m8E73cVSj6wCdWNKukmO/3HXxOkQ3JsaA6i4xUxQQnvJoPiVEcLk2pLd9p6hYjD
+jRKgQJX3nQ8ZanwMm+XUYN15wP2pfdykCYh5zb5WYwvLOtyZwaNj8UUiaoMSA4KrwaZQEY8uIln
AVkKrNkzTbfh1mzZpzIYKuqtkBIYecZ+KZiZk4z0k4QEkuJ5+pb8mLnx6R33uq35pXjRoT5mzKWm
wR1OCnHf1fE+/epvk0dHEA5NoUMVITPXVn4ITzYxuSfUhK4QuXChNu9bES5B1E4DyZlz2qLcVxJ6
CvS+/gmXvB900+Nmcz2MZbwjNoosx37JT8RShGd7LzoqlZVP0CtfLz3RsOpauurUgAl4Jn8HF8I9
C6Uj7x+m3QrinGoJkrYiDx8pDbEWppthbEU9+mmNrXrxIup+QAVNg4ZzdDgN4CXCQs2LXJJO14Ls
tsUGtWEcAqcQxkcYbJX4xAxS/sHBetwu2mycz4gbCjUQGKxm3H0XX8FP2DLCStetLs0UygUJln6n
2KoMTOya6pjXV74tDlNarg9ZHMlsSrAWFXdyoqYN1pAcqLXbMyC4PEj3J60dWlI9ueQqAIa7j14x
FRNIpfJHFFNdirz8vpKQnCT9c6kt+oFmiqexX4C7sn0hZrLFnEi8jZ8MXpkanoa9QlROeir8zgRY
VaPOtO05/GXVjjAluWKQeM27sa8IpbOXFwbXzSJAYLwrKsQOn5yf9BytE6TuL9E9LGh+GyZ/pbVl
b87D776+Kwbxb8ZffPQuAfFDaQ+83SMh0PRgFB5e5GSNdmJccBGzjRe+UN5nx2NfBBmY9zkmrYo1
3KZrQLePbVA1lfi+tVavs21l6wXK+hnrYFQ5ySx+gW4QJqlalmeggXHQvWM48BdZVEWIj6yTGkDS
Goo+ZV1XP8SeSpmaGVI+rOqna36NvfTi0y8dAkR2YntaO+wfUppn7MRlafcdhO6vY428S1I4udoU
x5ucEmtB6ilZskXn6+LICfpqgSpy8H1H1gAD0aXiQ84t1zF+2+IS2A3IY4sydp1YeNKzdK5eE5Tm
gq4/AUnJS3LZPgiUQvjtzqbMgEs69X94pPH8FLp3W1O8WhJSE5MjuoLyJ/it/c8TJlDWWFIs3tBE
0uaofZ9M9HPgZb9EDIRRZad7ceEjkv/4KltN22fCe5J0H4JIpIUHQ8oJp+Reqcx7ZG/9tgK73VZ8
FiW5mOpME4BHcvaPwvy2CdXvZBEnRQW2J4D5QdzM+H4Dhpq1tyEpOW1el3KoBw3SXeTPshJVFYD2
V2hJZxnSGAyAzb350jsdHbneCu0A6OJJ6fMlslnYtojbhwxfePZQpWA7QbYClylZs/ms6b3B+ank
NwIyE9LFZ0JJGUe07sdG6V+j+sX731mZkObraBVyPXFHTb69f1Tz4xSb1LdrlDY3UcY5bPw/o/yi
xcvk1TWFga8YDqkxaaY9U/KwJC8eP+pfowNTxCn34yEf8T/SjxkAvtjAduoceTStenxjG16HMirP
eWebqEgU9c4u4sGn/qNZX2uOw22TjiRgrBcrvMyn79UXli5G2xGqyscpG9Ygg0BrIDwPGwi24ha6
Nx/FU4XPsmO3fNSbzbORivwblmkrOjQwtFp69VxsVPlZ/D+N3Tuj23befjeCwmCEigu/P2Gdo8wd
KXMmzHlptaEQXkrDSbv9XWw2XiRBvQWt0bcR/Uv2s9bulhS269mkIU+XyYKyxO5U6tdTExfeTjwj
cyBA4oPvpNOZvfsCER4+rz+pO+UNW50bkTcAcaP6O6RUjAjjNRNQIZ8PZoBlNsyNm3LC3O8+JMfZ
/52whsiaq0BIkWkD0rImNbhW9e0HcQqz1fc1CdBDEpTJ903qJhPaVwzW4M/O7YGP9KPtRB6wbCkI
+XVL1eYycssuFGWqp9lXe3+je2ivPw4Mc0yf4JMxjHExtpYAtB13LPi4P6O5uApAvsxPe/ZNCl2n
h7Rz8WIW+PFuRyhmgGKjUyegiRyz2mFEft2koFRJQDxV/1VtB+LyevNW4z83Swyod2x4t9m1aD8+
YLvBBweyF6rEv2nJNkAxeOaNUwPsLD+GbKGw15Hpn1mRWsVtBvOW8b2N3jveTmSbMU0Ub0gy9IQM
cX49cCyvLBECzmQ78amArg0tp0x0dAia9j3mv4wRL1tqz4NG3OKt9T1qvkYXVb/vEfYjVzMkP53f
CpTnJX4TYnQG7oQAiqCPHPrHgbLmAWeRf7zkQeU4yIa0EepunLWWpOvMIWrreGzncK+ghVUDpwrH
6eBYvuvfVAkpd+BgNqM2R2DakL1A5fMhTvc+cgU8f62w8t9iQgE+8ENVv7O5RGGU5cMKZWe+LIEo
iZQmbUq6Zy2/v00Eo3bgN2bUqYChTqW0FOAzNTaBtFPSonqPuBt2/BXJFOBybcRGkSsdLtn7J2tl
+S0YSQLW5fYLD/cC0XEazO9ALRLe4P4ddq8yoqWhgp1/EUur6k2EdeUtaUdBsOr56eJUTKc/lnC9
UPec+GarSOU+IOUfoOB+IBVrAnm8GDmKFZQgCkNfMv15RC6tdxVzzCuZ6HFEenz4Qh6AVt67El2+
1i1JG7Febv1Nd5Z+xmLWAl/OzTyt1SMz78/pOCapGhtqk9QXZdaVeN5hjB3AqcmGdctv2DIKG31V
9lPtS+7kcm/GTk3rxUixM/iNBf0lXDbR+4z/SCYoVtGfHESVHk8TLwxeCNdCOg5xE27mZ2bOnxD6
vZQLNsK2qDPEW8jPYlRHP25ATaorPW/FPYfx8BTWp4ViXDReQKMAIgZsXobfyyAPhH9v6oza/mgj
BpayBfpcMNiPenwGF5AhkXCB4CYPtY85tmw/D/YzOX1bqEZ26tatfWaRGQVWT47xjaWzg1wNnKyw
c5gEkcJ8LvRp1MXLp4JNUSyeDXgEjJAJoN10GT6b2O44mn9YHeHCBEARJlxR/nWoMPoslvN5Rahb
3+jH27W4TC9DQJvG5g9OVwXmBENcG3CqnPOzwbxFzZttYne7Mul+4hYE1t+lAzCtNP/UXS2jbMIF
OAchTfo/AVheDz80NMVnCJ1vE0S48A6KwQ3WQqBBnUKu6hi4Wz/yKtL8Vy/n4peOCkDMVRS5+o1G
UjUG+RFPWcGMvTdiKE00qfgrdB7Bh/ZibFrDIuDJbkTnSE3xPQVv8EX8EvdBxr8ngBjl4855yYyh
KUVhrNY3htgIuVBv8DMYzHGmtUkwm9oNf51KOzapuMFnb09fvxSMJ1oDhFMiVTQBtMkn2JIFwpZD
S3VsMD2PjaNUxUj5uKUPS1m27wpI88d2QvOR2m6YvRZgPR9QhNdL8+JMz57sHkoWc9TuCpto3g0v
m5swUirxUSxLkvV6+UKiysY4FuIY6YJamFh4d0DujvW+wzNcW35ayVIs9+O9NCJbsVgU6nFIpkSM
hdhMdyoJHqzU/MD2fy8iRBHoY8/YaXf/Hd1x+H+U70gnqogbAs1rf/vHY30H/T8DLbaPo5RsUOQg
GqTCc9v74CeB3zXM4cwJE6PK01r9EZQXlsbV6qZeXorSlXUMBl5OFfLYWrFEQRIIUq4Z+hMnUNh8
nSP4C1Mi1KoAcupo4vNlvrantRkcerLomr2pRZ1uch8M59OjKLBiuVYKGRkefAaW7CI3W0hY7510
/h1fjM7WdC6R/7Qbl4EQocUBQRvI81daYz1hiARbP4VlB9rLDT12DQxjjnWVKxfyI5Rb7f+P92U+
WNA+E7OJos2bn7Eki7wClz6EEELSY6lZM77n6Vew7dPAlQE2yZ/wSD/Y93KNeypIMjKyVpIGrjB5
jNDtkj08BObbsKUKKiXoSbD8ypmxNRj5FvxAvfIkN/3Lc6w/o1cKOyvf7RM41hX5e3MDsAA0FG2W
AmSsoyUJvKoOyx8Leb2PvMhvGshojyz70SGXpG/GHxyG0BAeTkvhYv3I80JVF86ylSSzozBCTVTy
wBmh+O9i7gjbsBVuZvoYVGzHdPjbgFg1kK7bXbjgxtJeOpYwuJ3hAY+UVOFZXyqdGf9HIXx0dGgN
ReQtedzKJ/BK4uOXNiScn4p5di9thMbScNGpMM6L7dGa94jgFeKTo3WUpz0cHN8n/7KBomu0IvvM
/Nt18PLFKM6csUkkxd/aGcj080J8d6GAnIod2Pkox53rsBxjZ0s/8LVdPjTNCdjpOAoh94uhTZRi
oKHyEypcVt6QaKtaq+e7Emnrc6BgZTzxnPW0xEUMuyKVY+vI272K/dpowPfsOqIUbX4T8TtxaGgt
wv5L8U0RGAALwpv+ucnT5TwYi3J9qKCS1r9RyWutcM37swH30RFmGA0WgaPbLk1+Q0P5CEkpa9AZ
SG3a2K2Tre5AxJpeyvJ5dCnYomtJ4ORnaQGlY1KS4xzkrbtSHEDmuag34sz/vgLV2ME/VtmGqfjU
4F8sw7YnCOeRQ1jyXQh+XXkFrLzbOAv6rCZBBgZxCjArDV/rNGuv6DQo38frmRK5l6wU5g0Obeus
OeCkgPhS/AG5S7jTjnacYGwnGF+0SPEYxvrmKHV5TcABRGoH8wCduZGWgGzSmh3xS7l7Ugq1nERW
9zf55kUEBxyqsCliJ1fYwaj20CnrLd/liFl3XkHMkc35WzOIxibGSrIbtyNpBvP1ZIkBm+DX3ufG
HsRqqq3z4W6VqCPh2Nxk3N6Tqi81M3QEErqJMaZNNtijN750eIvOXGDkcbrCEDmuXOoYTBcUYZSd
IbZICGl+Z8kxbPGrBHzZhN3ww5zCT1rTFS2lNQQWioW2ir/3l7F1Wo0tp/7OBMQXtxOeAyX0EGEa
MlrpwzKWGwbJ/HT9SRiXzzMU5VOz1dgBDqZ9NHNLBefpzGi+x43Ft0jhZXtKSEX/mCRl3k1VQQCV
HRmvPDkRFFkBkrpJsDd8zZP767UWzWwgOqSNaEQCnC1q+X6BPuJJF70OULja6BwOyCRpnB9VNnWK
uqN9oD5WqBGF1oLuOMPllA2p6G/J/tPwDPSE2dEX1VqqNc9SYesdl5Xit5+tStgfuYK/0VeslkN/
L4D9etv3fm5FWo2EbC7N0vzrsOEBzxkW90OsCzHBSqi6Vwr1U0rVZXxY8wSUuNpM26ucvdBaJ+2K
R3kHU8143jdnG4hogr2+oLXZPfcXD8ezltKwPW6fBGRHk/Y0+ObEO1JgI7CHHl04Wh7IUcbycOym
vf8aC/Lg08ukk6fDHl+OkFtJql23oA+xucXeDugeYI2+pFO5lPDFV4hCYrY+NKSwD9QKwctoey41
W6Vm/jNgZd+rh44sRYbAVJyIDmbZrTz9fviFfy6mmi515UJ2aVQvG/6V2/2UB2VtISnNHcVTHBMQ
OD8fRSPScOcLfRmyf3jEvfCurRchJMGFLf/TNDvEqzSU7yvwHhU2l8E9W1E/r3N/cw7rgS7GzX3C
XSr2i8rRDJBp7UIlJUJfpFXjfqm2euMMlyeITMqJUfSZmF+69L7PtIifukNct1La9h6YIecxeG7G
yGPtmnoynLb0B/t16s0DACjKu4OpW8J16EFXbHWLatZ4j8OlzU5susfhqI2AK5BezHKA1qdH/PkK
FaBEqKIaFxkNoZZx32NhTaw0fTKLw3rXZDOuM0qluhOuHwpueuwRO22chWDVk8GiqY1hvnoNQNkB
+euBE96Ldn/2RdSz5QMQzbA/IPCfOIohETp3dWutx43Me62gza2XV+a4aHhThLYpofZK3KWO+XUy
5TAvVedmTFGVLLqlz/OqiAmi/DZLWerTyupbVGfK1TwQrp5hmm6KoQQmnv6aSrwwlAuLjImEbowO
720itbv0MQNFf/WoScn64/pN9EX4EVqpO9ZlhH4CmewJwaOcJ9NItd3nJbh/VVQnNBniBV5ucoqY
MiezBUCocXWT5+Cofvl24HGnsN94U4/AsHoa+RyheVvB+MisYwUCCucjU4SSjtFwEhUubgum5BHo
zqnJouyuUKzmc13VZWWZ3PDZpdSKQTmS6sro95SJcfZ/jnQ+43nHW+/R5gRjIMXCbTERUNWJv52Z
/QUMLRPcPASRpomwjBD9zRvMhQeFLlmQAiz9PSfHMuJobuUbe9KVxwvwednMMBGcJ9CCJDcvotrh
e0dQlE+Ln955LTYaOnJfZqGy2vI+4vhWevFYksXWz56AE2pmtNlg0g4K7a+StGqSNtxIi9oF/KnN
4nd28K/TsRdjw1Ji1qnbgL2u544y8210xMiD6JQDTgr5kXs7tTZGUgB5PZetsYMp7caoDXz1zycP
X3c08tgxHOHXbLGSvyj2HCZqFWpwqibLZwcVlfOszI7lTFes76UTgKD8WDoSxkBcfltlpzpkpkxY
zGw5Ica2OcCoIZPkxyT72BqBin7KDtQ2LnrU4bIvDLv9FnJBLM5RkNEvek9ucCj6bJoKdqHrBpCo
+KMhByd55VzToNLuA/nJSeDu4rCvipxC43XC7VCrzwgPAeJCmjWXJ3h9WFX4mDUGS+03Q9mtfBMs
shD51zh1LP9QfeFOOcW3t5zuthtYiKhJ2Kju8HU9tkeLdqNoARRI6vwKCXtypqpectSjRjnbC3Rb
/pQQswX/bAuGHwwWktuaOgbvsEipJEROah2u/tH029MlUaiY6SH8v5XNijNAI+buXiK3VDDhy8Dp
MJSWhbNpknNxdbhXLdohSfK+Z2mjXW4LsV7O3Txtdm5B/POCe+jsK3JgdXcxa+eCBOaB94k14MkO
Sk6s24029xkENcbTuxD5Tm3S7Q1MSjW82uOyT10SdPFT3U7q+uT8NWPHBbz8+OOQIr3/YKtdX8F4
lkOOdNHAo1fq0WmBbL944KG1jxNY+eSIIg3OGey6qSZCf6Rry6NqibQq11iG/ONuUIJEWeSbHgUg
70ObiwrPnZmKbdgQO0zkTZ0bMxRjAYatXVgxDvuCDvBpxZB/Jobctp4d/OSKPzp6cyYi/LvqtWof
p416bAGYRv/1U1FCLYQNrZNGAxOhxBs0Yds9HrchHxN3vGGIideJBQ5e7BQvgMceL9RakDCjagr/
4EijqIQqibjwxvz49pjClIrHnnJ3Ose/LMk+vM9ncQ/icGJ9Pl63WPsCBPb51lGeHBZ593pw+//8
Jd3DAZvhF1a4v4y73+LQBnR/IRWbhSfJsWSqr4Une88rLqj3LyoNUUa6jrkXdEbCjm30EL5/mawc
N6LZUkC7TEnmIrlW2YiKC/OwiNVETXTl1Zr4zwS5wk+iBCESEK/nQQ8iWfpCY6QFYJIwZ9rKgxiu
gYhRx/OVqgP1DMiGvlFFmrJZgNF7UGkk6hw3zucdu3g1qSpRboFFjdmuZounctkKgI2xwooO0F/T
Qg8lztXbOQAUYsyecJ2KuQ+x12OAU7vPFkUCZhGyZ3lyx5pMc2M6niO7gi2wru7V+8Ve4hCOsczU
zqhQWtp0v9Rfg0rVFZtLPVYUOvt2m9/XdwTZo/omeuUHrw5KLtMyHuo8iKl8E87PYMzNVB/x9QTc
gUk2njsmaySiZdmJwZ0Hei2B6WAXCpSo6Ek93PPZLSTZF7lApC3J0KQl8uZxIX1J/m0a62jpnusk
Q3Dka0LpfkmW95yY/L8oS8vKL8L1RhV/x6BUt+mvKQDGmHs/IAmGIMAeIU7opnMuPmFqIoDimM7J
asc7Uxmq50sHzjhiP8m1FB3K8HkFvCGCMIKSghBPiVwA0eUzPNIUUSavt/3ktNT2X+vehiUb+Nx1
l8ofXf/YPOYD/FctOrEQY6BfqpsqAfUK7rVbOcAE8BAU0Q5gC/Ia6cA7ymY/D6Hha+/lw8wH9G0V
IjJT9GHjaAsVSchoBgNwiBwWvGPgzM8Fw2SECrMSfgk1vFNuen6FpAd5iPCvrbvmK1tkcyk+6Sn2
w0ZnZh5PRnlh+O0dSc941kbf4fxZ+nH24dh9d6bcG7kl0QWZVk9G0emd9+cW4lmJ6Tlh9ZE42yd5
SkVfTFHEvACycrQZDyA3bc0h0RNynavh4AwvKkEiBSWo3CQ7Q3yZlhwpSE+w85x1sTObpCHKUdgg
uoUYPel6vhX8fsypdbA6MInHfR3n181VPVnG4/BjWcGq2lL3VIMuin0rNHDABo/EgPB2kry4LnNH
fkX5+sDBQ/2TIPySTM0pGXQEgfDu09SHmNK8YrKDP/0RcF37PlLl3gXU4tP9qCZfo1FGMnDfugA+
rgUCP7tPWLGfRFFLy4yIDRBSO1fQjfT2LccU6MO0W+KNICpgmbm4Y/Rl0T40BqmsWya9bBiTo+qS
FcWSlG4rjBGip1VcGfb3CDH5s1LX5m1refUTYPFal3JrBWEhl2RYDPLUqayxQdmO7mQLqBhdNwdN
ooJpxHS4sKD2FY2IKFCLcgfuFBitxNua1jIk0gBmh9KVQZkgCY+4FeGsrGvlZEdV2bjhzkgq1Jec
mwCbp6s7YoCf/t6lDQspSs3kTUosQEC5/mT3+AAeElFv0urWGDUD/lZLSxJMwWgyJN1jp8JOdAOz
YkUEVRQKV11c+SVClzfBFuueKXry07O4ZuIAxkDZ+awqeaWjXcUfhsRHOMAFrh6IzwuRCFaPUdhw
xm0YPjNQX/suCY70qivbJeeFC+iEbsQc/jYc3AxOlHvKObyJN3nckcWJtcs+tbO4yv8ryaBfcekj
kB43cweuqCd2rOzQ3ZInED5dJJXSk4d6nlFC54gZUWVLBSkdhr4TIMB99oF2X3/C4+a73Ktlny5z
Jj3mn76dQPfT1g+EHDhKlOPxHqN7Z2i0b3WBLe4/PVqy4qbyChCKtq1prP0/5CCsibW2xwvIH3yt
zl4IlRue+aAwVMT45cQNJYVUcyBy5m4osSn3rXc4Y7Hk6VjwdpaYq76zkCftfRIlRNy+4jylOvuR
jsNEVwHGNzYxl0Ly6HUN7edECl//okwPrumH6cd+qFqKc7TM1pmYlC1M0uwgLs5IfnBXsaTZHzw/
CGK7OCziGhFu1o5D5YOvNPj0hJht4XpKHERyd7NgeAljD7Vx59WDuApI6bMehsF2b98DoePNJ/lH
WAN42fTTzZNGHa0pgTbs6+Gtb+/KHZ053JYX/EJFBE/Iac2wqwnXd5LsWxiLkv3nJVjCFnhygEpM
5YhAbAWcQ9cQ7Kv5kwkkh2X0E3cAKrE4Xg1SqudjDr3dQALgkJqJXQl0LLQ4MbkZBOHn4jNUYLnR
CoNmKJsWvWrEFMpaSlrwwVvmfC2NpQHsEm1MrhyS9e/TgFKEyJCjzSvwdLFoPYYX61cgpuk8hNEl
Wv1tAdTTGslxrHzPZn7cMbPN/Z8PWu7I8G23DlZUcWG+scjyKmheNeEua+q28HEm6I1FUiQrGzVJ
/hbgoO9eijmfnjnN/2+gOPDWrJ1j5EP+AX51osjum83rPBbmW1/FPBcuF73V8uNbDYCQGtBCOBVh
HoZZJyAnXpCoVNTc051YF2b22oWqPVRRkqC8yqBuwTl4BnO69J3CYyajvb05O80wVl8uk2K7+l3R
zsPy4BzUfDd64+yTLjigEfZTVETEE5FoC95NoMPP6rVjqNN1NqriGv7HaJg4Gd5uB3kmhDLdZ6ZM
J/+sIwF/l4q1mbk57xrQcsh8vZWg1UC/fPK0I1LZqOFNKhZYrrF7KpowWy3F252xanruZ635e+6X
iBtfAUTB7Ke8Lr3aAWXFmyUyIab0OrnqiZ0xjUxQoOQY9DNX6XqvuoO9I9j3FSSyofoPbfLQqmoU
8TcE/h+Ox2k1oBtk0620Pu3TvyH09EvWLKA83UKYw+PewocKcIUj9R/wj/xLk3RKdzD7TvaiEYlB
aZELGbJ5oos2ZR1YH0MD/LX5LSIu+ejEebpjfkxnhTDe8QmDAmIs4iHkvpe5mDWZsSXEEUu0wR/E
UizU+z4hTDwBeZE8hNzu+cfqZctT2FRufdagkfoKD3eXilBzk3WQ1ecZ9w8HK1F5ybOSO5sv7hUn
MKcDg4NysaTKigjH4xvxddiGfJ9Ei5yJnhIJf8pTdQKsqj1yAnWOVQeE6ojix7d+fEMFyvGFabzx
/2oRG2d/eDdSKtmhQywvjP7HD+0Zoy/5+6zMfRYtNaHyQYYASQ6HY/qv1uAbNKIJ4T8b05Ku/Oq4
/3TT3911Q/EQvkfPbQSjqoPEh3yCxlap4ZpRcNauzi24lneNBKx1VK3XOSpwgOzP8Lo/1ZRpHUT0
zG1fLdqlGsjGq1YlqqSQF99BNup8WXPy9iqJXkILQmN8FCLKK1AqUPk8mRcpc6jpS3vFMyWrJjSI
REYhK6ZNjWsJJEWlFj4yyd/LLz6EEvcxhMns1FQTj3B/h1RLVhCIxOIJh5TeG5WYTF72k8MRSgCT
ft/1lZPxyUlUIKK6zaxfnoxUVHwIyKll6Z4Q4njqL9hWhVP/Ve3sKlGBSiqOQPy9qt+32bnQdo9Z
J5aAT1g4Xp3nUAUFU+E1lAKcnmTyTyY5+hc00ce4nqsHQGRuQraMHwXc1UOn7WcunWupJ467LAT/
9MrHkIDeYFiJQd6jEcqfSEzskbQxRzHqvchoyGlK8nteSiEMZRyuOybq07s9pA6b4X1XO+vdJyEB
VK9drUl8lnqeyXQzhtXZNypg1GqjFnjDHVidE8qmEkHCilVYYL7CqW9vEKIDbMEJPOQiQP+4maVb
OYiaJeRQ5ki78LQGffGn2qgoL9V78xOwnZQDky96lCjAd8Ba7U9RpPAI7rGjgvL3aVR48mQeEAih
P02sFbGyKi9XbADZFOAV20D33kYbClnpskSUmB1ZOJCpspUUVSAOGKkMk1afGuEyFahokK0Y8iWY
Wuv6/I+GpL+FFoA3YGOLpzNQ2uvvdUCA3IcC5yFutamfS9hcElBX8tXECf0bPYJlzjj0xpyoUpMo
TnuDrr4ju06qh++MK3beaKixBSiKc/n0jmDHuIur54BF2m434GYpzjFrEP6d8iuh2mfb5eDQeDEm
hkTcsZeBlwEHB7dtQW1eTRs8vdzEhuHRRD6yksZwW5YfaQOQOHdDSkE8zB2tXQjhekE9C2UuyjCy
soaf6mxDwAF4vJH+7Emq2G5KtZytuQUyIiPOCbD4VsJW+LkcjplZW1ufyTNDr+25Nu24z2Q3LB0i
fhQAzV8E2Pmlubmvh9AHgcONk1pZpDChqjmySd3RVlCP0fEa9CSQtSwkmSRjb4O10aMoh4b0vnKV
b0yLIkhpHG0DxTBUYUEU5AtEOyMRc7dZnrYUOYZvIjYw/y4ekcjRxvJEEAc5zkEDoViLoHWkdi/i
xnbqJ8HcNXmzEXl1GdvMsGHZucQ58nYxgRTzWquR0qnxIh26mfLkieYHpwJd1gAn+LKoagtoPfUq
eIKDvhudqPe2izfe3pZP35h1v84F5XTi5mVrxCVZVW8m1fO2sSiZGFp2sMhRSmqZ2b6wcGy3V+Ch
B7lWljBIRzbQfzkzzriX+gEpLXKGNVMyx30ww+yslpoKRWp9W0rtL4tP4PkiheAhb6nUrGP8ieiK
/xYvdT6kbRhsIXtXjpE7qnyWcoDCy0QDmrKPT6O/q2LQ0INQ5APwbzAL0rUVFdZkmzoWBkCHSKIa
OOnxWvMDZLuD9S/hLxjJBS8DT2vGs8HOugnxnCE4QwpxEu6q7cZH0gIn0TCpkRQQTvWaNv4Mj1Dj
OAJ/ppsYNQfepDRr4yKccdD/jAz5Iaf6iJvGssE80sNks8tzwH6/pd4omGXhgW8VbMVEovjryHZN
yWPJAjtrSbeV24cBQAlZomvECfVbWsoHKyEyulVspm3pO4XkG+lqQdA9TpbmGL7C0tvXvi2fmF58
uew+r4+IinPfB9UWFWv4/uxQ6fkxWOco4eqWAq9+hPxGtASH4YK85r4HmCyiwHTudHCH8toqfWTQ
pMhG5XAGCHRTa17FpX41sUlFVt/VXIk/flGM81HUaB9Ctw7GJzXCxoZ+hwMa4mKgOKeHQY//HJM8
ulSNBKXyLse4lUGkOHLj2vLG6Qn4ZzNuZHyf52TpUoDkvRd09Ur8EDO43uqUueu8szyoeo/ukq+9
2XsgzTszTImnbNONtkkOA5xblLrHKyG3PnlH7aAyB1Llu4oI7mlj0LsmXD8F4HYYwKOY0VqJiVcZ
eaqU0fU01QYO+0ss6dFs1WeamJRihMOdO20r/BaKA/2xm0FlWUq+qggwcIIs73HZTOpaLEbyllK7
Rxkd0Z7Fvy9fI6AC8ZaSPh6YCj1Z78xbSAsCY8IgD52i7XndgAfr6Nd/yQlSDdlkSuysVpnmYn6b
jmTZ2bKBcd/wfzVCLkudX+5WaymeS4obd38JcVgjEAUbVLcB1PTXGPNqIEvJ9Xkh8ITpUmeN5Ndk
IhtZcUJxEgEpREbp9BW0wz/yFNHdaDeAzRTpHyPcnIdvjYl25ufeKgvWDaKcxmpI92A12CvvWVBE
0AQJB5oJcew9fNdJ5FwYLgnb42cAK1FMFHoVDjYgcYmZ41Ct2whCpsak8lKhM188q7gecdf/W+Er
RqIxfj2h8fQfB80wfv/rCF3J4mLVuvirBOfdjm1XcrHhL4a2MKdBikgiwfkx11cxw2BUd0VAySRq
IHae+lnOw0Qlkc027vonBbDA2G5/CjRT+Oy+HmCR6ShneqHrr93QGRUy4xdNjnumfrY0N8vc8NJ6
3wXWNk44lIf8svR56h1gda7I7YyXGwVh8tj9lxrAaM20NPDI+Jg99WdG6zT/vL5tCg/RSv4LQ8Of
cj+0j/qybMEkTO4/zng/K4aiJENH/oh92gX6lDg0AeXfQleoriQq77V6MVLyvDVmq5RMVg07QMKs
BKvRcG1+GeRp8l6rVnkibuhfBEzO/wR306RQC2sS+mp6laA1wCbg2ANykcwEYL8tEAmHXDzey4An
ZoB7lbjPcRoiXM4DYcZR5Z0g9NZ0b02aofOepAoFRtX9xrn+YL3CPryQiYWVjKCDdNJk0lwIrWVx
0GMwI9ujk+hx9twNvRezdbr0memG0ErWDH32c8ZjzN8C6a4Ua6ItikmE0N0MBu+OAUd6lt2KXKDP
qc2Nu2o3U/RdSC+PRWsdaQHepVDo0bDNJFPZwbjGGj87/iK247/BSFCIB2hOH/gTkbccNAkB2//4
if8R+5Iw/6KEtAQRIA8/eB9+Sbbjml3sS8U1j9HeQGEflPo5onWkInCVcU5xaW6bVOLpgOL4CcGU
qq5SL6HKNO+ReVWmE65bspuXJA9y6wFVQ7YTC0XM0bGxIhWPb2h6ZaG5Ad7U9+v06fo0Tujrl8EI
p/etD9FOnkzBpRXODBas1vmOi5DA3h2HUTGwkgfx1erxq1/lA5OCkTsW7piwJTygZMc5tE7xlzFs
Tehs0cH67U18/F7LQ6F8VHMeTQIkOpMrTiGfktRcOKPiEbh0PCJN3aGaWLzJ07BLC0qn4Xy5uTAv
ntu54McK7mOgN4yGi/rcZV1cEyBc8GeI+YC7lKd2FXYz4ZJWwxwuwOTWcY9kFJcNlwpq41/DXd7d
TSnkJXHW3gzkoPZWf9KIQvfSqfEL7RyMe8I5uMcIJJt4vohX0FVLbePylOCDmse6E+RDZm/0ruES
k3rSlL4sc13A1juqHcOiDf9QuoBqDXfpX/F7jBtyCUsKA4AxkCYqA6wFvX6fKsPdfuyPgCqFvQfe
2jRGvzpRqXCcrtq8zaXwpb8rEw0W4So20hCww7PckZ6pYPZZjjvpA7Q9miEp/ndNQUrlDpFBVIdR
Wem+MNwEzVPDTLvVTdu2hlWS+dD609BbBCgNyty6gkCdKrLhLSa25/vodkAhfMxE3xLdtJOT+ygC
YHIq6P50rsqbk12S7u/dVGbMXuN0u3/UWgJRYojHbj/rHCEQXeY/vN26ZULSwNRA1BuoEiVbd4lr
LURytDIImCqEvKHF2ueg4iVgf5eD/eNriwDisTpg3sLSG2Az3om69KG4QkiAukHQ4d/V6riIwPBK
k6HEWeZONFKuBRcydTRG6WcGaBXYQs1vgqg4S5w3ftj/VVoGEyp8GLmkoIvGf8pSCWKyYSsmmXeN
OAwHcy/UM1atys6ATBpwVyW0dqLAz4QtL6ac+0/YkA3O/yx3WF2C2AdvKaiCKSjjbmkxjoAkA6bh
dyEEWq1mGkY5ZrwUDizabbENoVZyx6lwOTf9g45uwxzfVpMIbYdToqcTyIwhvJ6Wj93XVJCz1VC4
gH6NbcHNeYpTba059PvgDTBjBBT3mDWt/U+tbgrsWrbgUZ98lTTETVB6PXHHwgBKbnTfeGTMIwzS
FN7D2bdYF2lr81qoePpcrtFQNPsuwuvtFMON+XWzmwQ+qZspgZ9aAKcPzrHctZjJcoBXCdT+deIa
vHKnA9yEw7J6scAjgC43c7okBWrQVHYGNempcvW2KmGqq7tDSn+lNmy5ju1oPGHFlSZlXziCgw7F
mcLfWhhJOArjr0Wi4TS+aShBdJE4Uuu2uVNnKSylMc+1/YnzHYU2Wd3v3kyCb7v/fnI8/e/ASTXv
UkbN5NR2AvyJpeKTxAm7lMXlNMJ9slC7ArUTVgpH48xLQYsRNNCHtBVCaQdEKorlj64J9OlxYp9y
Mv2RGPVlWYDHQkeqQCZa8PZyyLKKxjRzC3kCpkcCvZ7t1KVuwRKw48CZ/pz+iDldsXksLvNF0xxg
FBssD4BtlS8ARRg7TkHa5eIuV6y1pTDUIpHn3wFd7vbSJ4gioBTkHAFR+oV/OrzYsDQ50W27TYIR
XgT5T014mwIKZVLi3h26N5VxWxBtDl6F4pADM4CdMiLXHklSzc/+jPTWxWyZrAf90eXTh21WeBNr
DYaR9dChF3vNlErOlMSJK/ivN1lTEWm3kmNyuPXSC21OAF3Bk7ZdfSHGE8QleopGECtifUNi7SgX
8K2JNVN9J9U/vssYPy2l5MJXNchwUVi2UOBg4/YD7JL0eNeU24SA9MS4cBxm8ySYtbtp7TdyNicC
JrOgNuWB1VzUkS0jRmn85A7jvw3Vzr/bAMxeIpsWU7c20tCbAn0UJ/ypaqN/RP7CnGMZp9/tj8/p
YIQ4qS5GGUYiWYmI40R95mH8CBD6jyAa8+4fRz6Wpa4PBRB03bP2n1PgvY49DDTscKzj21fksOJC
aqPunHLsSSspyX0maok4YNdM0QpuccYXLwHTZlWXgNEReU+e8sb/UwHB76oLJZ0po6xs4xRTFlkD
NmEUOngVFhgnqnPP/tQPLEzNgYmPRhNY7UTWn9FOcVbQbAJ9xERyFL2xBU1PlAEnjnv8qs8K/dpg
FKfrT+LAse91YECX4zsoMu9Wv3Jf82kn17OAJDjiSSgOTEm7jdqHWQBKyyrgod3/C2+AFOEvR/Bg
Xm0YGYEdZUmp91eFJgajP0xgy0mOzqYJZwbqgbHyucCIbQ/s7gtQqEqRFNqZCpjrVgt5lfwNb/bw
Tl8h0pgi1H1gh77mMFJKtZP1pY1lK5m1PRXp4TSzL6BQM0G8EuRUbHqROSMYxBEuPbWIrBluBVGp
Nim1OxILYoD/YcFumKmn3HVfQ3cnENzKfp/zUJSekWPtKwhiW4ncQvvOl9JjSjEzia1Hgb6V/Tiy
uHdM6Qdnz3S5tlP7jUTpLF08DeushzF3Kk1Gh5dmFRJOlm9Y/ri1jdV7ACZvUYWLTq9x0R7ErqVk
0fqoAoGtQ0MvNLbCjw97vBR9OFIvIb2ufEN9lVCn5CFwP31p0GNPR5hNhcltT8GaNtq6fOEpZhmL
QkBr40VYkNaaH6ZeWfJ2K6lXrORmDr0v1Bz57AdFotMsQOXxtrvH1xyJQLjB0zCQFgdAvicqFDUB
2hFgVR4SF/MOR4U51wV7tnLqE+A9RwaF3Ryp9SbRDs19GHWb3ZQMnYHEpXFAzP1O2N31U1ODT0cC
2miLYfXad5PF+ThLZFBlYzcPnzxBUhlJMJDKEwAVVXr4OIBA3iy2pVsk5crmuYCwH2dUA72vN58N
BWYFFgT7W2jS7gOfhS8oc2G83/nUcG2Fi4V9/kMpCqcJ0HiJyNBMix6ozY4U4Zr7qullyCEP5dcx
Rd29pZW6tQxsVy39XaFIUdq1Ht+m9zKi1PlahXuhu9WmAME1XBoSwYSoKB6GN/HVOKjJkzFXHgTi
aAxhwaVmWgLTa2eeYFcJdAQbWjhqDtYeC4fw6xkpLRL6x7vQR3zzAeCP9gK41MuZjwAm5SdQxAk7
HhjCAOWa8rRj0P2cOhIiy/97EkcbmNpe2j98p1nlu1uz/Li7mrDztr3RO1x1zC8/kDXBhVBPKpMj
4MrAVN3H71OJcblLMN9Gnk4BWZ7ualVxl0Gf47aUW+AY43cHsjw8gSQmdi3KKdGf9vzMKdJy4PmJ
E734edqHhXS9rvxwmAhhjT1mhqJA0jmzDFI3dzPEWF6HH3AOAofbk7QylwX78HAKj1fL2S0URFHO
jw7K8XF3MJM+qzEuo2QaNB1Rw5PMNW+VE5CjtHkACENv45vYYteqh7fRaSSz7DmpsrXWcg7Lbgj5
JyXlfqKKPWSFNp0NtL8idtA2VZ+Fv2cmVi4A71NX3qNcPyBNyuM0RIubRKGHZcoC7nKdV+Azm6mp
OSbphrkXTXAt0YpIpWxrC3kV0c7lje+Ce549546dWOXFuFaShiyXuiTwhNO9JNgaIDxcj/buUsQb
CpAYrK8NMoeKW0ScbvBa2MKkxOtkxGzWm8zVryRVo8Y99ltSziq7u8O8bb21xfNch3MxBYSuuStC
QRbu6RtiZk7w9LM778ZBC7nrnpnaMbcOn1pDyIoxDPMF+zFJRYFHdmCux5ILOjEZnREChJ0zpgKK
/hTgRSuPlaVWPE1lplofge19lqVFmWM8IJqYb0HSErAJaItW21I/pGfv6QG6n0+GRYUYAE9/PTv3
8SpdEyYqFVQ6vzMxGT+p6RdyrPFYPtWUz44pWXx810Nc1Ls7YK5XitgOxi4To+5MsBxl26L0p1bz
avP0WleKzNGJgR1lTSuDnDDwIxvbhewEO33gZUZs1+AX5Ghb+ED43j8uCxwiijgIbIR5nL9TzHYo
5LwMvgos/TLHdKiuXcdCVxIhDGh8JtfmftzhsrQhdX1tJz6RzrBJOSmaFhP4Yg9KCIUkAvSglvH6
af7wsWBdqF0KC2U1mUyqcJD39/CIs/K+PNlykxqF/rAp9dKuvlpq/78k9ZPHVcANn6c6MPt/ZFZg
ZjA1x9xo90l0Q8Jz7nIEypXt5Y3DaLMvDERfopNAhSbH54PBSU4QzlLjGB4VCfVHY/shMq4tQ2it
Nic8DwpA/z45c9MsTYx3aG79D6UWvcMNc0ArBqAEn0OAjvwRb6rJhikmb2tg2rb1DQYbs35yV5QM
y1KndsQL01IaZtE4bnQLcO4OIcOIRsbxT9pPwmhFgjjCrpvHDm10SLVtPF+U4nRL9lI3NKNuYXNB
0HuBHrOioHkVKbtSee5T4L7a3n1UIWctVX80K1S3aoVZybQR5b3Wnli8y2nrA1f2PgtqJkzZZcZ9
i3lccbdeMUmrYBkgBYog7U5l5kwDYaxezVe/M0cgy4N7GT2FtTAJW0pSAkmxJsIXUlebzAJnPoLX
Z+KI1Zi/C7fd62u+QDMX8i4eI+KL0i0kNkOEbM0S/8VD7WMORV1YTssIZCvLNiIi5JGzhHbYan9c
VUNOCjT9qaJA6Xe51H6+z9ASy3zP9FwAhxuXM+JAqFSmEISIdMNbviyMUNv5OzAeEIsqZsFr1SG3
McqNohcd/tUHXTBJVW692gdCLmK4G8a/Atm4lTboSz2gSHQXIQtOxRu0NM8764IgE1lCu6zuWFx/
90cmgvfl4bj+r7xtVbgzLlEkEPq7t0M396DNKnZb3DfFtjuBhD7Vbow+cxri+XcZVo6N9cKm5bWw
zVZZmj2/bB7rU8rbYWou9jQ32+lSsYqPSA83EAKDtZDTL0wUfCM5wS8raQaH9O9De9fotmkZbNuv
mMDDW6Rdlso9vwggefVvkbShUSuJ492+dG0ifr8jdG37crEHntjP2oWYr6X8NSvx6C9H7v2mNW+r
DtYK1Iuadux1HJPVcUg9V7Ote+y3lO9uVdLhfulcd2kkyWGQr4EG8hN37DzoNLtCBhXmH3G21FGd
3rf8rTBSkaT5V8iOoYPUAkU5w8Hbo4nPEQoUlApbRU8xqC/apWYP3ZWpwd9zzuLPYeCKtEOt5wJz
9/9GHZ3saE2i0NToPI0Hu582WLKrT1bzrcWKd44ZoMYdG790WQH9p2JsZyp5nc9+duvNQa8DO/Cl
f4+NLwD4OUDSH3K9/KWcIWhDc+vIrw6rVhm47bsKpUcGwG1NdrAwAh8H7rKDF5hPN5IgTbgKV+eq
SshhCtZORMiBF2QFs7loWHVF+hfATv8KRpQ0nE2Evy3IGoIiEx9EdDwwZta33NPltZqF/hJLQ96y
FWrfe3XWBkVRvWEQrXyosIQjO/EamFSAWAIdYa07kBfbgSmjQk+r3CXJm3INPtLqTEjbRAuII6U5
n/bQj8wFxUaxIjlY3aJDGf3lnaJHBhXW1HezL12SL7g026o6H1bz2c33dVB1D8CceMPWfH5NIZwg
BXvGm2TJE12qUVE6Opw/aEI8SCuySl2ZH+HVcfIUAGTxONhZzdK1S8xkuMU6V5+0sltTEwaDSxvn
qUvrQnkPYMNgsqjrkMOK8h1XrAOFbT3KtxcdGkxQiin4yAvmJ0N9xGVdOtZHwMCsJi7W59RYEPxK
POVAv2NKodbmMtpmtmJOxkuIUFkdG3J6wbX7PMGUfYW/pCQ45C3ao6GOSdhkd+r2VO+lB60FAuNr
IZvb0gbESrWmB0bNVLWHtuldIewlBAO+ePp1MHLL/QdvdCQWIdJPqfk1rj6u8l7vq9r5I5NAXIIV
zEo2FEqsh/lcFJBAqXF5bq1Iik3BOejpLwp4TqWtcA3va+ZC9ytZnMVECCgicm4tK+GmXH74sa5O
rcU8iRbnvLC+JBCyiq+7s2SddAB9nvaQIcJ4M66DBzcPf2EbCQGOLLFVf2HROcGqj5UUPZdAm1ek
z+wSh1xyLcoFq4HpOtpNc2A4Ziolc87dP3ypV2GrStbE5TZnO04YmXHEDwbXzH2oz16fGCYJ7Y6C
xDcOiQtUHoFNRfq4sOlDag3g9ZwVqwhk3YTUu+Oi1zAbIdD/XeFzhiFRAi9MjVzSpevVDJUSKiRw
L2xZeMLacQUDVBWgwZ48ynFh5GzP4tuJn44+uzu8iGRvX4hSqqelzfQh2udf9d9opVycUIwTOFeb
TpHi1CbhP7x5Z7oc7PQawbmsqVNLWrRdUX63kNvpoqja+k/3LEdX43OiBTAoTaqX4UZOgfThT3sI
1w1o4w43t+QT9NHylMZC2NxuGkhpRdKA9eBLUCa7KG6063+QAqrN8zQlZOLRlj8ed54C0pXvb/bT
KRgOnWP5thUX6RZvFIAtH4ovrGck+PZq9A3WAzJYprzPnYIj9beE5IFfVg5hIbK5V8tKwh8yRnwF
ICQUh4WphmV5G1I5tH8PekYn52MS16T7792zq2IGV2YW8fuwaCR2Fg7AXFLht7vMvBZLm2NUPq4t
wApKyJCJnhifVHTFqi49XS7XU4kA2c8dfbpXt95Vt/9xuQv6okP40i3PofBojFsemefXVNuAjJFU
gmEPu7gkxVSnEM383fzM0ZLYZ5kc/vFkUyYCSRnaYZzcPOdreeZZnzbhvmJevPOA4vhwCVNaGT/3
3vzQoNrNk6a3QAG/ucC8ylKB24QngEtBb439KxtfDcOGpz/OMljrJW1UDvR5k4dr71IgY//ogRRg
Xf/xA1u8fwd5OEBIO6m+lLUf9H0JoyS5cEIqC+qKpT05HKsoIovmOg6jLlqtn/GkuPo+IuwXS4Qo
+uLf9usKKu+MjFeKvEOh00uumq0ZSHtOouwCYe/hrHzUYl9HBhocfQn2bppPNKRMeYvIGC8t+Ezp
q1WpuCB2etundbSTLxR27uAZezU65RHYY3NX+qPcKVKeOM2gORisGRIRlnND/MkJDLLh4PGH4ctt
wcupfp8fECcLbr9pRpLX3amUg9bsGmVI9HgZDK3FCzI/42vcOEPhSdiB37fx/p4d6yCM5O1mIHV4
uJNDdk3Pknb2cTaIzi+cK3vVMyVddImNfo3U2Q1zADJ3MPt/AGaZWYA5LttsAcg0kD3Qh9o59qMl
ibtqnh/De4qbWpOAKHYXf/jqCnvG9KjIzjZJLfnBaOvFWNHzINNvYKPja/EfbUI7uHpSY+0wirmo
djgEJch9JH+K8oIEmFZ//kcXb77IC4XyKnQ0vseTifrgsvp63y8v5qtNfSXSg2ebuzLl2HEgWaBa
OOeJCQjEwTZdn13ulNldDZKqIzc8V3H74mJKG9S/h6OhHCjkltyGbTCjUooph5gNe4FtWTd5dovY
QtaDwBw3RmfSViqDuXdQ8fhqluykKkReTOLIGaREC5AFaOje5GWRKU1ZOzxIKngiME4Wz/uKRY+A
GT8ki9eWDNXX2lq3s/urQocUfDUVinhwDbp5o9slOTwZH51eSDowu9SXqClPoyj1UMZsqfk/EgOO
E2BHG9UbaERlimwcbfCwK1oluHdX1ZHUc52+q4sgXqpnmzrQ3NnWJKD3tKOqnKWpNSsIjYgxY2J5
KecAjun/n+RSGJO6ZcZT/Mk6uMToT3C3cf2LBv7N93jjQEd0uogoG41D7kuA69TcqmedR/M1+Mx8
J9n64Fy95OuyjuhXouKJVs2irJOdecRVXOucR11LADB7m195iZkOcnc18I6Y9ZKHF1QnESRnMavV
wDOkxS342UQEi0jcRtyExajCbjVZ4r6M+8QnhVgfQe5rh+CrjtTRDkMljeNOR4GlJohWRRPlNTTs
zp0IbLVdiBbW/hmiGIuyJ8Plbs8nuqQWf9SUnuAg3YI8XVrnkZGcrdR2Aa5X9q5r+/0iL5xbc6VK
uqscCseboFeIeU1wHSnw5hawGOSLeVij8xfdVvYvgIUDBPzXRLsRRGRM6I/FxWjC6ZmV3R4gOdyr
GC8w2LITFQ7H7GwtA4dJ/AET7dVavnmz8MmoZIHfJd4XN8JlPgt9+SBU11i1swFLmnyM/YBrlGSj
Tk7RCl15+oKtXzAqHmh+NFVIWU26AITBZceCxewNb490EO0AR2sCbDfXhEWuWMdn4QGoVAgpQ/9y
FodYE0oZwOygYWLEcudXMVCm+HNcix9qzMTQBzerUlNs7lodbHFO2q086eQbffQZe0F5+2F2L41B
ZaGz5V7MEd1a4tHomSlPRkNWyRJW5eegAxKDwW2PTB6RKCP6jjlYKLYRk7Oo4og3xEGjDuqrw7AS
1Dq6aFxE8l3SdrK/hMlGJm+edA7RfyyvyHXIEG+NkuUW1lhecfNBtN2Eu74e5FVYPM6l4w4YzsWf
Ox3UIT+fX2JwYlMqvwqbBw99LQuPPaj1EnlIZvARp7+Rf4yU26KG97/bW/eVTohr2EZb5CeppVt2
1z4SaGb56HmFgWpVScyYb/zUMbLMXHihxwG2wZCAwt7ur5iPojrb32UbB58O6/c2qk8IcIW8/J05
HLLjY5fBia5BuHieAKJZXBha80C1ltIVkQbTKqf7Kq/ttoFZB6q6aWVgfkCjOvvV1qnN9Dq9aRgq
u9HP9MqY4xl0NBI4BysdNAvzmVOKR3QaOwI9h+uJgWEcqKx4towOkWx8m+lwliZ5nCsF+ZQY94kd
xsbYfkQknk/F7xvet+/slhy+XHWFB5hNQgR0jZQmnfTQxabeay0lhiVbnoOCid5Dj4Lg9dCpXL8k
V08v6Z6wNFAImwCcCd8ZTJ1Aau1q8J++jQhk0RyyWGBCJMx2IOFpJc3JiJCgxOOjC5gHxCSH6kQx
aRsnKLtz0NWDZUdVQT/wSSR8AsHeThvatERWeA7T59WZKQsEWARsbaLI/jw4AKvSF79Auzhve13r
9Rv3yS8MXpqK1OhtYje0rE8HbQGxboJKTt6p0wDyRgXOE/zqWKHs6TNWYcwfgtsSWPNJiLj150f0
mojlNi+rcgsuWow2I0Rr2YA+33mPjmqdJEiYosUESnGBASdyWQeNzgU6uHVOJv9SFRI6DEGIJuKF
wlIkQWxnAYYJZGLsBGILoMHRXW8Hgbw4vaedxWoa90fsrz+Lh2wy8i+YAcpWxzSnHNOAlNWq5gYE
9fn5k8EX5ltzol317nX75Vq03YwJNf7YCmKSuXngtD+ceKvbr1ho/BwxxpAkOdIq5iTVnYu6fmtG
9t83jlvu3R0KmV4eD+5RqxUMrmwM2RA8+hmWFiRN+GVzdcLgvcyjkr9UEBO105X8XwJcGaP6IwuJ
Ksxz3uAkXF92W9ldcGGuM9ujBPc3xLfIJYlDVUSZaH+TBD1JnxqMxTWThl5ptQ/OkY8BqLL+ImKj
mWcDssaRQaUVeu9Y6dhBdQ4HeTSi9VHa6PidYpcASMqk3V9EX/WDfMcNWZDdLZGVoHWjQjdqRF9H
69kvRa9oFtWdQKKkZwaUGnUBqJ4k+SjUbJo7FTQTTQh30ttDyLKYPEemmI6XeRkitkmA8+M3ClCL
MScKxLRWCQtx6P31PMDTHUIBoutbQ+9FkfPPbn81zYTE1p9S4uUysqeFV4iH8aFMDBhT04k2LO2A
gjBbPTOmwIYyqTybbulCj88UPFU0gVo4FXPMtnZb8MXbOaRHs5T3nmdPDB85RX8mPGaA5p4muuI1
2ZSW35Hf+e0XiIAhlgfVQMdkC4lurJZCVjj67sZF1L2vQveJmXucw7mGzgCwTzqbTo3yraGIlLa9
Qg0lUWfIF1d4JCO3vDmGy/75PmACKBm/GoAi7esjg+4CjehQPsfzsnyi00ag2K1gflZIwbr4iHDs
ogcqMWwXrjRnDcc19DvkHs0KkTUmz5167pImCf2YNNqXeoUqsOR7E20ITnU3FqeQXZJuNd5ZmXj5
jSn0IcxvpE5XKVdBF0gccp4rMrKlmpjSFzA0cfhDVwQpcEo3c4+nEjbBhZ9DauV0VGNWXO/dItqI
Iz6OM9w0bTSvPhzO03zcI9zHHolBDEjCnTDGf2VhbMLz6Kq/m5R1jmo2E3ErHSLOxibWKmrqNM7h
vJMi2Uhz2J7GaIpel2i9I+4YLm9/8vHnuyCAy8M6P4uXNx2fOUmVrxsrVVrkq+9cUou1TxDkGwCv
5UdE/s+/nVt9R0D3qQp6RPo85Qcx7QG43KQF+CKFlxyfD6DJdEl3yd5CcmPibSfCiwz9f9SXtEXo
QIFm9uvNWzuDdnfbd52AqPnJodCuq6c/0MG5d+YGtESryurOfzpCpV1n8j2V+4i6y7x8ewCLliq4
Rp1k6I4ed/mCGvsVuZbVXfZElMSPF6KGS3tgVQ+gBo6Z2gwmUPQKzD92wqOc6uT4tHPInr7SgpI8
Gz6a2lz7Wte3+woT8c4OhVArJu2kbgfizSC6fZEizbxApeZL2a8vt0/vLLYG8UNG9yu4rDGG/38X
ZmdL7WMzmiimjh/TqUpyr3o036u9Hd+oh92Zg0hAQMUPz1A3cHJiW8tzOYjTEPP6TpiZ2NKgqVTe
jdPtkBOLwl9K63B7Zop+bM/4dURAWo/h5a9Rf8j4Hl+Qsti794FDm+IIDvSCreigoB/XhRHN1e1e
1zH8vyQpJq0o0zSsO2uNNyQQgV/cMZ5JXoYSxgcuyB4mYibv+fvI5qnNW1pfw722dHkkhmpiWCYR
iLQSmPcqM2igdSBu9WE36k29+mYT73fpe4SSiVaaO0EwFhhnnFWUq3JT6+j9FVNHzSjl3XOutd5b
31S86RfwOptr6dkn3Feqr9FfWh3kSh2iF3zeo++tqboNajRFBZsTFxp5Su8eJ+aLaTyhZSH1Ln3q
OLUQcxU8yS39O+4IH+QcENdLfZybd3falVmL47DV+DcCEQGN1LG1rRmg4zGkOowcm8VVAB8bMUF6
SleJU0hRuHdBF+GtE2BUOI60uiyw4N+8YA8qy7Kj4yk+g8lXjMFQXAsYzp2lsJaYumISXNuWTsHu
Cx/763P0bNuNTknr0spBVI8F311b4K+NFgGAChAOJ3desMhoo7GfPAE/YRV0CiyPHS47mgdXm5kp
jbQp+g3l1IHDBrTtZ7aKehE2/onFzGAM2owGBgKJRnii8hFiyHa1zU93U6WRT/qYnDbI1ZYZRuWy
lmmgBtjpcg736Kq7MkkISkNLioho5jEqR+0RPoYBVIb44o+Jgth4c9eX+oowPMXdqrMqVgNg/SQv
D2/Bi5jjK0J5QDgTlL83kgoD7EUEmeN5HRg66qeb8arZpVGctEwrLjATacrTG/+PgM4c2daQULzF
SgjaY2bNMOYolpukxqw+fPpL2cqWTVofRMvILfg9WQIZUgWRjVD9d5TFnFurlTBAdVBx8OPBYGto
DLDIuuuUIokt/U2+tqAbibmXOnJoZuLqCKJRrSVlWw2COaAim32qhSuUMbrgDvj9MSLclLnmxmYg
PmDX94vP+a8L4/40//kYOL9n/c8/V9r9n2cYdL2Azl5Rwvy5pFzUBm513i1FFELe/k+F4p5aCF9E
3ht+4m5IDa4XDNxMe0FAlNIG20ZTbZQFxs8bVIrMQJCdRW93oBc+nA3LHcKzWChLRxKMfbYbW664
E+ZXm3ovstXfljtHrBHzCTmcMlQgjZRxwU+l7KZifH5xOs0wkPSrT7BGr4xoTrhxL8/K01zGMro5
frRdkjt7NZJ9UOAMpGDt3IJj2KuEyMH0oTExVP5nsI9HM3kNLg2PpnTrPGGxWZ86zHLWZI+/EAuB
97xHZPtpMWmt8xiHYHiiwx41mquKP4/1HBLjrd5m89uTcQe4USyhvC3Fkg3VR7cyAO6/m/Y4t/fK
Ez3wxYW0+IzbqPhMCeoxIouTKrW5RG7dt3bV9fZDjny85qziUQ7S/1sdzvPLmTHfFhf/yQw7bHON
srGZCoUl6kW6qcAuYNpLVjLEUMT6ogUHzNNq9ZsnNL1zsRMKShFp8sLcwnfl5KsEtfjtV7hR6psa
qBw3q4wBQQu2eCkMq9EffS0mBzY7ozSvwuuiPI7FBPrtc22cjPWC1gmmCcCRStDidTVPkpK7HrZo
tWJONi4C97hLUYOgKctKgV/tH+aEvjxtNrLWBF3dTbflioXO9UkhNPZNDiTxgJL0VWfuKhngKmNy
JOOZTyocqu4I7YdQCHSVIDeieilYUwXKYP3x2szYL0e9B7GRGZ/dOZQ+FhqSkG5uq4IF1CVQnARe
Vyd+bK5OUMNKcuNCgx0bqus3Xn8MBYmTIW3iuLdtGVyKlbe0LbLgPj6CmEh7Y80DSKRB+wFaMFYi
fo9JZRAR20cV3diCXeJZlXoaBmzZXjdOQTnTB4YqxFjOVOPz6/s/3gbylfJepFEav4wJdtk4ofFh
WHvjkfhCI4EAsVaFk/DIAq7l5SF6M8b0JEG4U5s+zDsc5mDJRyy46t2+Eo7K2ea3tOQcdEEJli6P
p6pz+1tJ1qHJ/Hnji4Iif+skkvFf5VSwff4ZDG4AcU8kAFWUlnhijsWByIwsG0jMJ2adnUGvVM87
5QDyL9vEo95Jt9mIzEmXlkIo26Xu7ovMPBW7RVXj3K2ocZwudX0W6u9IS0u/R3g1K7kvwtgqDiVD
PGjDIJpPdlKfQfzDGHRYmntPMN7ST9DWST2ZEJMm8dqWpNF8QPs1EjBvb851JBHSkHpVYl1PD0ab
o5oEa3tujilP/+KY9g0Vj8tusRsuJgqXnRV1+o4qPSReHKoK89nuQrP7vt4wleSMjf3qu8hV5MA6
jzEWBpzujKhl1M59Pa+O/nIjmAxcJ8qew4Hlsjcl+x8p65dKQadyIzA7xTOZ+frw+TzQsbClKN9A
O5YTvw4Q/koq9F7ksLDw1ykLYTgVsH7QAHG2UIv6MRuWzUkICAvCo50fCSqud8gRcF4wKg2DZaAZ
uFz8T/2Cw3K9RSG29es+ZE6ClN7Y5HHDXpfCQNNBc/AttzcrhPnGvZ9MsOLA1QEJoiiPBh1X/tFT
hJZ/FzioKAmVK2F8pNkvLLsVZnQYSiqRYer9n2O5e0fhdqDYkwjBtAXRCqmVcQJz7uHfaBMcc3Rh
5GYfwOykxHdgR+LeMRKyMXzeUu2zR2+2kYMdLrDulxSE9tZO4AWObiz2hQq9acKha6qos8remDA9
y5VtaxR94TDvQCCNioVY17p5OKAFBBGyJ4nnREjaJYBka4liTL3WLUT/CZJxZdmoIwVxIVeir0kU
HrIDianmU8hR9ePV6AXZCsRBQowhxUbUsIvnrNuZyDpea+B02BqF92CJ2SB3KPOkyZS0srZaQ9fi
pwXNrXiNsJWR2Yj2JyeNUOqttQZDQFLEMEwM3SxSv1s0zXYgf6EuVIzuq3X0GsVc42GUR1Ql+ppl
s/VYXHOGumQkYz4bEymwJPZRh4OAZakkHMcKo2ixkYGEI050pzrTufjfF7ypyZ3ZmOZEuadRv1Ru
UT6pzIucrDQPij/h64jVWZmS0BMb2aX1jRHtO2iUfXwwgzNyXEUJjeH2dW/HjkVpikp4ymOUoM5O
3fwk1PzSSJjbFrQ+A32s2G43FS+uhp9cLx/NUkiHIo/DcOot8bvC1Sy9j+BTKuNYJJ1XHORRBvU+
tH9taY6pLfrAvdsd09WJvviWzHpBsqmmkLEATKnUVAipGBEtcUU+dP8pyFS5hkyLQkpzb+8JRwsE
sdUy0rU1JSlaIkidSydlj6lha5ktU+tJfRYpR8Vy5ilPOOI2Q6uXhHJ5W9PgzeO0/wSCnA2XWaLI
rhRt0nNHd1BlFqJUlkfwlqPfAdezd1gFRLv7iqzSIwo9vc7bgoyWUr7LU+2HNt2uRJaPtuMCnI1D
1RGB5tIp6Ekn5XNywBsTACiaC5OKIljtG2lqAW7iWZ0qHQ9jXXpR09YOpo62WQon70TEBMQ7NAa8
17Ef/BY2HIPKgVKojS96KZ0HIifixS2gW06YVdXkZ1/moyaNahwfkbWztIaeaN7ndZggnwzJArXB
OC3jRbJ+xz7+fByty3PJy+ByfSxo0LF38P1+X2/7WlVPRUkSYG7MZaqN9eE3K+rgRpD68EWzCL2M
firvTbx4MKSV8zyewyItXrJ3zWyeObEaZJ4d2tHSni64xGNKAsUEMzpBXxDoFu/LSHw1Gl/dg6v3
BodZAW1qQ+IsP0SBBHHK6Vi5q2rWsa0DfAP1V84/HlEAXED1b7RTmKH1uwgVSFpfDYhSujGyCNdb
InTdDInqJ1MQvJI9X6IWrMUwtjkPkSZ8//Yl18l9Bxm2q6I+QLuWbEOjFmE/lcuyD3iNMvHH/PIU
ejNCev6DrqJG2YwtS/vy5iZJa9HvPbUGNqsSZQ983Aun/h9qX8g5bchuxo9VCbI/mixtsjaLNbxk
8w+Mp0eG41GqZzbVf4H44Wrs/kDM+6yVUDFrFD5C9D4XyL+XJrscWVCN0zM4/i7bwr5uMaIcuy6s
fHKa++N0bG0OnLiSamGISZTait1iXDK7KLNsIHIXzXPm28FcWmjHQys/cvdjOHXYiD04ir6drfc5
Qe4xuCWVTRJbAX/v6w10bfjCfu2Q9lahGVImnp4oD1ev41YfmPhdsqhk6OpbzTipGlw17y3BV5vH
vVvSqK9IjuCkDP87Vh6/41MpcrLbSkZ+leCCQWdunyHb4zND5M8BToj4RERUkMniyxC/wArkKbdZ
0RRQ7zsTVVs3Ty96+FL4HOIgfYY9bL1A7Pled2wp6Il3N5IUvpuDlCBdfp670jQhggVX8Fbinj7z
5k5gK1vxrCvHIAqatbvIVZ9IcIpO0uws0yjPWgj8yN3edDT7+67GV1ziJ1SdVIvrTzmV7cjWGQeH
SuslLXiHxNUtw5Urugw1O/ezF289ojcviN/00lVUkdpw/PRt482BbGuvJV2SZVdxArzFqGg1kJtH
xlvHk2DdZLZ1zFD/sTkOjVq39/WfmwVJKBmUdD/s7sjsEeGlf2wBvqwhx/rvWycpjECK+FIGKHuw
wCEqibQwnQqrxQgzXD/sTscEp8viZJIgEO7IbUtN4xbs6gHIVGQ9AC9dkUQLsNlqdRNGNO8nRqIS
8klzZ5hzzkgCTjIU5ZdhoVJ+/2KqRvpMpWDhj+srqHgTicKs+IAPHp9hwZhw9kYuUOCpYtZgLopF
Xu+J1E5OgJg6pZzh48Grq4SY8WTs+iHDJqM/E4mwN5hpcVI6dwbvszQJWePMZy2ltLklVsyc4EkN
xtSwCsYzB5CTxG2aWniRsKN0OPYkSMOQ0Wq9agk9nvPLPGDPzHHx6p5U3BC4gwV2WLn1tnvaV6aK
CMRT3KWSDeU6cO+x9fa9LGmo2/ThZZBw/HVtbPvsLRg1aEE89xHbLSc3F4nBZ/hm6IvU4y+fC4jE
Nh/AkpOSOwacWfbizslD9P3YKnm90waCxEOh+tgZ5LTFcc8+VAXhYPaMh3pT2mVZonVBMmC27oaG
74kfL5hkmEY9ZrTb98rkyEF5ZItYpyDTMizbMCk7VizUYCdd2FNIolmTvidxc+gqJeTKwqx+XlDB
fXOI4BoO3stW0xsdcs7f06z5HcsIoVzE4ZvRyVyaSUxaKpFBKxE8Os9ZOuj6uRXth1rMpPZs445f
OuO76LX3rGY5mcuo++u+fpgv0qo4avoWJmIFTThttqu08PiMex1VPpAlJ+pzIwaKnLDlGzToeFvq
F0/bCHOO3ytSC1pNqlKEOHdLm0MroMjn0XEwXJj78sxVxiLpTtfkvq9nNTtT0k61c9gZvNGrb1uK
eNUmyyl/ztg+p/rMtl7iw96OuNklTr6Ks6x11Xi1x/521IzKt46Z1Be+rGkv2YZi/wzm2OhRXYzc
87dkONLwMDDiWB/ILAn5rwmzcKfx3eEvm5xftz4nYtUw3U8K+Jsi0QufvOqOe/65BXoE7WTxFHo9
aEYyWcXjnSY9VQM6Ld0Aym8hAhjN0izMVYysKmmDl/PfYj0GBH2ILo+Nz9myr+/8VZUi0EMC5ZHk
8ldqcL7fLWghigTYF1cxlr4wU0EHve7Jjfa6IIpQcZ8YN0mkQiaNuUQpwh+1cBJr8W/Q5JlcipzS
ofNkCEpCzweZJmnAWo3TmaH12TwojT+Sgmr5EDhCRCLKMaCms0eBAe9illCW356z5tFapanWxMCh
APs0kfyDwwuoZUInCHuC6iLeGrLABxB/c0GGTMK0Q1XkvwZODxpETLiQMvI/+dJ3HHKwWKRf06zT
Gt965ilM+q74AfBrlbqEeHfFv4fPwIZ2IR9SAIhPnog2jvIel9eQ6R9TzHczXVGGV12CNwcorAUy
gb2FU3OSQ6s+2jfbdSOCveDkJv8vMH8ZPDhNKOKITZMnyG2ialI7bpol68AeqArmsBAK0peWFu4p
6tGOGhfbD/n6f828B1lbpQ150EKVLuU3KvfqTF5plVuXWKoGtJozhUjm9bTbksWH76Lbm1WSFQMn
lJIRZDpG8xS4OdfqjZqalRrIvCXsm0Scs0yB9pEFIqJOStw04QxeC8CV4pUslo0sNnomQE5QL0aR
hg/t6topdNRPeQhNGCbyCeW5q7DiJ92ntvXAYtWfsOXIbJEyyBXL4QjzClQpfEv5E1UIPQ21xEJH
tJ/YYbiqFoLftjExJU5jh/4Uyw/zUT18Ozgvw0migdn+97mDiivKqbNq7l0Pw8z/f5nVQ0DoSPAl
P9knDXqph6FzEDJxo/awoalaPAHWe+gwERYUdcJFUIBL/ojOn8amYkijiApsHdk1gjChUu1iKJu/
5OO28OAxBcPyXKZvBv2wXkGcHz7QLiBddQvew0srAzjIx/PQzsYqvZDYopSVyg7WXnUbEZqQo73B
zbqKRA5e+N6kVNuL/4RndbKaHB+qtSspPAauFPomnKdOStYADLKUGegr2mKF9+bp8eXxP3cwpotV
Gq1yttRHTPUwMTTXmgdILCUWfTApTlAk5anOdmZi9dqw4lLoUJB+aLXHVJFjajh5B79hUws46pEN
A1OghY8Ln966iAaei5C48BisW4+SSzwn3sZ5qXdg/WpM223yJg/DEEtrRPCEnUR6qIMH7b3w6t9U
LB6QIXzfqLXlQF8gb97w81j+i/GQDhLlhVErPEHBZteZW/8TiGGDWAEIApV9Cgh6owtyhnt5JVw2
cceYm1s+OkUw5SQZ8TxCBlc/3nD7HovHX1QSDCumhMEACCZrKbgyvm/o2HMKCw27XgBaZAm0bm+x
iBAJwaXXhmeG3P+RNBtbTCazmHrtIQrl8unjc7cZQ1JRRzYexvTrkmER9sGHHaHMGPjF1dhje/5k
hmSJgChF7/ZXvvqCIXVdo+crCRZsGAjzIDxe7Te29f+jq9HLBbh9TKMFGCGZZdhLOv8UyaQ32ql3
55teQUNBmgGaNoFpF/2P/Hg0foWweKvyBq4tOk2FeY8r+ig3kMcGbVEGBeA3lA+mroQqfxn/pYjp
lp+HbW29CQifD4rbGOsBMk3XplvDR/KVgcP/ariF+GrGZImsWk9NLw0SorjyimrWlVWI/ZCODeOO
lDsh8XdiBXQzApbkWSVwBZGhBtToZhkKAsL0suvk2Ccd9Lbgnp4Xvqr4Gf8FfCODWrnw0ik6Y5nu
Z2ZZuWGSXJUJVu4F6tu+2TCvGwqvk94KPVFIDKN7xioqGfBrT8VZPBPU6Wf0vZx7pwz0ROieDs6j
9sob1NClKxsJ13lwnJy8r5XT7GA93Yvm/Pvq34kjwK2dOrrfyYW+QS3rtWnqdnvu6KhhrX7L9pwK
pfvR9AsjyKmEC+xOvgnKGlTrBsJpuHLBJunEaA75y6kXemNy5tGenH+hNMS9UTNESIq/HJs/mhn0
BuD8RL0YPKWI3Y51c/EsMonySSW8iKNnAFbV7lAv50fY1nPi5tQVjSlZ/MRzJRjnF82YEpxvcqro
1F+GGi5ObhAfJXx9MjZhMraCciE/aBYyYaZWERr0jeOxR8KiJ+WnR4rpVdA25+7nAd2dlA9QAP6L
Fr7zbFMqnDugXEq9QKR7GgaJXy/0YGBrf6EnXo1a1thmbaHI4aK9md/7g57Y5sscd3HKu1gaBoK3
Fd4Hf5n/TB1ake4LhrT5yqp4P3Q2msY/ZWpXwzGHAPu+bzyIhqRBHJ5TyIfaD96GtqTUhQaqY4RU
Qouxnk6OLAbB+Hboj+vP1POeoa/IosUpPGUjXwoWsKk5fcQZfT636AGpCGBtfAnWr8bbUjDVAh5h
qpmQuXKwDq4eyqLGNgNjsb0N5Z+CRiXlXHjcXGimk+87F7NHO5UOSs74PyHhJDdN5Mgwc6WxV5F8
IeY6TN5OECkP6MFmEUxc7nUyaiqAQkLwBKpLo1wYdNlmjygp2nFKDCeIbJpbIv+12wxO5TTzm8FI
WFUVIfgccUE3BgcdkF6BIe7zlgm3rUMGi4fW4qrF3f87W0WIhlDh82DbqVrhT+FLhon32XELbNdf
ZnGmhFTjLFQ49GEJXZl9XW9b7AFkj6zFWgPPT/+Ow7CG5PKrz8sLg60Q1XI9+wyW9rRBvD040mVG
D0VjunnImpu21PfSxj8I0DCq6kmsJrJraLqhu8znwqad/xCO/jHmeY4Vp8xb2K2MyKv1v0BIWaA+
xNaBN0GrjRsKE9u5tCmPlT3qtLJnWl0VzkS4SQx2DGbI1VmWzfsgLyKbjdqc4XuVszTyZJvPt/qA
9AElLrVYgBJC6IEkHVRURTKWlbF0AqAdu2N7TpqIZ/1CV5Ang2wRpgG9hmkVtW8Ir3ZbIJDlOzUz
R27Hl6rc2kxTPkUt8Z9ci2aKbDAV8Cx8Y/2ExbRVfDm6+wzchrdj8tcbol+4ol7eO+7n4PVApKYy
fXM++wkcZzD1w5d0jh02wBmJ2AwFfGnJZ0hrqppmnpv1WAmFQx97l22SX1mf39nNLK2sTQ7JMk6G
JUGXxkcOHynki6tllw99N5N64CINcrlujGr2pFXMUkpoYYQO4e5e4yAtIWm+H3LZxSyO9OZ//NyW
L3lTV7mvSUX/e+Iy4EZg64wljkw7JhSs5L9qvak2JctUh7a2k6TcSfzj572FWCkTztci0qGcMsfa
sxCqBW6S7jD4V0oEq5OV17vOYqaw18r6w99tJIoAP1mXEwFooKFd8JWqQ4ZoeJhIeDAYC0q0s59S
sT83V4rhaFgSdxnV7zZyrh7joaBK/wg41B2Y4wBIPPyc4prSSIot1c2gUX7CRUzA38ntcJRgwNWB
GN8Wgx4MHnpGncscuoUk5pOWtCLAMl9pFmSQ/VZ/AasGSkbAgJVjGcrBJO517j4UYSWVbGQcNQRw
sGS08yd15OWEfYiptzsRdxwXeByDn72DWuTAbc6GOWQowQpLxv0cUaguKNzpNxZQQce5BbtVY5fS
prXnLot7WSHpDW6yGf5srNJPhW9qPP8SJIyh+2fMGGvOvlL+YBP4puaeQocHySB9OE7rgZ7vKZAA
A8lpxoJ5DfSZr6jUmV+fSGksjSurHMsH27cRh4V3BH2xz7KayxtvcX6BADoAQ/wu+r6tjggLIouo
K3yq+FDB14U5SeOqFUo6ceX1D4hA2WQ3bd+8oqGeLoL2Zdeyp6aJTBpQ0yC0/gBbAURGeY0r6aho
+2gap6/cyAqd48RXpqzApa+zLEFCF6O0RBRm49hCVDNi3PB3C9nmdA/TuGoXZ9e3mb7r5yYhNHzc
VDDIK0EvD2J72CUK+mMi/UGt3eWTmwcDJZdD8yDMIcwhdWra1sJauy7EGKuvRredf8+aMCjT4DdI
GsI5ASfPCbZSPVGqub36V2HwViDhNyaUHNfP/cWEmvgh5IdsEjPXIl2o0UWFA7FOhQoHvv+jgQ9Q
q7a5RLnNQk2zO9anSNdlvIk3i0XWREuSNa/awVOeBEMger2Ff+bzuzSPrucaF5MmRxFZ5fGj8WoJ
S66wXJFX7dcu0lBc9nZisQhdNX7nbGR3AIpcWEiVnFTohdefo3lagrZeIuJfoomhuPQnDm2ZAH1J
+kfMXVWeXgLIgQiRd1IeNFuH9cgKr17yBb/1Z4eELqHtJHosOAOSL6MnH070a0qbCF4ycibpE6qV
WT/HDLbBQ6b+qxSBDrdgtcBaUH0bFTHF7VcvaApbboqd5ysRqZYjAc9dxTj3tbUw9W4UHUI8GsOG
SRN/1Wqo4Da+MTvQIL8P52suth1cw+gXtJq6sEZxvvEH340ePYgWGQ0KU51EXlxSBziCF3npHp7x
20VtoJc1BSfQieImNfolJwreswqLeKnEoptlFMkZMRY3SGKKpBwEjYGjW02WJf+eYZ+D70wks3Qh
YBH4jYsEVi+Sg6hn49R4ytWgDJ/o4eMaY7lQwAAjdPCRi1sW1MPzSFF+CrxH+mj0Stt/QsMlVroD
k/fdOTQIYFvSQ7PQ6vGS/xS48jpl4f1IRAYwA1upoTwo33JMAplv/imAMBJKUFpcrHAowRvKyXbL
HHCxUZYUpKzza2BTbWvc64Ov16d0qvKa2wAD3G7rcs+07ycZEsj/rXfZoFcUOhdgn4etOLMT8xfK
7TOhf1Qyw2gFXIYRCeJPI6WwxP5TR8rCn2Wh/ix8L8Fh4PszIf80zEuvMxX+qDZlynezatxvteJ6
/bPNds0ngEc2NxFbBNm8kSBbSawSbqbeDqHjSVlpkzEYU3C8LCXME4wXPY9xWbCTc7qTmH0bi5N9
eEC0PoBqn4stzCr7zsBc9pNp5fVzI+XbZx3tC3daGofjxf2aOwL3EqlKa15I3/AW+bssFijNO/2n
Xam5h7vhGxIDBEw0Yhhl1E4HG8UJ+ZvAAQYl2PNVzY2rdTqOW1VWrKeasvir5EzxyCDrKQ+86TUh
L6TBdmQmrAziSXoJxViy7/9jw2TUKLnL0xRif2peTPlF3TEBeLSqjmExeOheIir+I3bqOVNKBa7Y
JGc9b611rqiKNMSiFPTxezbjDPxHVeu68PhhhAl1W8CdwRw7g3Qco4lxa4LYncBzEHXprVxICk/J
a7G4X6DVnJ+lciUQs+Ux93E1uleK7o4ddaoK8O7Jcm5kpTYR+TY9Y+US2L1wEkAlvQMoarIIVxm2
AYytqG4PuIFLamRrKnLxzS9tXY18BrkYcTO5Jc5a/BNtxdv+81umq7iB5GmAzXY1RvuiW68M6rHd
YChfC3qPJGHJJ3Slt+c8vEfFXi+fsuUUJYjpku0GM68imrNKnygQqLcITXnpQbw1L6uuAWSgXwZB
zjsVzB6lGIiFnj27IMUjj1vyGV5B6a/BCGhM5ppu2Ex2WlDkYLbFF09OsV99iENClh1z+bVDsaIJ
ab0bsL0Wahg7O468rhtnX0Dbp0Zjq0qvAFzAKQ6ok1Amr4kTt1tQTexaQ5cD/JrchvgVeASH4gg2
qDKJSoR039k+GspzEknU6Z2OzTIfbgyI88LMfoxIYZJaqDgo76fKm50OiClaYdF8vD98daw9vrVU
EPokR/9UyeY8K0r3/1VSOCtEvnJA6knwHwZ35iPNRYGhwYuqUIL/jeljYW5Ds08Yfe3s+MW08gNb
Oven5iSCx9QVGOz2EndYq8nLp10dt+60HwI3KwBdZ8F0Qcq4OY8z6xgqHSzKOauG0tAQ7Xx1nr5b
OU0lV0+wdNJPGhO9C3YuvVzc8i0VEtmR05+JGAeAHJlsxqNEUAYfc5s7NONJId7eZREvoIq04W3w
Tu+190pygWjFuJgF/GfJEz1VfVYinJM0mUDrF7fM3ovgzPGx1AvU7SG+sX1fbqN0WHAdi+1gj5y/
cY0a4RYJC+1b574q7QARMoD/7tlkbpvxi8epkwDQTNy9T/d1fCbHqMEG8l4Ad3Fh1/zoB+/JrkmA
EYLEjUAPQrzXU1wQn1pYwe3hhbb7gBsWt/bZ5Hs8WngLgewmk/TSKdamu/oPMhZoDQBiQrFwWnYW
HC+a70RW3FAbs3dhdFTLmc2mEMG8fXZARgf88aBq/ifJGf3NnWPX6ObWdCC2XffZ/W0b6LnFD2rU
d1MJzWwmQM7K8zkwrkKUsfui2FJ6MalsLEymamCPK264Mnz9+KvxPxjJzveydm6ZOumVID4Yktsq
WEq3zi1HklXhkurkRsBJ8yERYJt1wg1FsHaOBKBj7WzAoFZ3JsfHF7DU8F9zGIf2FRn2llnYXHO4
Cg8tSxpzjemaRz+G/pbsMlTTZYZeg93gO2QiNPDgIOexXG2vlbMas2SjSIFo1A6d1gqHP0LUcanF
iuDYOu0ajxiP6U4GtHtVts421l/4MYUfhqVAv2RQ2Qm3K35dycdVtu0xxQl0wkk6EgndQY5wf5ZP
ZN6zrqL7c0xp1xYtDQycnLu+IVdrO0+9vyGYbcfjuZSSHp1kqXps94tlKhhh48MSJIY1F8EoyEdF
HO+mKpGjZunQ9dnxmaUSGAfrbu8royc1yc9Dus7PRceES76ULIgnvZvZAuhMeFbWzh3KsKlWGn9Z
US/3nczwp6hhaoM2OXd7tYPa/EqruoVSsgMzHKqF7dg+Sj/c3U6D5tZlzPl71uCLwX+QV/cb5XML
z+EukDgLC8d/nIt8RwxUq4WitFN3DBg6B1ySZgFSWVlSliN876br4J3rRkkrJxICfAtO/+JItQeB
g9rZHDY+nJTg9vqjFwAzMoZL7QBpZQwFULUICHBIoTqUv8pcOkoxSzy89ANcTb4C8p9Iq+64Vj0p
wxffPsVbS7ZVn7LM4sUNL42pDhmElW472epg7owVspUi7f6cB34LOZv/g/Pm1dI2SiuD+IwoxJaV
E20BwSw+U+ubrzA+oftQAtnRcZrpf8kf0JJQZ289VrROeA+E6FIDZM/L08rr6lwXxR/AzmYyH9eC
pu0hFGnBrSb03wXVaezBeaSqnCvGxPqFhIL6PZLglUxMncUX911DQzL6A+6LFLK14aTg2MNhc5gk
pql7+6zSG8jA/yDJxBbqqwumZvWggbHMK/FdImh5CKrUSbGTvahwrMc7nCLa9zT9PfNMKbnWTwuf
Yc8Te5xNzG2e6oCCg/fX98SlpZVrRePvet+jePsjHFnd+qx55T28fj4jW2YKH19xaZMrmNvGEmsF
ZTKcFPmBrFkY1fIbYgqwYWCvbBatc1N9RE3sP2YjwgH2B+ffz7AvAADwmo7NBXxm7es9yl8fZVCq
+wtj4EssWf9DSjF+wYBdhHcnoH/W5Mt09GHZcDykgAzYf8Pq3iYTb5PtaICBHdxloZIzebGnFtMH
wFrHpOiGIhOw38YPHR0kHXeoqStO0wFRE9wb7gW35FweePsxba9M8+wZGaJsm98g2XV+6lIuXd3o
v9JOzR9L49DxpPTvA9cv163rLwCCBvxyQeNCKWXb8U16hQU/mV0SGmpofqo8FzVFhvpI5grN/59o
5aJifSBiuBcd+RqPMS7LzE+WeSjiVXaNf6CsmXPM0At/QFlPWtJDMFsbhslEYKR9AG7bTkGcBEzu
WiHxGyTAjvm3g3lxgZZWuyEDopQ8aBdGIbhcZzjQ67+nfbolwrIaYcpBGKaq/BEl1+rx6hDguMm/
//oFLhEF1Y6IxbeJO6Sm9n3oT9Jv35Mvn+5Qxa7Ko6J8S0pF6GglVNA/ozVLx6ZFY9onbizoU0sy
uWd+/p84rZUgPtAPL7f2aARd6QTqC24OGpLfDgMFvHm5gubnSQo6Q8aP2lVqqKSHIbIopuj/tLZE
skdwbkvs0QqRWNa5sY452l1NuR3iplC2liJK4wx0SNraT9DuGomHbUtOyT6INvDouB5FZbFfQPZZ
Wmzlvol7u+FFBZ22CWja5C4miF7brhj1jX3JwcfaR/5haNk5beQLVT7VGsJRHFvmlTBG9NmPwKhH
818L/MxsamebiPJYpxSRUHagaggbOHpYJ5gj1BU5bGzQRvlN7M/mJb3BH5lvapE2MKM6wBluuVev
orEQnbwOR2XwPlLLmA5xMKTejZicACF5aJnArUYPcaOpFCecaAgcKi3p2FGkVHBYHKefgg0syqo3
0Ef9ftmqFKSzwummoh19Cml7FwA4Vl+SYSEixcxjAFDP7tfaS3LqC449s0YlGXUM9lX76nMh5ROK
H1GEws1iJ+ACdIIKpaeuSUbMdbAwml2aXOCrocABMTAnP35211BbiteHc5b311A+7jjwoITopCrd
EhKtjdamnRx95RoN07U+USQ2oalJMlFi/cSEonJnjkgOr9mpe8iDqaslAi6VtmGltjrtWUDnj2Wo
HKNo+9LuxoRpD0uegd882+w/Ef5uEkiFwHu/NfE1N8+bmBq93F729mCFUI7xlR+3dSLLY0QbM0NL
3cMpVt2z8+a0FJVMvyvcdArDxf7AieGJ+Km6a5j62KsViM6shI1kU9XgF8RXq2suPqLTVPBJB9DN
1mfRIa2hb5aigNBOw32zbe+RIBWgoqdwZkE+z0FNBF/F4ZW5925HSwL/dYq9UkKb5oXA5qhAkbWS
Ky5ZcoysTx+uS1Yl9A82Nnx/ULl9spnvCKBdlEZD45DaRPUQyMNBAIQRJZHlRxUxDyOxJdIcSEmx
QEaDOjDStvkaVJM5myl5wJMZmanPyihKiYrwbwE1gqADgIJVCrP04176VUFeh4Nk0INi3MUOilW8
LYV8w6NSG1QK1B+UxcPtoVuKFTuPXlc4xAIs56vrT5j/40nQtKX1RjFXzx6K4Svu8vI2Aeej608p
jZ64QI2H8L5oScP3s2CVKHbucW9kVOivNli+IAzAAIhJSmicP1d6fkw2Xg/FbxFL3gkUz+de4LjC
twrQMvrEzMZrI1w6F9ua9TK8ayqQluLmDCM6g33hjNCfSKO/IIkglnoOcRJgggTPZJ16vPQG3vRS
NX6v66SNFK+2pSzJ3pMJrdYLkt9OemCMK8G/iYvMeF5+trx7tG4IMW/Y1i9zSpdSk1jear1sWLlv
wcak5V7UR2hhs+ZkaOkZU0E/9HGtrWU5yuX3HyBTXg6HCSYteKVJ9kpFfBpoY1dQJWyIl+V5iqBF
v6ZHuXEN7LJopcJ4L2KG9PswoWvGGoyfcsNdHSc7yigDpfGA01AQ2q9ugmgq3eZDTidcJVSFVrmb
1yjICKs67f3P59LLMFKaMTeYggFCMGivKwwuoGMyV3dfA8i3AeJyfUnFDZjMJmTslntEJp+FZ+7S
WzyJQ/qW7CBpoFowdNw1Fov90eNFlSRaB/oVwimv2oZeRCPD/lDlyiUOslP1skiI4yXkGz0wF/+P
WYvFZBuD9pHQpdCNPuly8pYvAqmv9MyEi0pfcKhLd1KKV7tamkL7a+EN4/I1z1Ig4cG6P2nDqUXz
8l4AqO8dEiRPTuOUdlbqrwQo8/o5po7JJz6PxTpCjo0R2g7brQskCL72lFEQtqKLA+RHg+oS/4l7
vEc9U/8xnfIXwleQG3SK1KykljkF0vJ7BCuY+UGzNEYMXUQpWEkAAC2kh6S5Okic3up4zmxXJ1YR
HOHASTU8g2nqtnsmOTCuRy8x2lYoygX1KVH4a7HMbf7vHELDhX0sE+nypj2/RuoziNAxxrWWwSao
szJPsG9DVOcUaD3vKTKzHyQ4PxYlVeLnIElCbVVSr2nxZZuZ0d6uNdC1NyRBZOXsq6T3fatFhWnG
LZXgvBGv4Pz9Yfm0374O7eJypR0lLN+baKHkLYtfHeJP7dkwmPbP/yqOneUmJIIDywYqrqVtMhTF
xn0X4pSx36sg5AiJ2+gP9VGYFKqW4WgqFkfcU3GZk/GUcaL3b9wWUwMiS2C3HthZ0E29/ZA/uA7F
cRTFrlxAiY+EBCfELvNc+IlnSakWK7HXpuBffsxAsCJ1FOZqg0xcSXRBN4gHIdehzjFtBU95dKS1
C6agtY3TSHkj7Bi6QcVou+DCCzkCvctbullZoPRx/pq2bOgbjQGHU1gh19bpwz6Ur/MtEUyB3EPX
k3uM6GWEbiUXGn98YmEiTKWg+2MTvQPuehGAvPznHKrPddq1LPrlsIU4LdYugTqCnyQp8DZnLVTW
U62MFDzY4gCuI/SuLiuXxrpOXxIRNdignrdu5Yz4oCWhXKUtOveR82XREqZ6AOLqbasLCLvwzNr0
M+b8S/IMtd98sdkluc2n5LQl+TysyhM+I/532a01Bph78XvkRpCM/F+wFnOOjXvs8+ZCdBmkO7lK
wouLgKMIo3tFFlPwWBGo8M8fTNQOR80UqBZaumfLtDZNigLpCHCZXfqrHzh+oXDKU62dRtEIZxdY
7xNZr5saw2yTRa0BmPRMEBV3luEoKMU0velGnekk0SVrwxh7ZFJBVCK75tfgh/j9k7Ok7B/S+UYh
SgrqxdF4BC7WsPhqPwhkDtt8JeuQ/yICMduiUtlaAj+/jRGsxTf9UcqZdI0zEYJ+omaZJgZYE7WE
JC4WLep1WXlNw4IV04FhqTm/0JKDphmxm+I8f00eMJFsfIp68sRFQru+B+9yNoQZCdzm2T9RZjOk
ChhGwJrewp87uBP+dHKsC4i0rAcQK4tjDjxhqVcPBto9AknbXrWI9528aIztqOz8EfXNvajZi8Qt
qmGFcCSe1ND+4xbXkOL0sGm+pFq21Sg9R5lQ7a23FMbT6MSrnbbnqbMbnj+UvAFxlWskHTKo9Fjt
jy12kSCLHbRwkgMFgBOyS5PBZ2fPYmujkt5XKa/WIYRwFBso8lZY5M3ZRWqTbMydxvlqbpjIPz65
BvUIURDFSS1OOrbPkbmtInefbjYG6iBOEgRlhw1FbeV8hKoJgtWpvnBJnYV+V5Wb4AnjWv+fAqbK
9yV0ijjB5/OgfN3xzAQFF0BHwRuQi6Hg3DlSAyf+H7X4uniSGuIZFia7875n8XvBLfacpIf6c9FN
UlnMT2oQH10L14lYhFAEnp3ZxoM0zsir8tVD3iSVFAE8Nzg+UAz8RQ+X4r7oIeh0w6II6jzvQeLP
bx+SDpQuf1YmFukcChDyNVCHjH5eKY9cMj2EIt/agO8knJrGXI+tP14vg/+Gc/bY9Mk5KujWilmA
viYGdg+XYLfadNep4rVHW6MuywtTe459JSlqcnJBkGjQCvXjkVCXjBwtImrsgHBSLIgBdsV6gc3F
AkYvc4LTnEUvzk9LeiAnIrIIRGCRHch8CAVPAkekaXYwSKo+PHTI4HrSFtq1H2ytV4pJznvjJpOT
R+RZ/tg+Pf5ilUz8cse57E2u84iAYz+NYw/y/8d70GA1/PBkQZZXN+K4uQyhORbiIbMVhZbBi4pX
G4+J3Vj3XjfG9abLGh/o550JMjd1ZCqLAa1raS2oHKJXZQHj5+/KyLCIL/SRFpXLmtYQuQK+zxMG
u05q//phFAQ8Ujz56em+aG6pkvDp5hZNil9mSqEUpX7DtMC3N5WEpPWrYYdCD1H0pnoTXBu181yh
mUxgP4fgN3N5YtyaceUyb2z63SKPGkATaNr7for3pKXGBRG4I7W+nSt4ufvk0JTbIrKIISwyvGsC
6RbGIjHVI+Fvacs+KLCSPpJTdgdk59N8r7Fu/aHeNRFmFa8vq8OIUOo8g+oSE9Mmjehdv1I0FYsG
2Kc55yNWbqOCYKtWNZKkMCh2Ge0z2ycamU8hKq2AWEjYJwLJLTazxDyzvHivmu35FgPK+i9977om
nCI5z0JyVr+3HCL6KaxS10E5Uf/byw8ZCAD/155ATAMRbnkFfKU0I6vOXFzGQhrBcv15DNQghBCQ
XpmT+uuQl0O+Lw1jM/XXTvclACcgNmUwL+7yq07bv95az/ShlcjaonrGZYxYlyKeiPns1KuntVbI
t+c+9LGUV/LGwvFkbW2UFEfbdFrrYZOo6VrvJX0a6MS+P0s/QSqbmBqw/XeRQpTxPab936282hWC
eOgbCDuMTfJLwttxZ+hYpwKd9KOA3krQicfEpA7k+V6ahGZ4NicxCZLu4SOuLHPkZ6V8qVCJZxUV
4aI+EHawgIP3aYXpzUvjD7+hJ4VftW+XWS1oYctILZV4z3XtTxOcNpxCygfHdbZET1Ke5WiYAtDH
QJUHMnrgHHsdPSi8+nebKJ282jYeb3YZcXQy8FcIc3H5E1JSggxXgqoee9pJlP41h93OV07V9jBy
9qdxDo4xCOOGpViCpaVjdWuTVrCS5QIstf34/6be8icXh4VbueDEtJ4pBQvTXhFtf3QHqVKgGIdR
aLOsbvlN7OfT36Ic3vmRu6K135vnB/kruYkCfOqz8uA7dXmHY1tcUuizOfRbXD5DjfyFZaAZiP4f
bttEWARCvu7GZHtAVQkfUYJQ5yODbIsigG3AbNJftZka2rFSDXw/6ope6JVNMcJINihDFo3mbeyL
ZOBVBqqqThOij28RY6HmtdMic6JoueleCNJdR8gakXsyUvJsGBqEfLJc7H9+04RsuSvfH4fp/fyf
bvkmJOepQXykeRbuiHgNTw4Ok/7eXkJzaLwWV4Qy1vcjAH3zzBEF7OFvo0NWRcyawwp8WR989nF7
y7PFYtZwIH/UBxPhG8H/xCx6EfXbhnl86RavN01NMeEdMVU7QAJHAcZNJVCcw/CpbQKFKC2etAqz
IvlVRiFh2Mr/vbcgUpzA3olLqq/tVBayhX/FF8SqTmiN+U0fPBEB0sAUWMGFmNINSYW9oDPxWdfC
7dNmRzm7DJ4+6jw3BaZUK7M9fkKuACN0ho0+X7IwS7CBuz5ueBguBTAB0yubhIM5a4sXTTtMmQg7
xfvOWlSUvJoG30Myf3kZQJYADjBI4ImegjI1bUPbfMIeM/sljTu46dt+5DWKwdYhnhv6CEdOQgB2
z1lDlu/foBCJ8Ann+3xYsuV00EpZFRehWDCmOa1psr4YtiYBIsKYrm8mxCXygiibWkwgjhPmTsT0
B9HXeq0JUTNTVRJAwbkt2ydhBxvi9IIVRpIPpd22Xf9zlJPXTV+e+i7wBNdMm78B0VitH+ILrU5Y
sfZ8M6ijXLz3nBhZ8oSR/u4uuqHGUqguOHu3W5WpvBn8ZvHPpp0i4GdTemCDLr51ucoZXL5KKblm
Yjh1QmqqG7L1Vv7NGp142gh8drw+r9WuS9tnvz89wvuPymCzcvbBtaD773GeLgFxy/mVegyFAujG
8+RFVznaHJAyDryfONlRcBuy9jsfcitT1gML5bx8XZY4SzcsoUb77ZprzBS2FOP7o8VoMLkAhgYk
aaLvfShzb5fsfGXvQZgII03f81ab+uZs9/LIP1ieJWDSfntNgra72pQUUC4+EhxuTt1EqjUU84Cr
dFY1t5euiaDsPGT5TKj5uab3341Nl+e0EL4q+0dYhld5pBED60PcL6bPkCe45fRQktLQNSEMno0M
gtL2PnbCTxeXwnAiv+AuHj+6DokGGwx9f2uiZOWucsOWuIW2f2eDqvkcY6zHJIWmT9dpEYKEVk/s
pm7grd6vSG8nrSkee2YdAujKBCyY1sTSYqP30cg9xd6RqXvNmCiS3W9kWz9YnFyOg+I3XqcoSfae
GRVVwkAABAeE+TSprUtYQsnBKIK2Qc7QPxd42ut9VQaFv2Ego+DOVhzzlTA2E8ATePBxPA8iltzl
RnovU6eIEHZ82600bbCOPk30Av7D65T3jWRfPS0F4iUmmpAZPOBoW/4kRq/ndQEQWwUkHQRYTjgV
HkOctKMa0hpvui1vTHph0w/AIlsqM1GN8Ku9ma8bLqXFAZEB92SXHA9quj+iRvWGqmmjfuI1vImq
Jx3AXWiE+cWeU6pxH8jHATR73ZRshTTbkww/6bhkXutYo3VxgiUIjHUmoctAcxEvW8K6kzP5Hw5F
PeDGp/Mho/aqYGbkyLtZ3v23PXZ7xYc/JqcEmYxDPPabCRPGHsc9hlOF8Vd3677bwyuqup4sFgIb
J1YHM+7Y5M2wWKLYIaCD8bwJSTNoOY+jimkheJ60LjnEh8r7/tLuI0Db6bXWZkICqOS5f81JO9GT
EHJkxHCKxY0tOkoknLhdUNU5+anMXvBnu8zKIuiDtcgngou5EfXG9R8nhQrUyWDkuIHN/Y4utW9u
U07IYIZIKrVTxdA722oXG/YJQxwcIbqSuC6qCKmFkS7HXGivNpdiHrO3+1vLohLT822qiV0n9/7t
0lnnCA5aVYfmj1RUJwbotVh8XmYdOs0aZE4jyGn01k3M6QJuwieAHrrSXu3bZvqo2R83ITgKmgRR
x4JM/wcm/gdtCaMIPmcKDmbEpfMOfc/nlBSZajn1HGON6wltNs6BhTI+Z5lBWro7JB/zLfttghjk
8RLr1nUP6t6yInR4OzVpWkxGWih/sJ78XbPNZOMtW6sb0ifKXV6V/rYaH/dj+ftb9pIkK8z9ACHU
gztHWesPqQXGjNt2w4cEo+lcYIjwGeyOe4CAoFk8kyrR7yBtmgVn6YjUskGS580KH8lFRZevYNfs
XA5Y6bLebDh6+qDizmb6YotpqQdJYgcZNqqNRlzfUifYATFkbE7m1o+9DLrpVF8/SNoE9vuTBRqr
6n4mEpphTTKHBvCyNHNMVoy/QuvqaTDbcctvs/cXukF12UlfQDfYIFYn+56AtOjZGyw3VStet9oA
EMRxaDZbiS5LUhi9hxvLkTwYwA84o6/EkEjxdGy4vlZwTcpUbbFKdNM8rsJYGYaI7lOW0RX7qU8E
Q/sKqwXVGY1bg9ltAGJqTUu1hbi5yy/apKSWHZfhAov23DHTFIYdD0yEDzf9SEvehO6ozYzsx/dz
Vvk6EAhuxsVE/7tBJbtMGlnIF/LS/hvd8ZJnqG7BsF5ZGRe2ouk5D07gbFyFuYhsxcM61p2Y8gih
bHSQNWabkWVVwqQKtGxBntPSfTLo/R5poqobw2+QWnnVIrZhgL1pvNu8GfMtr62JHTvygcN5b+Dg
dPcbwhzeTG4SBM2x8Sqhs5gGwwlyrZfalp7F8YnjiJiBxrJ3ESwx8kG4pDQJbEEIcIaynIGRjnme
awjfnWa5qgJg+FlYgKUHRpQyllQpoAqm1S2MLowICi/Cd2D/bErDbeN/7p5ewTmLUOi87M/G8XVS
FX8n7sFZlweyfzwYUFHYDBY4EFjhlCbw4QAmGsX2TkhsBvgmBRe3AVBbJFF/3tGQ3x1yFO8xXuC9
s+2Bj5+HfCzfVCyhTw+Akwdt4dDJ5MPYusmMzd8RXMxp5hDpY0s3urfKQBo28HQVy4EHVo+/mMb6
khYPUg5TzoRUo9ssvYRu+uDGA4jy6PZS1ZQuYVbwD15ajgtwBm5UBmqnbbPJMw4P63Aivh7M1F46
3BUYM7CrLFrK7PiYdgTYm+fHsUHsp9T+qPP5hO8GnG2OfH1AU8UG9aIXNfCmDx58vdWHZIdGzdL1
5x35qGIvmjclDcTlf7GFcYL3TqYhAE3jYqXkk9/WCNH8/ivwepnek3Vwl+v+SA68cFkH2dcYbn3n
njtPzHD++3lJkP+Lt7ufcmur2Cix0i6gjOaywJXcV5ZeMb51QHPC8Nq0FwuIVxdZWYlhlb2B3XP9
I8N55sSD9QRgAXoLNkPouOYldKdkYOFIQNoh2Cl30piwo+I6fgRBldeo6fkO33fAlwpOPMjX/n32
81ZbzhJA0pq0SAFthoiLVbTpZe4QBU0DGMJEV4H4f+9Oli/g8lGUnpi1zkJWkXztJ0Z0N3+kskJx
kpklrpN7H32SHR11N9+rXxWAOhR8WXoc2Sdflo4mGQTMODGj7rf3hNkGpuWrs7P+XD7m5rSCjvRZ
5fyE2WVacrqq3UxSyaxV3CE691od8USDlrmae5SwXGSQTZoqpLbBMv8kNY7TuoPJoPRczThSIqAy
l9LnUxnMhYXUbROy+6vCyIdlLJgdg4r6MGuwzAuaAYKKbvK4wcjiny82LsYWCi/Ph9lHqpbQLBSq
5wLdksJOufUKNdKN+zagx+2YpiGpPrr3dCbA6sZKqoZOBNLWJTi1ETGp+jEtZUtuM/Zmh/3/7J1E
3XZ9I5AEfrhoKNxP/CyJ0BGgxeT7F6U9oJyEnM7j5hTX0f+HYF/7FzwXt4lBnBpgo5dnF2dat54b
U5S0sLVcz8uuflnxzJh4PdyBing2WopS8NZXS/tznMeCrUL0/GWp+AxEBNFNVsX8NNGkFoF6maVA
uKsCSyyHy0aOtUM9xCRbx0VGy2vFTEtV9UTezBYrL8twNRMNkD2rg2DUm/sokeSehtFcD4zETrNR
27M6+rWzjW+hYp7ITEcCdYu+Z5hR4noB0n58mXSfh385ByJor68N1N6zKkGCRHLxNyjqG2bpHZVh
GqyrjjzF9l4wAZ9FL1Zhuiv7c07tQbSidIw85AKC//tfTc73ju4+7XrC4fK6srSYXW2wGBTjZE+3
bbjhWDsDL1PQEtsyh5eqsfe6r6+qoH0bdufxgd/zM/eLED/FIEmdVkz6y4QN3ApyorRwN1JBUoLb
mk/0RQo86tlU6i+1HyFX1KQr2TgApWAv0UQPiGYasiIgi1MlhRC/hJQ9Ovb9/GUWN+aNFjRnIFGP
mw+DExcCJHMmoG2uarv+QoDbUU+yJ1i3UGmnVvaNatLeX54e6nn3twNH4FYX4sya4Lbp09Cp1vJ4
BvD97N8zfODimBYAZ7P2gzA4kM67EtHi7v6kDHDPLdKCX50NGZYnHwtMLwL+GDNSBdM4Mx9IQQD6
wpeh1f9c7z+FgarfIzoSL00UZ9HR/PBBgQE2ffow3SWstICppuGew7yDuRhG08sgVtjycL7R9n9Z
y4XL4lxmNkUPBb4KBDMQOplnooiuEip8oPklaNYkgywJ6w0HiuaViu198xRGo2urQnbmMWNjvM0E
NI2xFkhzfwZ3XlLIf6yn1G+xoweWkZTnxxZG3/SUVpSOJI/BZEmUWA0gpqOwf8vfiD2onCkDAItZ
ZrLd1MktznYjir0wOqnFjyPP51PcRXtrJbFDbzqL5y/SJuylac5ld7hnPtW+SRY1RiiO4FU2AJtK
mX8YnSMVYAxHaPF6jd/tX/RNnX60/hKLUlgRcV5zLiCwvWZWQ0liaXHxxX3cynlkxc1Ao5FvXYtA
h/nzqIl7MfyDFFZFC0cRLJ9OweqchMCcLQky2VBfmAIVN7N0+RafzdSqJgRiVE6enVZIfmaFpbAp
ENHeeZBKmaQ7QoLFgO92ntwnZWRWlFPP20nfTYlefehM2SJBENBL6zm0N/CZWwgR0VYkqZPNPV/L
aXqN0gdoEdUjhFttJy9nABf8/0gr7MLpBAtrTWrYPPSSdzeN6LAukTjNfxMn8pfotNan9tVClT6d
IqXrfJMYeDRgmHzt8Kasl+fWJZGsdrlwDLEKAV11g9/AWBdi8jhRtr/M1oO6iwN8lk2F9JrnceEx
6U5/CbDJP7JR0QDK+tGIEbjZOEKyRECFtgl5nfrw89CBQ9nMrYTfteAAlJL5yrT0SiQTAs3n3eOV
wIWx1jpg9vEd1Yff6qPAz1zMuXV3Z4by2/sbzWn/3NJbkJkU54RCL/zjrtfFuou6Ab7HX9Ztqjl3
fdpkb/RE2S58N6St7UU00SUt4/rMLdVhgd3s/ycE+WIGd50ptAKlcWFMrmYGyjVdHfLR8qzJG2W0
VZQWRipW1W/9CejMj0QoCG6uEhCGMNz/nxvrkTCln5gUUuctRCg0l3meugPjfKbCD96cdj7MsWvB
4yYQzAVJP7sAzB5ZsERHARZbn/QivU1MaSey5iWuEE6J9BK47vpbXs7Za1QnNsd3F8IJITFIFoE/
nV3082SsS70mMoG71twGuy7xNsAjyg24mNPzWuholSrj7/u1O7gEfQ6vNxi3J+FT+BFwSE93Hy4y
yt2axKp/zhzVry4g4ngYHAVpTnNxC5aENNBxhNbgm9ahfRBRHIRZh4OB0hjYnOXc63D1I/YG9in/
vZsTji3bw50uR1kOC+tEzRgrNEQlg1aFZJx/pEY5N5EaLPOfc5R+XoaxLwwSLpMpQOFHwb5DytD2
B4JkC9LvbSHxkPLCqblwpQWhZdUMGY1M5325vx0kI3+5yiXiyH7s08oMspZkMVuUxCLxHDtgAmeO
7LyU7vVCr2rQV5JWFz2uD+98cC5ax1S5lnWTzCu107QrNGk7dNbi1U+gogqTxXA/dhe7sD7WvGK+
JWieey48aF+QwDT0/cl2amJKHuOQasTWQUDRlgLuA5zKferiIfdDMjUZ7d75YCUeAxZw2HygSv9J
xZQBylJ5rNC7nf6X/r5xLBcnFsCGeFfpW4J1uNudgVeBXe7UElQxiEm7mwOVQ7G/2pwOnhkzF+EW
A6MSq/+DwR4E7WuiTDsVuZwVvj13c8Go1fvdLiZhyJ3J0gn7ldeVdFO+aXBXl89lcLeVonSWZmzl
AJidnzATzLAx537iOqCP2fIHKDqKRXDtQPhRkbyl/W32thBEL4/TUlGhVQN+iOsoV9rruxNH06hY
y12p91NjEWCo5RRMg/GK15RF4mCsNjdQrkdy1sQUA4s38/dIdO6ETggdbXdRnp6bmtyIKvscm5WV
TWMvBs2H2VgsJUvpLLJWhWU2q/LCdARMlD2rcYPHaKLZWT7VAr50MhNItMPvmxCrzt+ugOs9qbWT
4tXRoldzlJF8ylxGAx43QEWAxcQOdLMSk31QZCuqudzDW3iTyaRTWIHb6NBXN8/FLbkqynP1U7Li
YRLpUG5NIz+78L4XvFU0jrWTkUAqBr/UQEUu15jgXvl2hxA6J0PH1sa2TwEEBWTcBdgXewyKIYbc
zryEal3GSvvpj5ztRhqcgL2jtc0SkFvTLtu6Oi04VUF47I5Yg8aMer/rP8n6f9jU0ztHy71d4tT2
EycqsPi4tnRm8mFaCBfRuWU+XqMEMSaFB//IDq48CaMMSyggoSiH9aJq/Jb7WNHs/u52v4r2+MSA
ADHMXp2kqyZNowUstC01z6rzHQeth2jFc1IiNkyYB9Nc3/3/XkMo+FhYj0iKicIcKr7YR02lFbvz
0ShgCIB10ycsOUvIpVm/NokEgsnAti2+wb42FOcgK2xpQA+xaLY9b4XgWzkOxCRr44u3MAfC8NBS
h8WpHXn0qzV+28DSir8QGbPcA6Gg0kDvcr/r2xCQyES3iOh9GFW72hUj6RMjDGy/d5mFdw9ubCTT
l2ke0FWrDHhc1N+EHtmcDtF9/l2PVWbtC8EjGJtjAO2jK5xq4H8qJU474pDLk5d4h1NnE0brZICP
vuhdU2IgVMt9p6e/ozWbJ3LpKTqZ0CDLy2hZN2eWBnc2+wcYvMWcUrRTfVvzuIupjCUVclHcqbfa
6f8mshjRT3N359nAsqYdfzb3s9Ef2scN6CB/IY7doG/LbLhLRKNiKhDrtWv5eRhsKRUVflbmYs2P
Pi0h6XVdnGqRsxq3djPU/izFXLL295F/CGwLIHRfHlfMQmc3S7UFzSqLX88n6Kz9CgPE2y0EO6ZB
+jx62i+AqUcmcsTYpYAMrx17VdTpgESxFO/tqnRTdrwoeOxI2Tio7lwrjaomguAP7pzGpoM3i/KQ
10tz8Lfkx+O6tmXaMZ+f9xql6o3tYVa3TgR7NSPlRg/0TJSzI5TdkUE891tE8iBGaR9H9tq1Imma
EX0THnTC5usRHbH3h2Bolf+OU8Nz7+6HGLKwphBe7jmxKd6cDgzefX0XMeRz4i/nJ//Qev+C0iSD
FYNpVk2Rc9Pkf9cofnyMaRIjNGJhK2Fm58tsFQD9KgLvtZf7vTM7v29N4KBaqbfbUJMm5MBvcLrG
fDZxX4ShVyoViUiWhi1UebJrf9m9WlNMG7zYdhFQOcLV6NiT8Nobm51NOQIdIpeuBfJP7ZNC1ZGm
wXbDfk5S6MDutJvfuQO1yMdkWjPA8kw/ZPisIgpAsiKli/PN2RHpZ3TYhFEaSl/GIqMRsWRZIHRu
KRWvX7CWwavHPztN+phkXhgmbqYIE3+kuACzJH8SVIDXagbKPi9gaeX8/W/yRuZuy8aDECs3e1H5
k8K6MPlp0gTePk9Bspr88+g3sQ6PMR1GGRFdvJWiu0SjFD1FkFPJvH0o84WfRZ1LMPsKdMj1C6AC
lxuqPV5GauktegmVXGdHuW39Kocih23dG81zNWOE4g8s0AB+khkXEBNZUsOWdx+1sTQqEkb46n1g
SKJ4H7cM94+S2TLn1P6Lm6r+AxlP67ihiJO3Ghk7O+x8hV/dyooi6VJ1IN2eqtVhCZDE4A16b9U3
abZUXAFLem1+rRP+TCI7BNpcI3icN2BML+onlY+CA2JmqjqXsU6iYAvAvgxizZBqe316nNAFCtg3
29XSk4C6hQBRc8s+vj3VAWcFUAK7dEYA81jDgJylJOJXAi87PX4Q1/+WnANXapawqS8S/J00ciHX
QonSm0aula24W3YL55s6K7Nzlmns8PUT04yfsCB6SDWE6BdeVzYJJIrsYdceHe/27CtdhF5YLVjh
5tWUEhfuGC7UfZD7ZxnEYIr6Wx6h09Sk2GYgmVY2znAj0t7+uld7hzsZbO0QPa+b2T3US4zPwydu
GnYbJScmwF5VT/96T7d7Th2XmTxt5zzaNWQkYVlAZJKY2KY8kENKd0zXzfFNX5SB1Tf3nG/mYChK
T5wMJs+RI3uS5qAW9zoNNHBPXjorbhUCtTtOjSvmMInEgCKO+EyD0ncXcJa0vdmhil1SnsAt5Ywv
5Rw+ALaaqyFj7EN/Lil8CZ836xSrcVtXBGHWTLtnK26yiC0JiV48czA9zRZ2o+qpoURB/iRiTHXQ
xiZ8Guf0AsH410w2pZHxxg1x7/VSDVpX6uZ3wU1jqQAsyZv7llCxNA4irfd/BwYHigUIFL9xGW/k
EidqH3k2600rVEZiWBMHp2jRN0ahnn2jFHBCUwrDopHDXM78I8CzKiue7zrHsKhyi0qnqqqOB/OA
vKP9LZY7uLnmJ4WtBXl6E0DvEaRYYfGuvk3ASC3q1xdCiYBw4MgKnZ2/EQMV5DRJ1kTPGuOda8Kv
M7Q6SOE+zWKSSdngNibYM9O/W9v/hCkFRKtUJoVE7IE4/0solIj7A03CINXmVTCpruU4DVXB19qN
O3mzyxWIiQQFeqkOiX+e+3iZo5YZs9+0jSloKI6dK0+eIz3z+Rh/9yDNZF3YVFP7j9D4Upq+TkEy
2UfvbKaF1mjWFUsSMqIsbgpP50m5zxRryRNV0Zkox8OVVTi9iNv4Utywyhs2TBjh1rt3nG7odxIY
K/SDcbD7sGgFVWDKF1+npDOqSRf/Osck3X7WcARl++wSDc/iEa0WTl+Eq8QNY+ApeCSxqr7u6+1a
K+5JtNuF1qvBwpERG2gYvI4TsWu66rK8YOeEgiQJx+CZAh1n0as0mfdEcpbh3eGalMtBqHRAdg0E
STUKbjzum6UNj8uTHwtZUceIi2lskE9GvKQWOmv4U5GEqvKSQ96cAa6WwR/EyJRPSWx0lG/o4AWr
uNUuNUDn1jUXGA2iioXWiYlnCUJKaMgxWJk6diGa0xBhLQBIs1iB1mJXwnRF4g1YYXU8/2pq/t/v
1lSihbMoJ3IFYXBQi+1tErTOCprdfbHgjCR8Frj3cqCjBt5rSHfxHA8hzu3Xn+I/9Bjb7Haspzyy
3p8R/iCzhOPaT7OSMGW6cdGuKBnIA8mOOKemH4K3dGkz6EC56MEz5whksGlm9Q3/F48xtfNtP/By
6zeyUMrFfF/VvE6V/VWj+uSlO4t+HDIIDaT6Umb29yJeY8bdF9z7Ffnos+UEJ4YcE2oI7DhITbE0
TcKHnEsAJqIC7LeKh8tjST+Ib4Pmz7+2dHnsrMbqip7mlo/53eB22KLu1FVMnVk0/+/qSdn+3fa3
5lx3BbkIE9bbyLjXSWMy397VLxeQh74RmN1YykK5u6UocZ/RkvutYSA4a/2jiI4wvcu2RpFb/HP/
INe2t2g59xk2Jscu75hcfYe0aV2e4y44lKyXW0DEsYXgvDUXVeWgIhCnIbLfX9DbGfBcZvSy6MgG
1+HGLr4dk+0Sp+TV63Tzx+UyJR7fzxDkKUSrpmySyk7I4a+Gqgbvm8hU2bmRwUHp/GBoMokmBqma
Q0ou6VDqFEMX5nR/h+AnFpf/0Jp5aSxnMdLpg/Sf+OuHvK//6Qz+G+szrQ39SAna2yx0/kdCyCQd
k7RnzGJRMRshselgHxxjY6ukm+f6NILLafyQD6VaFeByzHMPyVv2CIdHnZTb+2rfvRYcrAcfxI/o
C3tOEy4iRRaEX6Kt294VQfDj/HFKHMRBLEv4K+dCZRqGcyQnWYKg2Yrk4LgK/fHhos55ieryHQHG
sTN/NcC53248xN208DmNthRfvPNeopHJIw3aLhDz0hZXZ97gyraQ7/+WKYfCpk7ppV+xELY2XkJe
cOMpGlbo4a8ZVVCypPIVRNao22XCpCx39Xa3s5bINI9wWQFzzKay6tU5HvkQbH73nCVgfKbDHcds
YfLIbBJK2CXjtA/kLuVA7pwT8teyPnpV/k9CEmeIcX7xxxtO+wKsUYOdtEcVHo7BKfp0NIMRbbSA
0HWjXhHz2qkbgQAxG2nRNssbjUmQ+B0WBIBbXuU0a4sfFiFNlNHsSGXhNvY8wZeQMhWYZBhS09UK
QfjyOMtobcC0uNRn/7RXYnvx9mWdMPn+bph7DMWP5pqiK6pBOWr8tcS0iLfD7i55U5sO/lFjinbh
GEftovl6WhNfcjY7kJdgLZxwQrQuMnhNZLZeVSAvraa4Y+F1r+lpz7ZOA7RZcX2yUaVMGklOdYkE
cxsw7icSE8TqYs2XMXaRFZQh4VDuCwS9ckj0GyDEIIyZAZBzg4iCs/Q/CF4BaBa3mz4KY8yzTGrs
hVio4VqcDzQw6bmjaK8nqi0sNjHAauWSNNVh2VtOZi0iCLs78GleD/9cHkGgUtUw1x1P4QznI45J
aOOwofXbLMDZrknaxZW6O//GKEmSywMXC8RVhwIF7n1b1KHVw2PD519+DA0P1F8+dLpMh02mWUjk
mvwnLivG6m0qkoUulJwyLv0avkiWybjijP2wKUQ3s/xaK1tVqYKInogBZzwndsyx75Nd0jN8CgLf
aKNfXN+OjdWoDjWynR4sHm/9GG/gl/xVdHPafX1dVXUVUcOAXIDQdX4UO3vwvLSPTf51MdCRTr1r
NmHODM9O+DEMJ9FVYzjFDDytrwf0N2X69GV6ctBY+dXh4BipdZ6LALIp3HfF214ZBuniBjU1SPmb
AgZqxoIjGSbuA/7i0FRRrtFGgctB2tnrR4Csa+NafQVEGCWjgaljMhft8MmCsK6mzRZBmKJdTRN+
WrgbmShiC5gWBQDt7Fu5iD7hekq5p6hpJ6ItzzD9nL8dTFKtHev87vyz3+wwAUld/Z7ImAw66KF1
XH2QFdlCLBaFJYP6H7n6Y6W8LhAp8OZGEduax02upedb190Pne52jNLA0GukEkF3F6dPI/2e8Gf/
iItcUe7Vspda4nHw3ZaX9P9tJ/kRMwynqCOdRvNrfeBT9J8rvNFJBzIeCtptrh0Bd2SEWab2OqE4
uchd3a9Dp0Cc1q2Ioj7W/a/5v/sgbP7uhgK2CJspQJ4ndse/YZb5qQ9IgGjO3Yp3Trmyk1qQtfPN
tajllbQk5Xgiwu/BtoHhHTwQNpWqXb8V1Zs/YyQLbtnvtL0dH13ugj5cOZBkKmcI0EhUkK2X5W7o
ovxp1Nh503Je65FlbxXZbyTEA4I0rhrQJbbwusGJ9SRJS1OVRAskInuj6tOyLkSgVFuG2oN/JyRR
UjLThxJkYlF6ob2kJdv8vf1scaKm90Yru65CawaS4t7jwZaxv6kZvPFfECr7AVrqn1fDPhevJKXO
+byVQqs0/+UOKGSil3ZDSublyt9o2lFadRF4JeP8r+dxsHbCzOWmwauqWR7GuQkVagPUnKmULKc6
5REtTUsS4wZBrs35W0zZNjanK+jUj6gcNNnCOa+FxmkXu37K36X9K4h/TxyAr0+vbgsAZA4tG2os
u8W4qPOmHT+XR+ITJeWQoa1U6hwGpTDK/LCrbkyI/VMkpaEa2b2gr0wk1rVFvw7cVCjV/6T2DSOG
PcTYPV3UA5IrTFa2SYBlR09xH6PiJ7tXmzHMs42oqe7LkWCV/vctDI2h9ZhA8koY6YfA9XFisFH+
SdzNwtAJaI2mHMZdV0fsHZZHbv6YM4nBXLeeuyQd4Bmsgc2kZuvItCj4i6leNe+2Ui9MdSxnvaJA
MYR8+ivNfmpVMdSIUTYhe+PzdgQucq4cuQdv9sug+kWm3Zg+GwSHlJrPKZ5f2rlGuwn8LFITJR31
Ez2KngDbfgxRXUQODY2yzow/HioTolS5L4FuUWLZn/fobTQd2KqYqVk9FOgJHVzcvsjOMRSOGlEx
PqZ2qRnk5PnyeZo2scvTUvUSW0dWWVvU7sE0LM0XMm43TMA3ij9n6yG1un/QJXRRdUeSMicD3SAQ
Ev+hzB2oaTx3FRZgW0B2APDLWy4YqFrqUV1g5vsqrXpcmHAZ0zIXgB8qslv45lp+cT2xeDAqKk0z
nlw3Oq63YB5ej4gY5zGCSsN6oiugCXpi4hEQBKDuScjj1K7iEOONyXeIaBXEhqNxMT/2+cJX+sxt
XAjrKMYYSD7HKugetpUuRWD3LCwTGdlWLgiJCh4vMaM03GUttcg8lAqi2VLuh1e8UQxWqJy3IyE/
/iLNphofilSYQTEVDYmKT+Dkm9Q8sx1EsCh/BkVFGx527xZk6rQIA10HNUXvQTDgFX7DlYwtb30Q
YxrsEraaZLQ5BdbCh85ICAjUsmPeFh2cUOT6BFtERC93vg9umiVhlPMFPGDzMqWaYCs4dDNDga5t
XdGD8hJyUxPQRGg6qf4qH+vV3bO2rlwX2p/V0uiTIUptb1rwb64Z9AUHvwsyqdyuLI1U1eXLIg9y
8aU+MFeurfpYamd2LqcsfxZhNKeKarLbKDXSrHtq9OPE2Ll99LC2QH6S4CD6cqjkcYqIRCVIeOv/
BN7QYwd5/YGiNXNsF3Z4bQ3hiHrSg7BFz1XRXoS8llTFkEEG9rDK5QzaWJTS4EgqSHQldRYjwvLv
UIpJOpWs4FJv9Jc2fqyGZQ/+r4/o8nwGdxfnJvtE4SIbYaS9grD5Pm8VDEL7Wml2KUdn3loVibyf
4PmYmJ1r+wUqj0n9mddI+c9gpynVy5I9gQ9wQYSQT1ohVKLlQNMNztebxObeWZsYioXaRonl38QN
VF3afsYzSaDi6i/WKYPRTe7KW2EFTI32K28bnrFop51ePM7KFy+VuPwp8gvVjrEJosbIuSMChjHF
e3L47NK136kt8bM3ensh111dkfc1R2Uw1eWeQkd3GxB8OJNHhDz21LV19pJ7u5NgEMQ6c1N19+tu
2dl42q0oFyQAsixyhA482gFoaxC1RAYzFhCgv0RrEpDzgUh0t3akbuKruVgXcw7p4ocgDP0FAalG
JhydMoikEwfXEr3GiHDOP0pwBeWmrTWGyo5ir3vqp4dloYnHJyJg6C75VW8jZUFxzyE1imMWd/y1
u4Tsf1ZOmSpVxjFtf8mQwHmIopj/YEeuhFPJC+QxdPXWrrC/xCVpEHX2qjQUdhh2ZsMKwMETOc3n
vww23Mua6fZNuNvZpsGWvxkq7riodnyQeM93cljPvXVXPk5JT6Ua1S2eA4ag1eihhpHDk3nPtEDV
0v13TFLhBmsa2U9rD9TKhAp4ZhJf6JzszZMG/7CFriS9hRfg0SfUUaoM62GgiZ50U9JTMHHMAhqf
/eATiy/BOzxx6mgy1dtDxiz1DZcnK5QnEMGwvd3PIejZTKQwB0bUJGmhinmlyuoDGwDfGeP5RBk3
unCMdGPW6nqKgMSdhmQCc7nnbOWIg3D1gIPsHZZidgtLQPDHrtAfaH9lV6zraPHyi7ooDV8aWQPc
HdzbUykoRLCD2XVLBNFsd1Gtr1XF0ExVAcfAOUuSpen7KSrGHaO+0OxDZAOJJV3ebGxmCRH49vdL
zglieApAKvosK+IXQAzFU6BkIlMv1V1V8VQgmekk3GkTudzNPAHat7eDmh85qaWZtb0iWbTYaUmi
K6cgRGXa57LhEYQ+22bctcW6zwj1TSLoRO7rdvJImBi3ZdgwnG7WWZCQYcV+iJ/EdtwDeRUzkAh8
X+IgboFTl8qAs9Dojm81cvsYM9ra07vR6Vev/nkxjkirsaeMBlcZZLItvNVTkpL4oB1ylbTrhUYr
XLXk5UlV9Ak3fhW6p2oeghM9ldxt1YMLmg303aaJdaBHYieTuzVSys2KMHIydIjqf2/CEZnVZejH
stxkKQFJCiiCaDpXOmuJZnP0RVqup9mobFzbv2RvSjvzlKJlJUbquz6OFDbXtWtuvc7yweuU0lux
Cu1APXcuif2qlWcOqE59CmhOb4tjnjWiVrnYOZcfELtDQ/Ia8UtXVUHBuUMOFkAZmjzGTn60LvjC
qmKx1hJN6+9TtJDiKE4RfvlTbrGZqV52FdXkyisPsOQH9jZ5bJRIEoYSwfMdow8KsUyllB0y8vjH
/NkrlNUpSKzewcp4FnV09eNXovbN3krf3Xjx2XWtp2jUcnxrvPm57dUC0aXB+ah3khKluHL+ix5M
jiNOTSnzyDY85XPxi6/aauLP1fKDT/XlAG6LteNnvF/STwBr7T3P7njcKpWt/H42gHgQMrW7h8oL
RTQ3hNz4wgI6UNKJa82i7b5fT3X+NfXAjNLbKZbgcNUhXFtIW2Ihvcl2JuGpVl4ysJK5G1bfJ9J7
68jfUMBUhwn/2IHvcbbY964Qhf01hMyuLNItIXd4Jgrd4w1v0PT0W3nWb1Sf7PQL3hP/rSxgbHpE
sM7vLfIaWzYBsbmfydG7Pzm2c3mChRMa8vrlt0SVH7TQZB094igwdhFNdPqE7GIatULau2EePn6w
WzPcXBzL5FuFVqANQ1fEUk+CLD/3dkIEmAkFcvTawjXTpLXCiZbFMgtl+k2fOihUiugGRUKZoiZ6
11mLpJaDgd0gA4fUaC1qrSwBr8WnX11yEbqkkablyPaUK9lUBOtstov7K5p8b+w+cTiKvdgpnEUR
ccBM1Yx9Www+GSgAnlgdBjR6xXIpfMDVjLKCJY4FsF7EOJ7PfPoEDN0wPKKBAvF+80tOv/Ddn2YT
JDzyr3zdXVEpbyT3IWuhrYzVnwGIDHQEvF9OSuVxmmI+LSTmLc8PyGed1kCib2xcvoqvrxuT4+71
XeWYi13vj0YCd+f3bz5TohzRhWrhXOR0ee/0ajSyhs9DP/I54P5MYMo8OzGTOUVY9do5i2he5JRu
i0Axs3sNsz/y8gLgDizhHkK12iUF7El3bdU85rWbxNo4WgIFfVAeQESll80sIAMW9634Lc8pfr8T
mySTyu0Ko2IWsx6NEx4ZTSrum+9E4rhInRixaDd0BLgtLbxWx3+jfHMreOIpXTd6VXnubUjjdhLk
tFbqXS6cWrp2oaZv8qNQy3iFqJC6091e996UW6WF2a6HuJtiotKog6Wcr91EZ45TLKa9OO9aK4On
EFxfCE5WqpBWhHduqeohmh1ahsQqrI3R6MLZ6A99Ft/dEJwTRstKV17rRA6teVMfTiqV4ScjIT1c
7+/YhrZedVKBHyliPiIgw6nxGpEjo4PyCkE8uyAk0l/+lSOMOOEm+FNdcKmweZIYWkUyfHVoVse1
IwtSG4tiDRNBsOKOQk5vQG9RlTEklSCrlL17vnd8y9Xnc8txwCkbhyKKwJNmbKDSUq3fcO5wkC3t
Gn6FvrRmrsHOLL3YhKJl7V0KwQvSKgXIkveABCmSP9QubGGScp5LebY5EKF3LO5VkcCHPNWh6KK7
USXlMUEk6J/r/kh/t37elVwWNL56jpxnj5EPGK7NrP8zJg/MArn8jtHJBqAPaPRaP7oLqCuhNcu2
5LjnOKsVLNk1amZCz+yeV05Bj7+dIDrWa89OaR4ZxoMhWeHLtUw1vyoi9eAqFlR5vSTfohs0NEKk
kQx3ychfaTob2Bj/IomccCO2ODGz7jGaoaFaklN7LOrDBavAfMjOmvDMAzsL46QQDXASutfk+0li
/RPgLkbBdHwz7O+UDwcd0859RcaPHdpRo+DEHXgeUn5rPRCPmFWp3BRNxTgs73sAB6R3Ogp+jsTB
r6P8ro9QnK1nxd/NgKPtFY1Txnyg+I6NGwNAa6DrVEPRmO1wKstwD1SGt7yyxq6ESsdsZiVb4Dkx
n5jrfOQ87RKHFgRhdf5WSwmY9byzzH1FigcNzEUxDA7qpDdLNYWK5aCs9/YJ2RiPFsmOGp7BBSu7
AB4l60bQjodYNX92fMHRGqG2mlZvwkyLnWgtdpj0SJXRyHKEuTxCRrZTK6pWocx5nd5p4385VA8p
dnUeWQT/pnEIbsSHR4mZClkv8LdrgDiB2nD8TpLWvB8emGKJLUroCKbqzGxf9JEXHBrQs7K2aWpB
rLu4R/xCkUJpeDpiGWhcJijh1neWQeT/O6ElS86scMZhla0y/zQYwPc+ZSUJf3Pbb2PVUKxseB76
Dbyj3WvYPk8eHgcRJGUcDVI2zyGvlco6GWU9MJYEMQQP9Sb3cR1MPq5nVNViaUD0OuiCzKjDUWH2
/ISLk0wH8NWtUV7uEsC7LHW2vgbBN6xIAD6LqHy+qMxe+WLLCEQeFTN5QAtUWvJh6mtD6iGNS/Ml
QuVRV7HEDGGIxtuj0avfNmHasEDUdwYoj2rya+hSAbVbRF875PAZh9+gM/AKW6SsqwdqN2FNe2z3
WdB3vRxBWRAFLDhvc0l1hGf8eZnYEyKvobYCubJiR67shN09/JQq8rxgNMfvVDZIHS7JDlmzUwOw
YJfI6epH/pgEDxilj+gGStLxsNrSO44y/jc4XPI9AnVhdstk5xGpAJg1lSpsKPvWCWw3U+pCfm03
XLuGvr4hoYkM89MQ37ceNlFWXxUuWGXOF2oCiKhmkr8FxNKlwXk5jJSvU0MhYYa/d4MO4/nN7LyZ
rlUEYsnIfbK3IRdDavknwby84X5Gg6WB5mNA8oVvq6uEzsvDFOVRRD05ppn8nwD49GxZE9kZSktX
8idvjhbLfCt3jobUkb2AlM7Emz1/wa4Z9n3lK0lc+ov/4Leoi65lcDnm4vDXfu10+3eTR6KIeNUP
Q26YF9+h7GKmOTzZpJZtpPIfDHZdhYb6gZcSlAXcLrnTHZje6EapoY2LkoKnJRYacSQpWbJ1xoeu
iFoYB/dkIM2HQC8PdUpgYh4pLx2G5kUkHuMtEbLdgObxbMvy5yOVkuYtkpH5VkzRWm1/BqiXwhZk
keT4mv54n19fIBbS/fxgDI8zCAl3pB0GxFVY1hhuFO0kQ4T0U1hND2zIiQO2QROHPYLYTKE77i+A
3ivl0oWq/AiJtxFNQLpDJ1VxzCeiGiq9ykP4xBo75qPVVvJc/oLd1gejqIQgsVUIJ7wPeM3sDwuJ
6exTEasgI414sSSJ8CidlHizGoh38ksoDFFhS+LBEzBrTA9brTb9BVmr23hcHMijjMOOvWgPe1Ll
yT5FZCSeX2lCH/Kf3Ze0R9Q7iWndEKlezO1ikfRGvVpMeoODxpwWaUvX0wTkEeRdisFbmQ1Ay4YM
GLKw7jqDDpJ3lzOy3xdi6EOXzGxSKx8RiDUkWYSMsqD5Q+p+wE4h1NyRTgXdhuPdghTMM8T1RY8o
R9YGvlTmAlrlJhK9MJi3UhE6k5g1p5KqmkuXlAY8q2rZ7LBrnDIkBLMiOZg9ZW58uMNBtkg0DqBV
JUOs4Ek2+/UDcBNXuUGJNP6GwMBFgRnLDShQRvM4yqLbFJpGOKrElvSafbo7zxwU7O2rTL8rlg5a
badD5n2qsXgGyjma8HHqWVjNXFAbPrbBQAe/uABKiarCyN6Z8+/6VLf5SL1vzSanPThGLFLKu2FD
iEtOcbA5cGu8jok55RGdY+Mnct2wwGrBfqMGxYBy+Vvc4lKjoCDABi8Ac8qjgroTRE3ar20Nbr3K
wRVjkmBfEkIKdVmF6uajO92gN/hlU2i++1KirdPrY2ywU/62NMKJtympaMa1lQAReK9lW+SH8m8U
Liso30l4IRja7nmjo+AgAIf3oKobyz4d8fsvp1gRLmNBYnyFAa1xV5ptcWqROg/3wmWbcIh3fxme
44Xdq1weAsUaxCTDv3NG/qE6wci2V4xAOqP4nDt8j26SQaPqflEPhcUdkv55NaoKE7oAxM1Q9V01
W9LGDGZ3GOMh5sifytOrqH9Lps3hfNX1WBfKvhzU+WArGefyA1Nmo852eqLmpsJ1MWVgOxm05eGi
PLlt+l3X+Lo47F/tjJocKIFnVyDlngPcDHHB/ZrKKxTIAvbNZDcX4aE56RJDm9SAxnScKHnMRyz2
ehFGgPlID1PlxA2djoY1DA/Anw+M4GFK0qXPg8KkH6j8SK+t8qDQA873O1AhLk4XdoG5nzlwbJq/
4c/LvUDnwCY89jQIHA4ol6n6o/BptBGx/QExwLY5t+Cxfq3o6Pg/uTBw9fgMf7agQ/Lvk+Gxc7iq
6qSiur2CBqn5mK8B6nElOVfYgXHH9GFm5xQwium/z/7Mq63niKuvHik7bf/78k6gAMDv2pmZaRYs
FZ8IKlYnGfE9gwbMakT7p8kEsH2UPCabuAKcbqbmw4Sbi3jTO7mVVDXuXcrZlwV8NSKoD5qXI5CV
fwMKZMWBIYdRQ1wN4YSR1JyQV0hk3a6euYgOzy/LLgf/s0+DsENlbvGhq48ZiqDBFQBTijpqTJXB
jTH8DZPAw0cLDohevKfWHSxkWoxyd3a7WTCB4MxrVdAVgoHj2Qw1aX6I2H8Yk5l4ndY/m/J35Y3t
amR1YOhNQaV4Jw5yPqTynU/ptoNfx9mT9JlqO1xYRA+n72/mrpOlREmG4R/vntFG/8Xqwd1qAXPJ
6NZvNVNYnYnSzql1f8HDyJOJXRRhcYyf0ybkvH39K+1LaZFNT/KcKdQuG8qtDuhjMBcrlo9TBwYo
LjbqO6sskS0Z7n9qnd28hcDMJOTQI14juwpZf6UZxFoWo8wpDe/TldqERwSyujHAsXqmX1GgdMIZ
oX5lreQDHDJcSX3/peFgxFqlw55XNZqbnOfGxk8au+CpEwvpnZklo7saiGpcV41KhLliVV49sVI+
YUHrVX/tSznIWNrNviHZoaJ1A+0B54T4U8E0TVJt/2wE03XKUDcJmVjwpaSZ5Xm6WxEuBxK1GaaC
a3Gdg0QhcU5F/ObCZLFAF/6mU+6egH074BB6L28nLmIQHeEFl07ESskOzxQMRMNP5+DkOMwdRd2C
uAKZ/999CijKsmszoa8WGCOEHCnrQ3XmaSC+jba0BXdQwIUke6Rz4S8fANl6PImW/11rJmM00MRT
onZjQEaOQwiYKD8V7a2ZHERrcGwXxrZoe1e2iix4jcldmVdRInbSCbpwJ/toFMFKC5LWhncXfU0D
y9IdvihzK6sDRprnkwyq39KsY+7plAsSlbxaDADe4cX+Oh9MePbXRkIWezWAjoZaAkszZ1N6jGm1
kA72ZeqPOlOpFVuS/cp8H4mBHZWNCevrqsMqh/cp12m/3HT/nJ80hOO4/ciMY0JZLyRuNp3RlI8Z
EFacqAMVpV7qS+9WPEKkQ3qY9P6jmSpp2wBIfW+/++1aX11vGbM11aqZxMhvf0Rt8hHUz2NiwBUA
+vaQbB3ylbly+SF418vCiW5OsnNfsoGnl66hlEzeqvJGbLP3FQ4og+LuNQ+HPSiJ03vs3arMQGbg
sSMXy9B6sdejddI+S3QLBRlItPp8exwQ1PkLz+L0WTvaHFoQ+kTQ+fHpo4QPyrFKfwV5lN+gOv63
1yZUNu/liuG5c5Za69ttdyp2mDsIyBDJ7eKvTv1UdOPLfDAFzQDqSQveRnLn45WzJnUyVklbUgd4
kaVH5H0R6dOhNz/i93i8Th0EF/rtIyvz1k5PeGEtEN85muOfDrqi5fuaMNpYwZNkyW1r6cEhclBK
kjokLzYOFuLPe2MdNgudtho+EI8FOVFQY9AsLz9ntwg9tj0yDgEXskCcAXwNXnnkRuEt2lADdt29
3H0doc97kBafSnk8pIap5Yxt8tW1WS7LgVHDN74GMvdz2J4nP5fGyU63yjm9ahgiH3tHs8f3vouw
FZpvONT4+W7RZ9MQb2aZ5kSGbIlx1aIOBCuYuLvsCVCdXGP9jtKU6u4s+xCAScfhSIKrgbM+0q/o
If+uh3Ew+DzKqILVOYRxMqs67Lfmk3f40OOAtvOCd8uIv0rZkj0IueUH1ZMnC2a3ehdMXVOOnJ59
ZQUNK5Kn2pDGEjgjlwYTfo2Dj9jId/2+p72xvLmVL5Cm/Y4hxIIbrHJlmvrMwgnlMu2KR1a+2ikP
2J1EyBvxat4Yg3GDS7l4EEbwLbNBNQoIcPsjoHwism6ZvUGwf5eRSia1tVle3FLhVlsd98vwY+SD
PnPGelCSdQJ1hrt/gmQJyY3UeprghD6hBeJFYE9Si+IAz3AlptVHOBsy6D9yer+y7jxh7cJXCrR6
SW9ODEphN08n0yr2SMrHrgXKznHvsCGsN/A0q40WaMwoajCQfIDwVFD3Jl+Wwcc5D5+S7XLcTEeA
i/DJugPuUvYFaOElKhOXSMmwXTLDSQJ7i8AotXab09QQeqljVySeqmYj7Z2n0HeuDPTYdtj3+NKR
r22CI9P4xx67je4B+D7qLlaVBgMowERR7d9R4uyfa57Mp537cQ2BY3PsNPedHfvzWvUcy13e6CdM
mECUF55fjFwc9lPCLJD4PiJqu5vnAx6uf5jtVw71Bi+0NLkrIJEGxdaMWRiyHDCedZtZKSb5V410
Xl+YtccYuGt8ZY2K3p9OCuMdjVAGD8/rLZO/yYIkl8s+G5Z5RvzzwNs17XQ3AKJtqjWs8SlGsyzs
cUlgHXugQO2Xf3jblBT8u8PCvpQYAqZndQdAwmDfALpcgTyNgU1Q5xk1qQ16sufZ4o5xpp3sD7HT
LeHXOfRmMbshpXXcX1oQ+OndcuRcIwXUU493HSSIsXsEwLVmfJzs8b006lbJxbDQ/0oN1XqKC1O0
N12WeEJzU+5Y3HAfy2Z/OaY/2HFY6zAJwXJs8Qe6z+5wulE3opZ02qMZVjFYpkkHZLzO8DY+U1xi
bsZE7Mvgj6YkK/UHaSECC1hRAo5OAv7G0nDk6i2AVpoDPqaEonX3MAE2PNgBAB/VQl0S1FwIIlyJ
AbyQt23NZ6f1Vg7iGHJ0LpnONUABXtUePg+sG6lNWoUt0uUe1VnynxQRa3JI4DWZoGuGMuHw+EuA
ZnikF491Zeord+GOaG5EyCrISunz+U8lph7ZMRzg0EyMdI4fsjsLf7P/MxnfWFRR8gYZFasWXeEu
5pB8Sz1dvToWEOTxgLjmhvGu6fGEaVHRi8oStFZrdmQIiywJQFD4KDNo10/r7Fi9ytGQjpKGHOP+
HurwQrlP4UCGf1iWdHQfJTSd0RT158GEm2j61YP+zpNbJlb9RrLN/ZQb0EVT303iLIUUAu937hIb
z15Lfo0IZ0oyoMrOMqF03lkqZTFivU8taoW6D/5bO8C+FrHpsiL5Bcwl+Pk1mkqrtAtHrfzJZMHf
95WOZW311s3nn0qJ3Ri68PY2DHFFymmXdpRTOSAOpm0tFTnsD1QrXv3NRl6ojo18Jy7+OI8VFb0r
wcL4k+83UxctWzpucmpTND8wWFQb8fqku33sK4NzHHkYvjHczfEDnoGulA4RO0P18wdzzHJnzHj9
jqmEMrZC8XuXm3nRFpuomOpmVcjtjmkLpLcDjCJcSrkBCtLUWFljCSsFgwE2NppZC0bdhfAaPcfT
C5QbfIbTo2Vs5fm0hw51lXQB9JkeHEyHf5uJkBrryxGmByn6Q7AfP08Ya33si1npYF6zfNDy9Vgc
BfDvGEyDwHoezt/rqhjiFI9cv1s/f6ux0l0+maMdltkx9Nx3AHbCCptReZ+L7QO+AXBg5gnNOGKy
S9iKGRk7K/AeEfO8MzLB0C638T9EE5tDtdhCcoI5KVYocpDuUtGioA5ok2Bg+TGdlCuJanjDcqBQ
PWyf2wTBzRrZjTKxi0PCrAghyDZKJCd43FlBBwfDbAI0zyywYd2H4wptcToiKjIKVTEWddlxGJ+z
hy0Euqq6fCRXG5Q+5dtVncK5GWEO5ifA6/f+A5BwCp+li3JOSVeh3cE7EWN0ClaXyPYa0+fixmTO
DPmer+p6HxokvsEfVkjKrViDWkReBa3GH5P1eOswrI0xMqiik0Z78Fjpyuszpby3jX1p0dagAR8U
Pcm7pER+x2QbcXxBrIFd0wkm1ZbBl5J95JtBppdhD3tFdDo6TNl8OsE8ySNvSQXlVoTmzmoPIPNJ
B9x/Ohwr15eAm9/nBKe0csJhYXYM5UTyyrTDphdhI5APRdn68rfdSAKmwxeLuc6Eu1rr17eOrHEv
WL5WWVE/og5ASMhp0RjscIHWIJK5m7Uqgv14kZsGlG4vYHhQsoesMCVmbTboWWCCjWgQPT2qpiJK
Y1Gqb/ByBz0lyFZJC0SFxNJb3oDivZXPsZORSvgGreOeD/nW+ot4Hxe6AtPgUdKJoEI3okK3jDtW
Qk75Wc5VmL4cITxkuqi4L3Fqh34hIrHkOvvfm+7zt0ReV7b/MT3I2yXojNAqqnn6yCD2YYgzYZAa
+pjMpbG0Ba9f+ZHiqr+45hAtKWkZ3xJfhcF+FzPRTsIegn76WduFJOtnoidCa3m6VxwRb0rji8bz
1Wbl/osYZlN/ehcHKxsicZeTVA2im5VEgJOuFP7BkJbALfwGoZ67Sv0UXE/FoJbw7yZxkdgzlCHG
jG4LjVy960olTUWvgvX7BJm2K0SjnU1zOeFoRuzeEj4xUDozMzC4nLi7dU3iBiAa8FXKtqCANcjQ
8nozB4ei+1KZjC/KL9IM62Foinnt56EpaSR5aOmEUah74HaleQPj6q8H7JZZQnZ4Gd9zkMwFm6MW
nbM6gcYTD7tYpP/A1IU4sjml3R0FJYfwznQU3skSFXjlzk2ZL4p79hwKGg9bapK9gpEaIWLXyM/h
91cveJuRjyS4HEsI0fwdg590qF2QvMX8XxEUVdZ/U4F7HZVUPf7kzsjMiYvZ2TECZAKJewKxddle
bCOfQLXzjM/CbXBZxPJBQPnvXATh7PPzRCYUX/fg4Y5sBIdyfdVaFestyFbs6q9Qb7TR54S8w1XB
a7GR1dXVPSytRsmxS28sGPNB5pywTl1n07s1pBnWx3z1z0B6aiyiehOHQWiYZh+Ym89ZiJZnbE73
6kQB/4ocfuVrS/fGEWrS6bgPb7073KL0DP/2+geXvVpqytVlslV7lHSQ82oK0sRDgykKgnUVA5/M
XOvpJ9oB0MRKdlUNnpbaOlQLifI56zUo4IfKhHgVcd76ex0uFJVX79CpYau05MQlo8Y0kW7zFjfs
mn0J5YujYVTJ9J/yVKrHYXPuaM3tHFrvFBdQzkhlCicunhUaChGzFzPsRmmilAgyyqNkaP7lHxDV
fjXnCqtRmrW+lDZW8/M3OTJwDauhJIgxyW/VlyUdqY3b0UtPYIiAIDiuBchN9IUOvjbg3OU1pLa1
5s1pNkfx6+Z6+hv4ktn/ztWhuyq+LNlwbCwpjRSVZ89VEXV+oyviwze0Youtoi3Hf3SXwEZHO/SM
AURFMauqHQt07irTO7gmSzIzo3xaL8wyiBStAaTuwT51ODuLrtwF/k7v3cLV6vsPJrB6jysC6Y5F
h0r0Uh4Lbws14hzg9bciz7ctdGDJhbgBJzWKmlpH/1K683Iv6kBQOH9sFrUgP8nP2f3WCudi2Rkh
4QyQdy4TjjUd/h3erXTxqxcXIaVyp+uyvjvDak/9Yv5QrUih6Eqg5nin9xohnh4CByeM5strz5Vo
ilVOggqb3dU4Q5uqSOVDgH1wjlWIZ9e7JpEnqzvvZCrlL+jhj9jVs1/nWdKrVuux708Vp9eY9NfQ
lCjuf1vXaHtr1xB3FCa0TF3ZSk200pomGefkFuYrnUHnJj0odc6V1MkBOzaiDlBeL6MVMQgLIw06
rYGleiAHziOdcpMmDW/XSDHWEkQ+kTp2GLYfZtQ/kTiFpF5ChQXq4+ULzFwZEECEPAqaudQ42dRp
KBvhnRq08JsG1SVi74DE7q0SCo4BV9hmUF9GuUTjcrIg9tq14QGpYgTicsplLUcS3NO7xFP6htcU
D4kaSXXtg3iwLVd24BbHZ9A+5SH895LzVCYSWEG2pT5LTJY+DPnAv1rwh/AzOK2RA4xCC1+pGGEC
L07IX6xjEnmWS4xBIrNM5J0oXp1lmocRCovP3ncqPEnMA3Vwp++/ummEgjRHPVoH4vqaNX/JHdTx
pwsOkyMWc5gkj9JY5UH86nW3fcVyT2OVXmlCmUFwLwwQLLb484A7zA2NgJW9Kpg+Rg2qU4JfmHqh
ZGdGnRch6ipuDN3glxkYDqHuJkJTks0ymQgYk1q42/QUIIuIfeNdgZ1DGXPfB+iTwpG0iX5CtND4
7QqKdGcZ9l3xyLEQ63bFqXIAPQ2o+N6KF3UIjUc6CPgvMFR1Et4s28GnJjv6JUKtyTRw1OCXfUWw
1wDfad4IsPSKUC/+i9VMyhVBnsxNvJPba6Hxeh1RB79AVXPIn+L6TtmHJh+eXbdSMLfF0d45wRvz
4HElrBoHW0aGihZ5ggDET4YRfbOMNzK+vLpH7jGBkTakxdH128kiTCbQNSw10V3sfHH0nzHnQ2y2
q5AVn54LfZLVnpDKtfE+a6op47vQB93kfoZ37lPNxVLKoh22EFvsFhWUaxCIoCwzbOXB2x1M0O1N
H+peJx34w8KXjBdh9/XqN+P27wn3qTVxS1W3hxvrck99sUFNEqDoYt/N3Dn3k0UDJcX9jF4sCcIm
+PBWM4L2yHZWw0yHHKJQBYj/cA2hEFeuqcaIO1BqewCLEQRs3mFPUe4EVtlCeYoz9sNJwt4xWxcg
wBe7oes1svvFZ6hKFm3IY8Pa6Msahz5IZwwSKr+tEf5P/QG0AqgUSb6lBEiWavmywW4VgukJtv0m
dqGAoLmi8P9cg9CYNKuOUOxOZqwbOKSGI8K5THMaNaFFCF+o7cANYvOMXDYqSnmYEPOXIeNpqPkY
QumSFP85K5RblttITeldTaY/cdDiXbQj7sQkLpPdqnXCQZOj1fXxUi3UJuZKscOVs1C7rLV//XpF
r3i/fcaT7/EgG/4wOoG9St9VVt6WKU6jr/dtR23f91sMEmK2KlZhBaaMtxo8wrDSl9iDnuqxhuX3
+6TbKdOAq2FsZJII0VxlqYf/Bpt5txNvXghp45LIEnKZfWPSxl9ig69tY7xRNgIajeS4exnl8Gvt
csiBprpNberKdjtT4fuGtDLnHnPciVfCKNEdalD64H5IDroRXOPTKehglUqXwfrKIuhAir+N41Yx
3eQ3uThUbzDWk7xhxwVgoPCAfbguWKOtZKLUjK9UBy8Ooammy2tcYvMo4mr5j0ju/KbfoQMvSWIb
xEHjDUTpU8ESrsa17j0sHcCd55Z1xAow2Kgl3Uw6melOLGd7HXf2aP+HlCvuNMNlwQYPFNBgj9bO
YuKbyVDigC99dwaB8wDj+bPkWq3yWU3kYrHh011dr7G9sIFHxgbrosO90yVAH8BdP4hD/SLN4GQO
ETN/ASBARJJAxmqnkJf6auVKuXhzd41Rnfk//OAa6EYvBDJb6AA0oN1MgsErF9XecUcnVe4ejR+y
WK0GuV0zem98wPXpxo6W74R5sjT9gaHdV77R8CvRI3q226bchH3P0rfTx8lpkfStt7VNE+g7/Wuz
KH/hhgSpfgrqD6H6pQSaHYvBXAbVHue5+WWFJwMgkdidLhKPSmMJAQ+RH4/8az6WcbXit/BZHQj+
orztaQ2+EUgAyBs6+ZcA5YkfXHpZjVqpfdE0DzEz1NYCvMlTjK9LSrH/ydC4zRTIrYGKQw2fscxB
6omuSYf+/5ovdr95h4GDvuAbsSbFHh+JC2Z9KdpQW4V36xoSEJKrtiD/1BrJjRY0/gsKCi8824/G
4hmqTUG6KeqYTHcYsr2h0WSL7Nv1IKwUay/oZdWF0PzGe6GmW1NGNJpzS++DD58OPnp52lHWRywW
q88EsQEaz4aHhGpF6uebllOFmzU6LwRbkXeO3t+LNHpZE0X5MvMbUftdKMLC6sNTLVf2fyiwiw+0
vF99NqfVPCFqAPMEW2XQJWykCPvubZqfsYI2WgvIvoEyRAANw4KzLtuhKI0xv32wAJZA7T5jKd8K
uvt2qdSrt/BDkvYZ3yi6xBdEGSPkCvc/b69/PFPVmlcwCj5OSOod69tiqtb4jWNmPV2Ky66nCJ8q
/eS7DECALlWIivJkO3TziIOJAvHDBrrUF4BZmCReu6smtBfjYqD9gXPH/PObZkgflBdFTJvfECkp
DsiNuH0mNMhl1Zway4lRIT0O5x4cczwpkoTBd7lgYjqW3YfsrRPfcekJ4oK6hZ+43IkiF/cM/Bmd
SmGNDofdp/dJOGFD6iyMXzCUqO70/LaOr5MZypAB83gCGmHLf78v6cMzxQiZPASczbiE+SXSlBrE
VlWCmb9BcqvHG6/0jWgnyJY6c6ocgJi8CxngSiJ4RGNgO9UikYLXmJA2DJFA7cG/w5yCXLXANqI5
Gqd9GieJlUe1/8uCrqzRW7mjfZxfwxBSb/Bf+3lV+HigqgineCHm2kVy0/iC05zw6MbshSaJCsuT
3/rnHZGKe4+Ca7f/MtGmf3BlYNkgaIqz7MmrQvNhVCZD3tNH59w4y91Log6fAvknH6wt5Y+/u+n7
+EEd0awg07m5rHw/AzH3eybdmobxSkwkipgsHNahI0mljnU84i9hRCqzYpX0kD6vX4tWUaP5JcJD
QsK/KcafUszPyJiDtV+mia5iATBZQ89p9PKY4dUtfj8H839FfwvkzvbrwdvO7EXqc1IWo5boBTTN
ZmDETCN+1tCP2HyWdIi6F9uLL9sA6ZPBUE95y9rJxLNFNBZayeN/U1/9ZAqj/UCB3J7BxDWslmzD
rpbf+ta8MkjUviC5NXuoGYD3CqDkvfRt0Lez+NtbbW1BNipOVw4dH6HQU0sZdwY4TpZpol1mcO5K
O7EFaahiZdWNECunzXyky0do0GsIOEd9fz6QuKTJVVOSgnsq2WvBCFVf7crVT9AUVu2TXNJFhO8j
m8QP+PjuYK5uaHBgljS2kIeJ92fanFrPAKDo35Cg82z4Rj+KYtaAd7EMQjEt8uv78OLNwAln9GLw
PU+gpiPPWo0S7kgKPm4XlYZo2Xd1nmYnxklsLH68wwRXZKCxMVE3c9eoVXkc4hNE/FwQl2/JX5Ue
neEXdbFxouFaNDyBCOmGeRFdHGBFiMvz9NdVYk9cDTwUu0pphB6Plhhc1ZBUe1mOj0TEJpMzR4p2
l7DA+f5BgPoQ9/nBcDJAFRdaiYwIWT18fDnMGbj6A3VP/5pdzDLgLYOyWI5K881yB58gwHMgMbyg
rVN0AGf7VhfJiO1c3y69gfjARF5m40unXCnV0BkcEOZvyuFdO9xp408nbM4B3tsvS91JQD62niaI
+AyVWWgEhxR1YamLwvRqAI70aLjforf6CncbmRPhZ3Xsh3hznTnvolIj4olN1/RbfyyjX0dAH8JU
tfq8bOnKjp1jx+H4r0kqkaPuRg73nO3s84GUPJk4ZGngp/JFpHFoYZrFMoSX48QtloNwNqxv3QAn
TyJiZaDA7bV7gTPZj9diCm2XY+aDlLXh7B0mHyEB77Nwti6TIGJai2/0lyqb2zmcNxYtNSgyhBL/
4+IArBxSv3P6zjkgTkrIDwsGeRy5XQEBBjZx1p/KgjZir9MGveEkjrRC0COg6L4QBMojglzYggTF
PPTrHklqPheHQulhnkvWPeCdqlcaq+uU1dvJw8exAaYGGlsJds5G3ZVcFUztodLoyBhdZQg6sBNI
2QuGFCMfIpnEBpu0rKwOszHWW4MTiEl34VR+lWuzyVb/eHMzzqKhOIHLEp8LEr10qcY31s4gYl9S
ow9wNVeLUV+3dOdTA9Rsb+jSrnMHElZDeAYLNlj8FE3C2crqvN+HrEPOEoye55+jiwOyWtixeQFt
v1k0qSilQ8SR/QKOvLGwkvoTZrV+07zAWaooNA5xAtnCsUe7pRI6RfqcGgiENnt5isxqCbLwVEdA
/aM54EitgHa7VACWVyhxWSrEUFQUHbyMzy9gJN8cfK+/fHPDyh1YpqycRli7/h2mosz2WWoC2jMy
V7R7rIF0IhMyvrDmoyute4t12X0EsLnhH178u482Z3nTHf8zxwbQWVnyhxYbAkLbyuZWbkJFiVJc
aHFiGV4q7NE2y1ged0HOm1z6WPQoExH/BjkCIqgD2pY+g5sglgJqr35gk5z7DUV4oRIaSXOgiEuw
SUsgN0dXzEY/9eVfzlDjhWh8NBQyDpIB+4/hxQSsZh2rrrKN1Xea7lCVvvayyRDaTmYkdynol6T0
hiP8iAYv0LCfLTaGLgS+7dHkyAwqazSsuJ2MFXKDYIJ/qyDUnk5C9FZkDQLRXmmLRWL9+hn2YB7q
4vUCbv/14yJBAAikA14OhY/ufDi5S6nji2Pq/vabIPChgWy1Lkj845KkTooS0bONVwAA/AtPgyu+
oydWgzASeNDy/y/79gfg0IkeWZTBl9IyAn61vdAGj/BxTfSimKNcxufUhiWmEScYkyYOpEOE9/NX
9AcXR+b9icRHeRWp4PxLOjOB0pB/T/VN6JUPGlV2cqT4Zz0s3+uXIHmwsdRWNHhNgWsyCN+B1+sg
XkW2i+n5A0v3cDqKFBeTamrpDXkrHDG2HJBNyfDbnc6w+iS0z+ny611LhiAYIDEiUa1GVYLW/LTd
SSLs0PFM7ljrG+9S249Ca8i0TwKX/wx8vjY/ZhxzsPmd2mx8Uesd9LFM27PpB+oKBP5ENhl6wFKw
xWwc3SyRdX2c4Osk45NGRc+g2w5R+Mcwwg7xZ3vdaRbG3pnTQdnkEkbhpFO6e1AaZ3Kax00mZJJb
BctAOMza8cCQjYpViGGzW9L1Zp71it+B2rnAr58azlYSroG+GUNoMVyrPhiECmZmFV8IJcPTDtlj
nweK9r79wMNKPWK3pP+cxJUHF9/U19uv0Cl4cvjEdLM5Sa9AzauEzVVKkONr5GvCMoHUZl2CkZYD
hAQd8UTS6glFbVFU4luOMpjJ28Q+uZtqaf0wXW5RGJ1+zFaHCSL7LeIpjoR71J+UZ/y6P7pwapGo
/BMiTi/QALN/Yv17QIuruNoiC5cmULH0netICTh1Lh1vO1HsR4irkV2jEbpUAp975zqGTWE1tkCa
hnRH3jwoljdIGerkMaYwZCNuKygYclqcQY/7ExYQeLZKy0ubdL/GrAaqIYtsrE7QXSzk57nrYRj4
LIpNMJX8BGu3R6qeXVSzagQRFUyz6ZRO0ju2drh7VWgZkNjhGh5vCuIveu07P9B2Uadq51OjcFut
FSyP3gBSFI4R15cMPeUZ4k2P7iJJ2fGAmQY5ZgqRIa/NZ55cfEAaI9CetJVLoaXMVqzlGqHFY6PC
yjn6G+ZK+xyJLrgtQANiIHGXfxIRNuTgAyaP7m0wHe2Iewd+cyfdB+yy5EYYW4oT2sc0EbnmGAAn
1ZyR9rlzflDEuvz5pjFNpDS8fxMTspLAz8l9MY70zPWb7KFAw8kOapE5NpMaA7TiWehHiiEssQGM
1YXzX4sQZw3B3pjKm30RftZ5nvEUc8kN5dZu7JPWpXrQvgC7w0lBNNF0L43v1M14ty85H5wZprwH
+nxLJz+f2P1V1YmjOL+4S4PFbzcWzQ9JuUeTsrd6cB48b3Mpn5HLIEK9R1aRVbP1GHD6jePFmAEw
oTsAC7GaFhKvwpYeMWcYFUNZWGankZj3/Arznd8f5K2UVehF4JMDAuQeNc9U30NeWHnjpEI5KgK9
098ScFI6JsNgAqMbEHT0ZEGce/BP5aJnNGPi5LvTgi6U8jptdkaMBlGk+94mSWx9SdBuEWGampQ9
LCIW3KJo/mLAebcNOUjMNyN49aIEPslleoAp0fX+0n7UkvR/oIxZTNIPKBHPg2160OFsu4UC8Tev
X6RsGYTLRq/JxxjJ7JGyKPxNDc54mvU7DLGSMkTBmtSk+NjGXoNhe+38f/9MjWaSTdAuHV7n/1SX
sSyyacFbIA88algbqFpLMq/TJqyeH3mNPNXhUxQb2UfK5+k8fgnmpaLmKNn9wimcaffoDZtyMr/G
6sRoNcK0adT/jrS5LY7TNhONU9LABanQW/ud0ctxmLBdSac8I/SlpO9XqqsF2DHIVRZworoc6FB1
4zEgPax2QMZQ+vV3xU89Nd5vg/w/wudJ/ZGVRlwCfgHyMgfKPU7AGMZAd6YLsFut07OGQzv8yW5Z
1ikUsxhogtbY1uCOFGiElz7WywyJ4YtSaZfEdiokKvMP1cz4loB2FUsCL+36fyGyxlP3agJilUMX
DUJ1cRLP0oH4NF36284Ycc/7HJZ5OE2D0CvOMG2mPM2Yiz8b3kOL14XYGGI5UDFegyIIzw03ClOP
9sK2CF3xwNVRwLyvvtY2KEEupPeiyrvmHwcbvgbppRY66vJOYGXfgUqh4NB46+dzu78+LVm5NTTS
83CGnSSIj68l542ax924KB0pldcN7DJ930rzmviPWCxi9/O6aCu1ZeGp7yCQAcJSdG3hQD4zshij
nwsXsMlaD5v4x+TH5+ICXlw6Gj4OhbD5mRZWGpaXfxoHAsdnQbGR65Wd2DvGAEzuOHUP5qo5KtVh
TCDRNwjiClKekK9tyn3bGzJYJ+z/nJmC4Hul4LuSbWN7rLgbKOFSXIlCuzHkMONakM4PjHuT3GlV
Vf+SjHfPaNwmzhiCyn5zBT6u8WtiLj7UDz1YhkCYN7O7Pg1mTqjwcPgAMHONTas3lRtV/2k51+7M
7/E9HehdSBvuO11/Nk4sZPJ2QnNYKhCp351fl8Tz/5dR1vTjsBTc5hnvPQJwNrNGylrZjM+WfX8P
ZVmvOdAjrBWzvInA+BzsWupsfIctFAxNUn/QdNsSaXRTqe5qRTx4O1SR2pikP8pdVkgGLZhxMFNc
q3rZTxBUy1wVvzgJkHt5g6pOSAQrEbR9Ziab1GleTYtLpt4YOo62sYMA33d0q/AkzkcmJzeTw37M
/r/8Oi9GPx7d8rrZNVqiGC74wigN7AT15YD/hwGc0iZlA/eJKEW4ysvVV01kFr6IxKnzF+4Z3TNo
mVsEedyisUA25ophF6Xw5YPf9nrqQbGomf+ALSTSxRvItponHNnDhaBVrmQnwJs1WkISF9/CPqIh
U8tdZ3+CNXpKmdtjH3iOHwNXGrm2RpbMexE6kKmEkIy81RMp25kZnYvsL7sBkshid16LG66WuVhE
G9Vz9EsaJ3A7GOpaHd51KzcPfKcBEt6io+dO/rKK/R60fm7Qlbh3XoOCIlhCK1QliUJ5joce9dDb
6Hgfdd03gM0YvQndgciI/A1nWVDhQG5VmPIwA9WHGlMVwH/e+48jTUoT2D8/y3EXnqlMmGi59oQq
sk3kQxBw+fvRhXoJ7+KitIuTfm34XrDG671tLQ8WT4VHuzlZyJsNk+TvYmXZ2fH2l+28yGFvAyCV
p3lgwhbEsmoKjsKLmpIVyw8YBH/CYl0b/YOBFAAbzSyLQ5I8v0zfwTYwkpnMRpwOey2x8J54FbIN
AK5LNgouGOull49NCK9CJqvlFFwb/rlavlB3LZ9wOaZMViuT87E5XPVuC4qrl4jjppF/4ZdZVaTv
GxNzg8TDcrStUNcmGI/2o1wWjP7skB9VwXn9apwzGbH+7NS0Z8fblmOCywtFuGbkt8AIwiQpq3uL
ic+G0c977l6QK/8v6l06Xo0ugTpuAHwEhnWzJEgwiYSAlrXaP2JZZZCfRUcgYuqLv/W5s1TXqFxG
Z45Nfx5yBd5eKZyYTwMJgbQ/U+eJ6kNmzprGiZUKZR6SYV+R10R6eZ5HI46PBVkZhC0i6NHvAGHY
yR50eYV8iw0n+vRt/+Cevn7BO2x5FvVmIuerEvOpcKpgMCYtT/tgq1k7qSf/n+FoJY9Hu5hRJMHf
1CbhYyJgM2N4c2CVPliKvI6HL5Qv8QBQnKHvtLz+6P8JF6LCbnVl8pe5dXCyszleGAh6dL7xgBpI
EZ40U0erhcDiwzN2OHEED8RtcyP2MaPOLJJbewFcSAI/b3R8LimsAhXBjpd6VZQH0cC7MQitvYED
vYABH62YObQ+7TgxFIfGBl4EuNplzn8fg80UnlRb59N74bu8yV3sUTGm5+cGmKsCji/DQqo+EPeG
RCbZB0DbeNKO+SDj4XeeLrnHUa6caL3ueK08t4tmwg6fZVdv9PWN1/DBSoZkw45vbJjjj98ggX8t
XQB/qH8JnSIFwdeT0fJEIxOOowo10UicKzDEaeAdrDV7ksJLAAbmvcq+Il9tDtPG02VFlsIBpZvU
Aa2NW7dilmDeIdWCy2Bz33oinPRewUg9i2OZTN5s0zBIHRo9j+mcHONvuK/WPsvD4CXNONE10lTR
9et+sMu1GD47uoViQy9rSM85+aJaG1Edsj5VlprMm//d3EDcH/duJQ964medlIs243eZF52/CZHa
UUnF0/1i4Gf4tW7eidakwhWa99uiW6gqv/zGSE2ljKJ/fWVgWFNLkTcVVfvCN07LEFOW+PmRFRzl
epUzjJoPZLdsEanjxuHZ7yIO9lS9vTKKmF8M0iVVru7X8toZD6wJMQvIjV0C1SbHcSyf1QFTD5Ig
BxTqUj5N9sZQV0pKUjobXoRx3sz2tQC5SL5Rungge1MEe7aZmw6LYFstrDr0iJtsgPADkajhkfhY
z9h0ZSGcOtniOKZ8bzGOSPkSCx7fP6+xC4A//EGONCBfW2xt5ldJeu83Gf6KEc4HKtfwqDJEZFGY
KHYBlmIIVhueWQ35KJfkus4DvzoX/0O26jN0Wyz+bfp/J/kyrnf7maiNIrfkAv2IsiRMbAExBtx7
lllf/jvA4hy1kV9r7TbDQyaPSSkLCooUB3I0UfwIukpN6pCRfepaI5HkpA91QWbDaeTHIvFmr/8k
qS6YuOlxD5+Is7G27Q+xTvYF7j4EemzahVVurTqp20ToHTAHuIkHBvMFkbysBSMF4n9v+x4fC2VC
l4oAr4frSoWHrMsfjwxrh6RGsY3KM3rO8i2XWyMUrfp1tTRhrkCdNUtkV6NjPeDlIv6QD4VNFWs1
8lcoIKApylarW3Ne0H5Xc7QU6DQQ0Du/A+xcvlm4/24tPPopWwEd4CuLUSEmczRePnWprjBVrUO7
7ld8FhzjhKWxLD5P+wwDEhQ1qPxwBHaA5kkezVCUiuTfg0FFCBZlIgE0/bRMq2eev+e2OK1rJ4Z/
KlfgnJRQqe9RiQahJi9He7UsLTDrEt6UyGhxkuXDzjwEFUOeqrHpdc6TDU8iDr0avGf68HrXBi+3
C2ggeM/eR7tM2EVhiZuPveLA71jyTTjT+t0MZi/+SGY1nOdc0D4gYx/4tvY6ayLJzsW+ke7KzuRX
9vXC7ZNCCNTEwYcX/fQd50QEz2xufYBZLIMQDCv2I8g3YvABdKexTKMmDiwAXQt30/vbq3icf+lB
o6YoA2SUMsOMuD0XUIiiXFycAJZ5BoNltDQP0jo97NlHyYCN5O6piJzcjKMf8nKzFN8OLORWNKhr
cAQfs4nrQt+XVe7BqEULRF2Ht4jfl3HhxHYCnhOPbkjI9/nClKxuq9idQocbmmS67EQfJkvMoZgl
bgDeu+rbUoFMIVCojWqfofXbaEVO7wBlOZ40b0fa/a5qy/bvj+wEBNNyM4clpod83y9GEVk/XFam
6eKwtuKLwUGEfjpmCsw2Yew4jrgcVm25a4hqt6eNCXkqlEtTjaBHpPX1GufICB1zY/lmdlSd/Lfw
70xB/uIl/C7K9sTyonQAUraJvLOUuSsJUm/ZTo8k+UmuA0K6PqDx6kXrFM6ziUCQ3YC+YdNioYNO
VVulvpYfIvCD3jjLkFlKz4SbjryqZhY+h6roTFED8foTs+v6h4OK+MRJ7E53pAdHh4wmNxZhdFKQ
V3JS4oYQ5sHXQs8XwP9q22/SLre/VE0G0UDmjplGhtCCqDdalhEwcIm91bKr6IBfvfJxGoQhbrgx
5Zz5C5I/V/odw/i9F9UgSZ/8h7oF157ZUfvedvY2oWR3a09HOVAN1IdBbsl2JAdtjnYYpfvvrNgT
HMxNDo+4sHMs1HW/zFgaHD7f2I2x3cYmK/0YboZe7HuLYbfNXy4LH1jE+dDNmJvxKVMOY1WG/C3q
Jf1qAjZCBDKmRH3/RdMQu2RZ0aB252P67pNK/4naSjPVZ6JRSzxiX0jJXpm/i9eYljgDQyzacDHE
uYgcEc/46w+nKGObyyfpK6D08/uEaP7taHTGCMcnOjgFLGrjLaOBKzGekw9GvU2cK5Y2zr5aUNMr
P4wwaVvgvzZynkSD5D7Pb2Op5I+CDGK4HrIZIOnOhXmPpHJN9Ksr/PGKo+ER+PPFOBuS4dS2jzLI
/CTWbS4EkLmFAuhT/iDMUXlf510Ebjg06g1j+oaxTWDtRepnuj0z3OrBjtPtpodyseD1Py61w4Nt
9BlqcIqFZsVSf7HfTynbYuTkqxadjMsOVZaAw3Oyr6NMDp8geYB955hYKEayxJBQoXaSD0FIcZ5g
NRCrS9S3ZfmP4MGD+HDWu2/QXTMvezzPPvk7kRFufvs7ilYdEfmP6bRxBbN4djD3Mcv8UxZr/xJg
SQ8LPviZNXvdn4z8ihEwzVtiQmPiRINzOdncszLPB3HWYmgok9HkJ+OqwU1754YSmG5A1MMGXmFX
+EJrdvs31Z5blDMin027qbUmsMVOCi5iUz285wH8FC/1pgGfEOCQrz0eKpmwEx9ZjWEdnaTTUC9L
8qZ1Im+cr+Z0AjgGgXlKp1xPX2fzXihavMIGcH2+cf5McN6HFgapszOelcK1rzuUylpK+wuk4W2S
C0Mfl2cyanCiZLP1bpM1rpxuOZ4CRHqYudw3Ri3SVzkKz6D3y/VJuPzBdDl1FoJAC079fHseQAYH
g0U+AiNmdnywXm9boCPic67qXSjvwIQ+2uQ36zWigl4Te/svOvSEhUguqh9MeDGZlh+u/nQBzZPl
g1OW/rnSxiI7dCia3Sc3Ojc4TWkRdFMjKtTHMwJTQk/g8pXebUWKyFSL6F9VsGXuHC7WRDc3Fp7n
Z8OZ4MGqxIXlObJU9HsYtxrqFaYu1TOctvXIAsapqykBminkgdLFktDd/e0n3eaRzTzi3HQZQhZd
rUyhvOWsP6wVhkZT0XCSZB4xnYb1/K9XpNfKCpzzTAidBUV0bKe9+vZPdnqPGGByrTdsut1ZiK5y
GcFWwHmihATOJljdnb7Vur/obVfYxJMLFfubvnsKJcdEP2YYmj61gFAMTMJnBcbEdALL+A5/nLF9
oj3CRwUqL502OWU5+xwOxVC8O1mPctj3nmKQhYkWb0KYNUiXbWKb+ubO5MyhEFwlKdO29cLS7h5q
wBi8USFwOMp42nWA+iCcU23oE/g8WbYI/ssWDWMYF3HFnNIXSNNs6ydksjP1n3uPld/PFxEN0H6n
DW6i1OB76+LyG3sNtONSxEGYiutGlZIMg4/odd1CPMOPFQ2L3zWWlDuvD9oNONdlGna+vCUTliwS
2d8oFM8JfUUus1ak/ooPm63CF8OH0SuIjJBxJ1bcsUIgsitS/OWIkNVAqh22yOM0CjW9CHGb/Fj+
YCFbbvyFDnozpb8IabJUdpMkGj5idWmTeMarfZwGpsNZWhuMs3hkouSfqoh5de9zAU1PoZ8Ghzf5
vnYhREExLJweeMACbjukCg/fdtXO/lnQ+5wI43YYOmSCxzjJZF8CJ0ZMNje4gyKq0A0UIfLB0lNe
b3q937vIx2RAtGTqLwOmH2k19Qb3hKHOc0MXdnUgzfg8LaZulXSZ4s4Z9MbdF9O7Xm0qsjIaH+DF
IzCE1IZp/fhRNNH4hh8bVe4nP5Dxovl8n1CXY8OJ/wcOpDHtDUx7sU6EPJF41MqnEroxqvLEqK0V
aORhQjlcrtyR+mJBnhjjkhKuOaNMw0MNPz+JW698BrWPmyVyazrmZk/H++AF5LDqQggNX8GgdDo+
JKyVl7IYz7gls3B/pgMh0agndmFn3vkyuZOSAsPWfrQoDn6/QRMAjv0cb7JR49JgYBN+PVzw7Qf4
Ne5ISG9j9bqyIv3mKD8ZWQCW/OFG6EP790IDCAdqw3mwuxK/tV2omrAnnv/hqHj/qNwcouMMsM4f
ma/3AcY6YugyYSpAzA5164aYJ29wCFudnSOX2GSyMUnxgCpSL+NscgHjMY9IubQzkQAFyqc6vUKm
WoyrKJcE41YVPTPl7YedLtbvNHRG9K35iKZVqNK13vdNCm6MH75bc9u8eosNkDkj8VeqdHDp/0Jl
o3gf8Adp8h17yM2Rpnri5FXONzqIXfiIipC7Wg/ku5ERG8rZ/l8WqUiRBYVxEOsptpiqN/2hBMGe
wZLNPepmW6Rj0kZOiP491YJ9aZ4t6NOEKcm+dE6/B9Pu8YOFCcw3KI0xwOqiACeySI3Ucii0BgDv
ck5u/0zv1tH7IhNAfUdwD6em5nKI6XfZwwU3eOVSoQduPUNYSDnz+YMZSGP0zLNebUNl5ID+qI/W
rjYfEcDT2vO3FNKLTLY8IGVPxBSeMMNIdNslaJdSolLACtbMTY4Iiq9tcwEn35KbFqgEMyrhxn15
lMcLfOkUoKZXosPOmBn5c6QIsxFahDyp/aSwmT5JZerZPqTJhjVP0SfdSlopQEYOkSgr4f/mtg6H
oq36Xh0uAsvKCiBA6lfdS7Y65XNCii5gSgbDXzd8yxAGa/3QtariQnvy4YfRsu1Id7/le5FNY/tG
qr35P0cGFeh5cEjF0QhlRnMyO5N5iCkO3nJAapsI3DVXN72ORfC+W3903LlyAFgheksodeZNOkOL
ISjHNvBWp8ltNBSrtMPD+76cRqlkNa7xDW/IKFNtrn5NnJjCdkxB6Wu90jdeWvs1UAqy2JRjize0
v7Wx6mXjz0mzHmfU38Zg0yGTIif2sn1Fj7C+fzY672B9a8thlX5a1MqCsUiaa5ylhCAYwkJmTjXA
4rfgDRZSbQ/3ONgM4jrR4tP83tUHUCpPguOPxicAjlKtNwyVhXKGwuFxdVUki7oO2w3WLiX5/Xq4
M7Xc/tAQXtL+oYdbwpMCvqvWYO217LjQJe1hTbV2yDa+YpJd8gx4jGQWZn3ZpwmQu4cjySr+037A
eO1owiureeFpASf7i9yi5gkzdqYwAIrVKN/ojm7pE1i6PWDvDNquDk2ibBgf67bJwvNQ134rfcLC
tqLYRx8pcLw7aXrEhFHZPDpMV5r1CXWi6CbSHIn+5tCdyTg+n96ooenkxPR1A6LElELnoeu8LKpk
vd8H01lhPqnbZgt8XnCbbsWQB6Q4W1n13oWGA5s63DVUQmk+hRPAilByCvPvgSuFnOxngGOjWI9P
C7HCFAk2xf34u8BKF1zJbHSmesRBlyGjauJ0xeJtDZ9fnzf54AMJR4LRd0mR7VspUCi24JmC8k/7
Pfyi7nyv+stPn5ge6ZJeImDtS155HFRiQv5wglcNaFUX/ATPh21Wa+eg+O3NPHcQ95D6CosgHxfb
eTUrbNp0y/1pSWDg1vdE9vPo/DDtFOX3D7iIA+08R1l8yREGd9VL371TS1GgxOyxugf2gl6yUqfh
YlmHayiZZx99r6f2a82sldKsATD7byiIl9eFTBQJjrtYnr/+LVnIJ8GfzNup8pg2IAkhYxJPAAPF
0pyXqQs2qvnhnc5X83Mkw9lNCF88Loi/UA/Blv80ORKRWJdaF0GCYkDEMQGa0LiKa8pghZ4GuBel
tzlmO3bitC9CANq+vf3Bco3WcyqwVQSlmWzALmPHfnw3ulQmVVNy1SFnrDjgQefTFwZJbKYpYHlS
otXrrLAFPa9lOfwA4YWuhpuw7VXTHw3eavDdy2J+jcFh8k510lAYdC1fea/T9w4EeOrBiQ85Q3ix
ksqEgw0YgqXR+/h34/NOLlgz63TxMXYsxfWesB+WS6Xb1RF2nDjSX2BwdmdmiWdgLvyp8yCDT6P4
xC+NdZlMdSu2tzWRqaT5MFIA5ubugvyNYMnm0IidcQGRAks7/pKMhC+p6HS0W21b2Sq8B/1rcOv5
sYncqhLNiJHAs8FLb62E8MubFzmqQ68fh7RitBzwHK7k91NVi5eHyqjW5cQVXck87ZQRs7gflFLY
aU7RcNE1hZfxANBXWLLQy2CrKS40RC4OUMsckBGNDsVUnDaB5Q5DMP9goj2JgY1ORxIn5lwl21zk
onNqdHRQWqNmDQP+TscmlX0hj63ZB/PrXtFBuzlV0xR67D7hfj5Cj3XfVO/dLWyrGyqu/SYKhgmq
L5NqmOCviIwKOVS3P9qo+0ENreaE19qk/CrPTqoL/001n/eyBVtDNRwMq8ZLA/x0U5psCG6MaGtA
v85nwU/Jrgx0nB5GTfGIkVRcRAaRkrnPzZekfMrLJwUBCZ88fMX0JYOk0LgYlcZoOLvJVCBbNEI1
W6NThVpHjer1EywLczpE5RUXWetuDZUYPffHczV7RQzfCq6IcHbZMsrYgLlw9l8SfngyjcE28aJz
O48ERmvU2t5TNnTXq6uJB5T3JPIc1ge2t/20NKMQI7sM02/grnF00x77r7oCu0XY8EaSCWe9rrND
iJpfOzf+gAGbXz+KCTMmKnCoDtSGYvuaLfFRSmwrZHJEWQWnNuVuF2zrAuOyf6IouiFcz52iZnof
RikpZ2YfihJTgSEDIrzeK/Tl8ETt5JVbYUEsGs/avXaeGq4MmDuBIqNjSBQFf8Zq2SN/lBv7NmqP
wCoqeFdrMLTb3tkDQXkkulkaT0etN6oTxNJYgoQv6dQ25rxQGP8ZcPkTjEz14zBvKvxqhCgEEQJW
c/4JWKYZrLk5W2KgMEb6K4hpBCATK1EwBTqrTURwiOWBLjGGZ200FIhs+sWxl0tqzVcD/4O1IdXu
15Ak4C2SNV7O6GChyN22V8fg2hteMT8DtGWRORcw2kEFhRkN21TujJ/eR4lqcHb3FxlpUyeSGlvS
Oe4Ja26eLMoWyTHWQBg6xRQ7TnoFDZydUxI7J9TFxEFj/NEnZgCrDQM/K2RdkdtUjVz6W6ryAT9o
sJsVZYYqMQXoBW+3syobr/e/Al77nvUSCsl0GJu5OpJI9yWybjEPc8wmys8FoPrubtVCluqGCw87
URywCzi1FS7HGKdFWfxyo5wDlwZm9XzKJtPPlC6WT4YG9EB5G/e93LrPGzZ6XYKBNJBIfxaRu4Bv
KUg2iv4qzABVSTU5fNU9F1pFp53hxNQRcffOAO7biA9vBpDjKTEs3iOvMNqZs5uXpYD3h7JQ4jc6
rczUvihE85VHftDCRiXNpj6BDEDF2pCf1Ro45xUaNYnpTudOE3g7cwiOMADXnoRNdAHwGzmhQ6BE
7ANzE1yjLjp3rhXetCC39IjSOwfWRO93Mvs848AwXgaFETToxUznwEAI9NRhVhWjNYRQvbU7FHwS
f4v+/O02EyJvzBvqm172cvrgMcWhUu3LpneMMILmfmgWKeekzXgsywbosp+iu37wt467G9WnyVF/
Skzsbh/f+rNMQ/K2i3eAjHar5dUpNrmu+GIKqquFrTje6D4bxRmcw75roEtnQnj8Saxiv9WA5fth
0SQLoAJXIJSeGFjUz+JaAcxDhJjGrTYeqLmNkdvD61DxqYAoa1sO6yPg5x54QGr9eZYk/5U91e5Y
x+rI8pzGVIqavZbF0+uTeMv9jNGQN+wwfyqqqlyf2Ngb3hi6U1vK/YJZmo7NiYxf7kU4KvV+19pY
KAVmzb+516tO3Rh6WsUnaFlWvs15w9qdYhAiJ3feF6/VV7YW1cKH7lkY+LqX61Zw1Shc/Lkxn+1d
LbjeMv9tnH//9GYD0rXwvPEilzGUz/2GHZsQ46li+V/kBVyZvnYuIziJfib7M2AMsL+oeSW3SvHa
dgA3gmwTvzvt4xkSyArU2Fl74n9o+ey2fHYZ6DQveQcfqii8OR/w0CeXG+MYPqYkbnhlBANb08R9
vTS9NXtEGIR4Rgtln7zHoqgqaxhYikgKq5BzVmm0SNx0uR6aTA/448L0R6NtoL2bbZOOkaqhtPeW
izNwTjwAzkwh1sfW4B1bmbP8XXFZlfaMpSBAzgrSFCm0TYqZ/dMWoCm2CG4zuM6+PRj7lWLLkAuM
ATsjXPPgt2pDeb9ozjn4Ouey/HNB7Pu4hmTUYm3A0Np5SHRzGpONnBkO0FIdqAEWLs2xylFzVSLq
rdx+iDAzU7JAf7aVCCjCEGIIxvA022RBXDxkyziQ4pHJa1L2/zC+Ie2dbR36V9JM9Apcyt5f0uzw
SmnuW5IN8N6O319nPUTIC8htc9/VSWJiXZq14rE3P6dveIQqqLXT7hpT5482AmGhnnaeO1w9bOzU
Pq8riPIYD9POeiDdTLbGsV/AKEF/6g2GHpXy6R7QwruNfANeyHID7KlbVmPzZ4+cEeJNGckPvcWy
6oRUDZRMdhK9oEnIwgQBtZRHWYcp47YTa/rupUrET1J7jNteK8+E8+luTmd48Csh8QjXDfQNYLrV
myUEylCM9JYAZuBd1Ux32/wEcD3wxZZ6dPWAvN0avAgDZ11n19M/hHNd5CBkl9npv1ZD4cjbl2Jh
KURW5Rvjapwm0yXoZ0Ehm183Y1sIUwD8AWPmtYDMLe8JdJPFs27da+3rdEG3Xdzg8Sqoyu6OXSBU
IYLN7HLpO8iHKxRFWKFQbODAJUp4sLwZBsmn57hx77Yhp4y03ZeX/oqWsTf4Iqq5Ht/5QmUmLDoX
prU4iIzEOb93sOW3KN8zXo749OkvC2qNXq3j7cPkiU7nYZ2GaWVs5dx7FGwA/ATicESVPHB0noaV
7gUIiQFW8ob7jCfQr7bA3iUjv8n6kUOJxsbbsoqAyJGxBWmB5pAdGnC31mRV6lEVavDp79EVyapc
hmPxe53qhpLcKFTRCXg4d1WfFh/Dr5rhWn0H4jMi0kmD2MSFHYcA1UxPydctgB6VUsE0bY9oGNYN
q3q4Yq8fMlZc6J7uHCivOYNfBG3o5+WCjtnU+yFQCDT9FlQyiYfF3kp39Mj1xv/W2lW7wL6cZs9E
WYHcKRL7+P3BT44uo6tOZP+LBW3oLdFCvlmTu3EW7NQyQiO4RTo/eGBKzHp6ujcVShjyUNqL0fTa
CxPBy096+Qxdmv7Id8pFrPxcsyBuAXvMDkLOyp0MAoAu2hIq1/urMy26/NJlSWlLLvEBjc+lKCNz
+b7QfpX3pRQKAI2I/wJBP0LKwOiXXqxhu5r1eeNjiP725hO+L3nEIGi+vDYlBkRdKZu25mELve0Q
whDK58gcsB0oCptd1aT4ojpoyeYgxpJAz+eG7t6x80C6Gt7+bVWnjxK4pYIHhcSV/aDgqepA/Pri
0iVmkdLjv/35K/NpBnYAOvZZLGZEel82uyp/l8iXiaT8BorcO9p3PkHMajrwVe36q3MHuGAHjmYB
hwyu89qAhwRK7/Jqn5myVI/Vr36HmKRyiPWVu0FVf459RVd+IyMGxL76QOTQ4C2WwbVbvuGaVDqa
+KcifkeI9KX4oKXgcWuF5BSkdYJjk9HstZNtjMSMkgQE2YKTh5bjkrmrLRSJRi7w09Mx6AhIc6Lk
c53+UVltdGJ4wJaGnPoqEy9YS/avFOInQDLPmRFScfP99SlXWa9nO633LnZVKJAxPnG4VI/xtfWH
MFPJd1qtsGc/fVP/WEtNUAbDisFC2xOt29+oXiVt1kyQePK2kivEBgKvwEBbfffdCB9AxqXpA4o6
gdSxE1EFDidHSgk4DZy3/ZxJnWEdB0o/uQ7V3fDiFAjlWWi8qNKcZidtfgnIkEMX7dEcIdAFVIvr
UhhgCzTHlRz4X4iYf5OBAlHmC6ort30+uORYbD5xkKjRwumKiGhgnUz+Jklj5N37ZuN2olgOEInZ
dLHSbjBf09yMYC6QWa7sU/dfkINYN7Jtg1uNnLEMFFYsmvOaNBiWZ5D9GXizlNJYihLVpiGMffwa
mRCav4jPmsk5ChfgPXy+ZwMrIQCtmnlCrVRznUKa0UgBFwfG9Fy4WRgUG+lkj51ApCAN5/Y/Fh4r
zhjJqJW1TgC9fgyTbt8ohIrpH4AXtR55VrerInO/Yt0wmaD59aC+HwiCBAQCJXl9tBI/g4NGKr9/
36KyWytpwSeUEbjeWBYeipnjp0Z5qR+VhI0Z3atj15I8JD+mDhHgqepMPK0sujiHnkOMoEbtM0UV
8UR6Gr69BDU/WdT72oiuJ5MMzxiIrnOaE2J641egRLw4uirslNcsKK6e4hDgot70+71GZf09Wi4w
Eg9vJT3LP6aVwiat6OIkLIREog2I2vhmoV/jrpn+IYqgLN7YX60cFQZeYZ6vcZ4q4KgasxsThlJE
7Z9dQeQvLtYD8Qhi11ZQOOOE0T9L87yd75VFYysZqyOu0MQMilaeibVe3z4DOdzI4yFk72h2jVJ9
aG3OlzrDMit5KE5mnx5ybX8VgZJcdMULs61hwWdsF0W6mXtlamk7RQPnVRCQeWsbsERUVZHwETht
h4I8XkpIl+uUem+v7PPjm/vXh2aAocxNDVZjJUBQDrdeVeTVr78rNpR2q7gC3PSQ6bJxjNI+M5RR
/Prq5nWNi9nkn6h+Qc0PEbWZyDgNHPQwjgBiL4iWI1va+to8UMaZr9Cbv99g0Gr2SUiq1IeLhs1r
3XmcPmR67ffBwa/y9N1SQdxxgvBeV7Gl1yBF8EAo91DqAI8ndGBhM8fEDOK6dvCXtwQOGmX6XhnE
iFZzDcc8Ujj+Djy0gapDLk1023z4NxuSP2Nq7b1K4yxVkqtU5BKIK6quKMFd9uDM/gurGGl1bbKI
V5eMMNg5jqFxJoAW0xyVKdnMBrhV3fPWJGwLe87dWhyo6vVffhhWMR1ZJMKfbIvWqUKoDU9GGhx1
Swp0ETwMthkESoannNbTOl5KbD/Qqlab1yChQMFyxtIa05VAIDUVohgTUZ7PlI9Ulx06jURuQH3i
j/VNdc9vnR70GdBUvxvKA6Ijg56x6GfJKtmhPmFeLvcO/iVcUo1+/n5pFdDYBWtHxVM4jdPejrf9
I2B+FeTcxYkH1LbjtZLDR/78tm4TrAsmQUAy0HJw4SBGX5SFNsslj1Lf1kpZGBr5pc5ySxfyvoX/
EiUQi2COM8KdaLfcS9fssT7TYotSIX/mzqyrvM50ymZZkEVAS19pcUaYbWq79pZ6pSzcEucYDXRm
UYGsB5udpxboIQuLHIb83G81uP89uxf9QeYg+1TPYeyvJwI3JWF/BZISU/fO/za1S4l6IuG7XOca
vvgMCze69B2UsMZno0nMookDDDJmz6y9ud70Ew3w/wGSBndOw9D4Q8exGfo1fa8SEJ2T+Z/+SeJ6
7GM1rImeY/RuoT0qNAU/jMyYnarmpUSMuo7E5/E/tv7DdGLwyvde4RbdRE0I3Zz9adZ3MwsYgwEl
ABIrJY1L4D1mzpCoAY4qYzAA2bCOXPNW38/UVI3uo21H4YWuPd4Mm1Xb60D1M/ciHO7J833LE+7H
7G8saYaUvF9Sq02U5P3spmz/iDFVlxeN94dfxlQhEy5aMhSjlbZYThXSTK4AP+Y6HqSIlYX3ToMq
lZ2qJ5cS0cdFDfVxpYmhHSGZgYfLiHfe2kqDYJ6ce/iDcccGquGJ8WcKPhbDqiaQ+VwNJvPbRuSs
oaewelh71wiNlDPbofyZnjU7P9Y9Y5PUUuGW45f577EF8rihWbgAzA6AaA5T89wzUPNxkaCMdFI2
ORkFJUq10PxAiLJnRNgyST7aX1/wS+DnNzZP2WVyt1Nwq+tuTUu4tENekp+rxvq2cr3aDSmK3fjh
s1fY9kxa5C9ve/yROV7QT5LYLN0bZiS24sJzwviai2cKwawcaYBOQkCeSrtrsXxpWO1hWQZBN9Nk
mY69zbkt/7H7QzWzlOEeGGsl5NjOweW4wxzEpWlQlSsq0yaNJWFzVCW/roAHEfuRzO77eQULaTui
BDdx57PN6wztlCMFixWj96xWAYCu53zXKoz//DvlF8uhwJjTzU1KGomFeAvmZ5sCa7ogokCLm+wd
14ML8sUKove70icthaFu5djKrqNyLjNPnj1DsvK97CglhxA4UeIi+faikU/UKA858Ry4CCJcc0oB
G4FttCHbygwjO6MJlw95WTaDQo6Q7SNXMAB8aM4VbLfcTxRSU90DFAXegwlKFQgDNN9IVVYyvu91
A/czX/oSuVvQUfxvZbwRAkZY8H/kJdYw7Y8ogs5ONEcM80s5z3ao/5RpYV5S0lw7EXjccUQclZp9
CAt9D1ft8n+pFt788/s7MUwf5Fk1jsI38OEkU9zwuYycieqbkKWHYELQEz8KCb+LUj26s2L9LDg/
mQnqnRMrqZeXrnsx5TPIQAni2Y3KxZTDonuYkYFNmPzSUkkb3Gtw0IzsrPZHYsNuCrhlL3Iabxy2
es2UwaOB2URIPXkbFKRGT8CoP970Kzl3UUaJcWvL9JskSQbttxCnMY7vHXwQcsH3nIIbmA/AhU5m
oqlDqEUeJYMJbshJtFp7WD9OFW3HIA5grgjin4Cb+1umFW5uh2xIgdUL11QAvT2DgeVFegzlrmhY
61rwEjj4hpZzPVOdhYZ4K2QG6RiE/oTN2Dp/5tNyexP+ruXF+vPWrEnUJIZ2OgsKzFNwuxcdktry
j5cWLoBvEOZDs7SLVBWUWwkHrYiCMd4bFI8Ax89V34bLZtbVFC4zLgQVY5MCHlXv7GxgSCbIPT7f
4YiilJAl0gJbsGrj1q4rRVaV3nrMaKYbtU3+vHa2FjvxAhsKuxa0Kjrd1MmRvsub48PEn1/6vc1v
p4lVk0E7aTYBIx3IS1jIEpSEFjr/CMzAAGtGcwmdKatlovMLBuVmCP7WcerBbW0jKFpeyNZsW9FE
LVbyDIaiDSOCXUWf4kpvFLNugZ8lSRXzjI4mHPh3lzp/UsZYNh7uWCRMNWis4hJd6Qn1LcQqBziu
mEq3FNjbZfRCwUtDJp9ZT9M3I19kaH69zvwPFgnb1Nv+l9l3A7GcL9SOMD8NepAREZxngQJrxsI8
/8VK/DDXK0oa/TMcsnD52siNDLTeAiUfkFHmxHIR9ZRyhh3olgBuKTB6H5HARnrh1Pi6/cbyC2Bu
5MozwEvZLCH9Sm00yv/E10y2Jv0evhYFybn56oG/RmTKF4Ozu6bhg7PQKxNyFPg9QgGtPTWuwhia
9WIBbbbz9AcuNrJCWwhmSf1pfwrJg3RkDYlPfIgxfI8XoVNGL7xIphqhKzvPwpnJnoCJqwAN4+5p
Np4cdmFnAhOagfQdrfHvqHWjEd+1lCgHs/NuVCqqAwNwjtcweXZhvRHlKS3Tc4zr/r4UMqcjvUm9
wNuwiAJ3OJAmJfkgRwGgkuW2OsbbRRejNgypBFRSuJFU10X55jahvwxNLRCKHzaGgx229mOQMQ9B
tgoMd5N8cgN1jmcc6LkYIbk+gvQuL//hEFiC4jHoohFKRwXQa/DHJDTzB4jbyhOgtC0ql4HkMu7Z
Ex2dQ+XkgvSqvU8ZzrAUz8o2RrU8SxPDo/aW7bMcOty0jDSTbqoFuE2I3OSb8B3yNrmxumHub1fh
RDwniVEcEENtb7LBfNIvrbUuCMqA58B7w/TzAoJOKBIVwLsGJ3eDxcG/eIV0FkkJRbn795k3sVDB
to0JMWRKx3Grkr6E4dY7RXThE6cdyVTlzcephtBEjA3F4iJBj2jIv+9Dym3lDccKzpZZckG5dHaf
QtnWlEtba84NYDW4fERKjRA5EtAyNpfkuuZhimc1s1g7WYbcnquBZu6wfXtqL1Y0Hnzif8CyVmmt
f2YH73v95X9JgoGKxQ1slFh7NSpWkiScvE/V4hUkaDEyupLzewo51wCAga/dG5Hyvz0B4V619+fD
LTfL1JOCg4qICVRPlq6R/Cay3M4CQGaP2kG8XSSEU9TGsd1cKfsds/d3h7Ano/XpkhGn//viRLeX
aAmKLXpRHMp12cjqPWCtP/AsZbjBIgPhw8Iq0n+W6hh1UmsLDR76joqfDSV/PziaPIWJMGZKAOAW
IQg07bq6rksBYbWcEvrCQmKJk7nn8CZlWVfl0q2oGaUmwbWkBp/ovTezxO3+R/IMJF4IMdxld3Rb
ly3Va3UaoYycc493Hm/H6O+xoWd10Kg9PFXtu3gyp2nFKIZXyruj5yyR/hrB2AmPuKptI0ven0Uq
8UBPZACHDnc8hvsJsF5DKsJzyRlLb1KCSw0aYO770OchwFJB3BZBNQ6KBAs+O11HBsqlcXeOqHF6
HzdBeYXhknq0ofu3x504BSQZeMCUSfrqKr9/qwOY6aATbVRPMAAaU28Z/InwNtiMY/FbBmpiQk9m
YklDy+uTqNxCuhi7dUirvKhSuj5hUIapF2tGC7qi7d5IC9PYx4pK4J0QF33eA7T/lMDf02bR83JP
teJUeVT0TtQZ8RqkumrBNjJBt5IOBKOPRP1bm5dLfOR2BtE0Acgl5ECuXQ21qsIBNaF7U0a+AVk3
n9znyiRxaR0ys0aH5w9zJutC+tdHvRNRDvDcxK+dTHPCQeCkwdf8N4XqOviNYBt4VbsK9SdidNQu
FGEFBOlsbhjaBoFVmsV9q/702Kffz/xdIF/6AxxGDOYD0hzlc0CrQ5lfdvqA8pLOuckC2ccE++kt
IRw6FLdqJ4rlsJB0sFwkJojpxdCK01pgCjahPlAPkYpDd/qR1/NnXzqs6u9JqanmHkmUSzhyHQ2E
dfe6d/8Zzap0Qo8GvFKC40h4hT+64k0Y+d/WbyO9eroFWbOz5/D0G79r+NBu5FFt+RCAOpFaiyTg
eEsrJQtA5zvbH6HlyYW+dEwGGzEGb3K0afZEHwJnbqThmw/eaLa8mUMvBo2hNykt6KsI/K3R4ymR
zI5PRU0Vp9GboY2qYnqQw9YpkmUavjsWsjEBA42RunkFGISujx8aWqAZPe6g8/7KqpOfYXwNMt5L
MZPTbnxolO1xFavIJHz4d7AsrI5+RJGwszZGyrCixNYo8odHVswA25cifC5tMz50Kw6vC87tWQD3
KU5sK2KwkQKE5fNAiTQpS+nGysENj3iC/zBO4Yho0lZfvLKP4dtDV9UWAKWiGsIMNESeVTadlUay
TBfU+pWVABYMlaXNtv5H7+TjERQGA+s/+lZThwGJoSnGT39UlWzh22DokCMvClAz7k8AhZ5fea0a
FUhcwQ9TTSEHQ94WazE2zVtpAeX42jX1ho/0DR0OR/udPK00LVx7UdloCmU8MkVAxi/Lym9s21V7
0WarApmCQjvKH4f7MJZDhH6Jmv1/rv8V1b1H6hTLHl5GTWxs4HgGdDky+sJAPYLVXIwayiOFl064
yaKzf+0NfR01O1G0vMggWCLHhhs43XQkwCngouyRUNTT+5czuM7nLuEH/VNpwfPRvnNtb7uhegn0
zMqIvSJZJrTfi5OPv/JE3ZWGFeBm2uDzFxj0wPCjpOY+Fwf0fa1Q8WSxiS1nOIIlpuqmLwcHGtyc
zIAPF73MN0lvSmSOLag1GiD3/OiC0h+I0wwjFv1yDvflmugDhu2R4R+UMCOstRfT00cOcbt3Xowp
eUhpp6zO5Bn3M7EHQdbGnTU6vS6FY+2C5u7lmyXu8gLkrWIp5gx2PLWQOP6aivaum3CMgUhrrmEV
6/HZF5ieMuT039wY1XLIMXpH+hxmYJKG0IzHEugMMARoWImKWmDIoRGu6lUj8ebd6aOTDs1H/+PL
uNzyx8U6jF0blYHePhpJC3vwx7QLtUwDJsrhg10o7Y75lWvmMFH2opvRMW13v/RpEjIQsIGx1w9K
E5oDvA5cyCcCWXnJ8/w+rWSfrzdTSxCaoMO4hPPPGa2QJ0cVtxTMqbiJY9tL0nRU+dexPnJOQ5dJ
8r8vMs693tj0puhflIhee2Y1ikeI0ZDMj4p79ZjvJsPZR8lyto689HjLZfRo6LUSQML/HW0Nftlw
8mcbIYYdgtZZCXJubhuwJ4aZlJrDXObknyWPwsybnZUtz4NyyVw0v1gW5SUtBpkT6REVdCcOVuUd
gT6p2Dq2H/Bd3Fx862qpjSidL1H7vb7dqQQwI2SE4RQWK96fAEIXC2ePe/5ccvaoN6UdVwXccI/u
XB5loFM3iP8Qri62LMZ+cyNsyYmqeTWBPYjkHseRoZrSZgAjhpxBu4MG1h71ulcsA6wcAGyxkWfA
VBeDQdOJxa3N9ovhJoofOp/vSTkvbyBnFPRt+d1septcX6akocAXvApUe28rI1ErCfi009TMSzKS
Bs31RHmhGcbr/yrY+knN1cvt26craw5zgUVSGpQy1+glWZ2QbGkd56rf4J9PR4Y/stL6ngRxoLVj
zmOHMfz5ea3WVtWfKThGJ9cYdeWklutQVWKi5wre5ZKdXZE3+/2RwZy3DReEJCuv4t8/k5Fs/Okz
oLW3grI5TMrEeurcA86CRjRpj432DO8tdFDzTo+DaBsAAs+sWNw4IKB9kQygPXSR/IiFA//3VVKD
+eeqwr8eIzTsZBXCIXi9oHYxpmmLFjtWnK8Zd2MHETs9oCo+3BTV3n98pEsqL2XiV0su6xak2CcN
uh6nnbIt/FimRwTampcT87oZGdXYzG5wlzc2HZZnsUMk+qsRGulSebCbfrv/Bu8O54/G+EDaR9Ij
lICEFaEgyCRFhx7S/e8FW5je31Kgkw3oopdP7wm66cih1CJVH9PmhMkQhgSIRu8XHTirBplaY6lG
xvUa7s6H5ncbopiA00bpyyjny+7sTB97pTyg7+cgZUXAa6M4MIjqbdBJJglpnHE6RJFZC1A5jKZx
OSTtQRQCLhLOGXtxLvMZo9U0DM4mnq5pSRevKHI6K/S524Co874CIZSKlpSPJH5wnPjHanPPVp7p
5bhFZt1ATeOKgkWFj/pZ7fTGIHz9Oupc7OQB07baDLYx4ACOH+wBb6ZheUUKJrNGZQEuDPmg7KsI
C+OsEvJ2S3baXvObCV0Sky1gUiHF3OmOSwryZK0TbJ6tcXNukvYmywd7zToGTAw63ho1Rjc0XKvf
YYc0373HhR2u0ONAfyaQQPr7EXw/CDBADgO3bGCC4r0/GbT7u+HIbygbTLU7Grzj9tSvSksS4oH5
9YGJkyZprijRmuRXTfdGeSaB+WPBez2ONFNAfR/Z7Sg+F9gNNLK1XYw9d1vWGS7H691/pTOacZgu
D0lQMkWqW7Ny0x9yxeXub5QboJjvUlKgLNoWqlanCfbPUawZ7V2CuUFMrWvX/E2bACl7cSNd3paR
IsHx+Iuwc7zivJpX1kwQwVFjCtTedl4BhiT8I/QsNU7+rQRPdWK/axPN6yj82O7ASkmg2BDxMgsc
7YKc+lZHy9GGsCYPLB6bQwhOQ6hNQ70pxYgfjRmtszfkK65RGbdiajhLWrqrWlAuwFM9w9jI65HQ
hLopESB8HWyLcaWKIMqov0sN0isCBakEZqD3Ss3vBrB8aH2HK9Kq7lBEbj9s4ZdGyh0I3qeZ14iO
V1i9Nxw/Ft7CJV1qZy+rEFONzOn14VPJfa7fZYk/Iku60TkkZ0zib7jjerws1KE8icysb1JqFBlF
lGFBuXs1T93A0Jq2IIEFPnKfWtSnTnk/hON1IGj46JlAO+8qi6ZI2FzysoFjIzmc+UvF12QgODMG
QXpsfd3wTcdGzKMzTIk17Y78rhPqYIbidiOHv/ldI+IIT/0BdjLQi+dVr/77VkbLqKcuzBTfvQ0S
JAYcJHJcozvL4WbOgI/9ifndqnluURKOEFxF5mC0YLtfBIMZRK9tgpIgKpRcGoz0DG8LJjgKmQ97
q1Xbq3s/pK8iVy54jkfbfYPBxcqWRAT0T+6tiAuQ12DbwVFDy6WaIaP9rERnfJRLOHgFhSp5u+v8
V+46CNzbGKbnul75NXr0Qt/imym1JzYckXT+lBzEqQXt18BigekCySU+K1ilUjRylwA4gTQecO78
2aPyEHHHxlnFKjv8tGmgFbkQycogTi6kwzXWpd83wo0Qsgnlwo4sAWyLe/JtrI8ThGofEDVf6rgf
Ak896l1oslIcB9vteO5BHEnrZJh2hGrWbRR9a+QCWAFgBwKhqehIH4lFpoDtdNxq7tEr9Bt1spsv
Wy8RvTSp4UJL0ZnvMtbaTzdY1Pf4SqW5dH7S4rpx10FwhIFsR9WsjTWGOEaxEoTC2OeLTmbp7/Rb
Xl/eW+EdNzJVDtODr2u+VaGmxBkk936tZCcxlqcvwtYTkVbZJXbHIPf6GeIXe2QItMDBMoIj0eo0
AHvOKAaIYtN2WzCcbRt+ed0ZlcrRqHH0XrFC4eQNwZSMwTsTwiTQ6qnwgi8i0cDpCbFDN/6WPCWH
JYo1ZVLXoEyCsalnkF8fwI+ZwJFquJMIg3BYw+b4E80QGeFWY4R1/48Tge6ecizNqb7t3zMDoA+y
Tq+whbXk3nSzjMN2F4hXHgUjV2ywMkMk6KtwQQCoLGo59zfMjVUOqfhsJhNLF4byV2cuu+gKfLsM
EENa/bORwyfWkwHtFnoLEXZOwmdPrKJHsXDPZ6BeWcQSfU1Apiz5QZfGOcfDq1wEM1tElmBuJxcf
f6JyR43O5S4XH8Pbkj51ZxwrFKKl0yB8EUqsq3k04LMXgN2sinczo18gmr8md9tigDpF5qGzP2CX
6FRuJnQTj5RXcBRvMmFiU1C8W6NyWeH0qCtoswmFp0knQLk+PLQfkbsE6P9Z6kn4TXxLf5CKAbRH
MvW0sQ4ZU+PUrgVJRLXdJoN2bzGw3nEuYiDfPs8GcGrN+zTh4y/mq/uOmSvTWD1CHeUOqpIfWg3q
UPkIe7p5ol8ZChbPB2wKRuN/GQw2HRtlkthmxkV6AF1/xbk74uTt9OD5emNdApa6Xb+X7zuoehVe
4z15UCXUTCWUmxxIZkF5ShZqpqT68nxe6M8G775SabQIsnjzPPhQ2nZah1G6t1Rmrp/7/Y7To92X
fTbXYD+d1jxiB+Qb7DXVgMMm3Oyp+QZbu3SOh/9l5jShzOVNTEgbyAC+0FbxvpiAzIfpcSGmzOgD
nQI3Pmad5JI0sBjaRlP9yUj3vvyx2/t/XrKohL1qWLX3LFVb1oclcwuebrwMxEauwOFpGVDFNJNH
m1LPt2nUTv7QuwbVGeoMVbVLMvC9eaMOK6P9hToUd8YICyTM2U6+Sthhym1Iz8j8dUh0wHw/6ByQ
e3CQSpa6d52fOOdJ1GSKBcUVbGGJ4uxqNxQYYc+VNyTT+3tqNy3CjPteXbSl5vLWASpPFDmh6GnP
DSp83j2R44akKabSmRLdYoh1UA6Z5sdKfPkQljohIGY/FmRUsFop/ZNZsF1ih+wD78ianQxiRECe
3fpmjhVcYTEnqcuMKXvWkVlpmCAEZJgsbjK9R0HjMiKT+3xYvhUvTNyVyTM9l6H7yR23gv38maHL
3r42W02s9Xswkn1whadmA57DzSs8iAGZ7ecYm3rdWoYaYOGi+YiNnNDODyAKyY8DnaXvN2IhIShA
NbNIsu706T71vgPhnxssomM9YstdspnqEnbqfzsIAnr8FOqUipdCtmEQNqFbPJeyJSc3SepXVZxJ
dvnnBru80RjiVOB0ZOplqB11ukFHLQJxcmfBQjeJEA5RxErHZ36+/xnMnOffGZzb2wSe/YusUawy
S9F/w5yJTT56z+uiyvNFPSsesOooFa4hccob4JCOarwZ29J5/0IbqiWVNbVxMb7peyR74jvxiM/J
01tfUMWlZ0ouVXcKLQkdBRG0lM+O5uuwBvtIvRaqEByRJjtXaQz2/0tl/ZeAgyWOu6kLcJ8tRcHm
S7yC20Rv2w1H4Ch36/vO7Beqzp4VQgfPnWLjP8lUPKr298BH5Rw222CmOXoI59Q/NWSAyKqKdn5j
hEtUIBLy/xtpr8FQ7VQpdxfwFKYrkDo5GX3AlaNgsnNgQ6jESuG939+/rIdmnyG07SmlwCD6C08T
AWa3thI9elg7zecoFzseur0uMW7hbjDCyppNaGyo5MbzD44gXjw41boNdZTG34KzJ0Y3HcRJkMQO
QtfcYjce7b7BjU7KIsZE0yyqJxjW30Dcf2kAlaPEFPZ7henJ8RNOt4ztXgLZyfCG86IYwzlMoCb+
Q/qVs7bTlCv4u0WLr4JauYD6Pi80k7L863mOkurwjkS03wKsfcnT9vYHlanxubDi9tT+l18EI0pt
AT9IVtRQgfTENOCot968mUJl5d1P46FGAyPUzhNC5JpDA0OWmsXUFQxHOK/tAUMCIKGZUJsX8T2p
Nsj/HyFY/cpowwN1A8+cSNTQAT99ZSKeAIQt8BBchss2dVWnCE4YXi6u4YeU0g7Q9QminZcKUwIB
7wOjxfutnShuVk7z8A4HRSSurT3NHVD4aX9pHN2xjuB82ewvmDmgFDmksO5VRdsNKXoIVXf707N5
BUU4hPfpEJ1xg8ZNnQeHI1jyogiV/T2fIWtR/DxxiB2/ngGUtZq3+MhrM3zjtL2Vk7vbodDYflUK
mSufdV0/wpxk1dn3yWje4ndArAGC3z5eV+hmvQG7sOGK2BQ4R91XL8vsjp16juDKt6IBAJWIn7NF
8cFpo81+a5W4KIyu7WiKk/oFZ/Xtt3x43RtuyECD6YcSsDFmOGfvCjBFKCaM1qhoAa/nFB/U3F74
va0fiozOKb/aBCP28FemFcMB6zbwmG8FPR2qa4D9pbGLHhPmHTOIG1Ny6ZA8sx2eYhb0tjy1cqgJ
KJJm4m5lPDEz9Cp96nOKuJkm4TVURFG/UWzrPXK7svBZkUu9E65y90SpJmsa0e9w6VCiii2IOch0
cWn5TSk/qXst+1D9pp3/OhFwV6OkWWFVFB7phuHZCa6zQornSU0rc8ZsUXTb6oUMtdx7pXYwiGUj
RwsXyWX54MDdJpFjx17KQtvuGKecNYXn18rRx9Es6flzHjtGM3MT7IK3mCuT7cDmjBmS+JNozLhS
Z9pKcawa341nriy8KCFVjNKRJHkaDbm5UP54bEBImAqQSNPxAdt0sLPQXJ/eOFIMxkL8meEp0RGh
h3KLKOD1VYACedqSoOp8pZLs7l3hdCGGI1WZrEbJVJ9aWyTTl6U6qwExU3SxHWHZM4LQITWkTqv5
R/DbMRc5C0bJYKVibkBYy7yoDYpfMqYmd+0K+s5RK73Iyk/VPHga+TZgWxg2M4X4rIgJS5OZSCTW
PMMEnBpa2qrcJOQnjXM6QkwJQ+9UEnJTjXAxNSZVMyspLhFiPiW/l9X/723qAB4U+ieFO3IhRR+5
5XDFgygAjFcnRYK4qwlwc3rflF9uUudGqvBRyVI5W3w46VcbcdYWJxWZx2hBfWijOkTjf7+gKTP5
rAATIUO9tZa1aPu6P2ZmX5W+yyw6zPcL46AoNompJOCH9VyALNOqewj7EFRsvyCMGf17W0AIF24S
HSUZuBSdtuLJ++8QRlwclVEdinhftpjNPfyJX0Z9zu1UgiKzyUlH5ZglMl28flg/v0VKp6aG41bX
NGQdyRA5BrBPR7xgrahHrAptOimRhasS6KbqMQDYiVXeP9+V01BhNzkcPcuAervv+SUXAM6YZnMS
kI82xbtBLa9wbNCzH3cuwr6SW48Q8UuBwD9m2CQO3TmrjvjxUgxW1Vlz2hqvU4FB0jUj3GAfv66R
VQ68iE4oaRYOaPXNvjguyLAKJueZkYJn29QuNuBrLfPVADDR0KxKApWNgqLeCJBkot8juSxbjwja
k9MZJERd4Vd/7DXUoXBo4vJMmG0Ao3zGm/2LX7Jzrt9raWhL9NLvva55wXmxnstkmxur+oH6Djk8
a3OjZrDkBFlp8yZM2UdjsZmncfdoyumbojGwNPslhnqMpH+TnQMEyj+JPkc2mEL0d39H0oQYxBeJ
KpD7sTvsw9qB38MglUGIe8xN8nM4P0qxxf4Mqsz1R5s/qZi6V/5EkrNf8WI9HcB6OhmF1g+bxgaF
OMMAlpA3sK69V4dRiv98q+NKCq1mIF02bTl7SykvQ7nt8PAlQfoFA9HXau/KkeLqeBVyG/8qh+Wu
yNw1kdlnaDXEq/Exnl4KDcH2eCzDSmiRA8slV6WoS8WA3xiYpD74jdInKAb72a6Co/asahzjbMFd
s/GC4bStJUgIg6AqsluAnP3/j8dkPiX6XvsE6b2URJL09IcrOomBMqQIeQTbACDd2wTI/UMOreqQ
uzFfYJg8t7/QBmZoSSgfjbT4x75a0mzAgqH6EphcMUBVibpYt64a4Wk57iHw9zbtzZb9M/KXtxK7
QRYIXecVjk0Z0NeuX8qie9TeFOGQL9XYI9RhP68YPHQjOLN+aEZCaXDLSB/nLdJtV/wlmb0EJxTA
lA+4r4b+6PcpyEUoZtuk26u4dTJRq3Vi76cgy01xqlijRK4mGD3UFuba63hUjMkK3bvtHlWnXcyp
J3Wz339TbZwWJrA9XdxoHfAI4c5XGtP6Sy5hFpZyzldbDH3UeAM3XZWI7OzVFsqntLEpEKgbtT3S
l/+AGeAtVplIa4DvtmYucS4FASMnhvt048MwIdXea+yATarzJ55vtPadKzhSJhmbbNRaZ+fdY94v
H7/xGTu/gOcff66qqPyczVwb43pE7Xa0+qRvoxcpOW2rsxPmnAu2uwPzeBO7JUIrNFxIXoD4qmHb
er5cPJXxl1ZMoIXs2Jqy2oLj/knzJzJ+CqUkEJFwS+SPdj9xLlfm3SE/sonm2Azubi8MWOY73IUQ
aMiP6nEgG474XsIPg7uO2XO0/gr8TGFpmqggYDaAZX6epIGSAht8CgYWnyJ5ZCu6yvECQDER4qjk
4I/eKqSB/juff0/FwDHmqap2GgNtJBcp/oH1KY2xSYsEyxZ7pIx38EHP+jKiKXH2lqXLF6Bsp1aP
WWgkh6AyyUiK4lyRQBIyZ92HPZiI6dFGrZvESdnDgECnMGY3sRahFppv8AiHTnxS9A+Fhf4CF/1l
1HMF0W+y6I6SdOv/DaJn3kyC8ocK7f3OM7XDClNieB45av9ExUjRJ5VTJ/6s1HD0MNlFOGzr18hu
93iUdumEwVwPZh4pcSFAYxpwSj4gW34BqxzsZbSzzFcEyZSg6eRVBZ5mhamf8VRFyjc5yV+tHTdR
1kCON4U13ttemGyUG2MHPmMEB15SMzCxY3KIIuy4NydFC5Vqi3Yiwz6OAiArtL9SLF8DpCt/zZWQ
w+Hi+x2VHrCjnf8NvGmsieAaGm5WbIQK+JhzQNxzEEG9oCLlm1k8bOGlD2Pl5X6zI5spPaQ0XAnz
R/rZ5J5DX5bdSkbldbkgfc5NjX2uEFlmN31/LFVFj/UZx3zDDYaza2rPP1sWDVRM/u93BC3j7CiX
e+cstnaqqlpOMWelEVF2LEgbjk2Q9EC/TEjcta2RShhakiT0O1Mjj/+jDPaaB02Co8ABPWVyNaPi
PCQ24zSQ22dTmWKAhj5cCnjqMGrHeZa8QJhE1FIDrJi1yoPbTfulhZmzXdmXkEwqvm0L/DjfuSGc
LWCtcqzxyYOK95Axbr/rqd+qLC/Gm8Z3msrZU3s59RfhwBk0Ek+TAetOXflifDS6QyW6NN+kuo/F
3u83XD7LrqT7WkInTQtu87E91YtpO0qmOVvwsWLw4I4AngvehNGs+g1wxGsAlRXgNjuOn66sz4bH
EI+fNuGz8eqb8LMw1DvgUwaPZnxkrhx+e8SBa7sbVifP8s6HQP0Xy5l4/nAOI638+Zu8eif8OGFi
oz5b7sjTb/iBBKf8ix85iz0SexH7gQL2xJzwZfv8gNey49h1s/vM/YXoppM4la2jZGVlZcUKSa2y
/XN3f1Ha/uCBbpn4uLTi/y715ZdD6ub91MAjSl9VRNGbi1GSRFrbkBhziepmbpblMMkblPsCvnfo
DIGCXEtQyseOMByeWg4d48JVzO8448/YBspMwSPlEr1JHmSUqslN5pFaS9vD5yanN/KkuJsAKYUJ
kFNUUMIYmQUN2CmXTYthHNd75Q1bgW5aKAy7CTaCwoDekr06R7k9RGVBc1D9El1vZZ1qkDh4srEU
1gy0QpzuMFmjv7NogmXfxMkcQmPKyOMnceSfu5C5WaqQLJZyjY/6T+lgyYhrojquWcAso3w/16pM
uQyZ2qCLIXtRyoTr1izhb8k4HaI6jbvEMldsLsOt4ZZF9SGrIbRhof7ve7aVH4Qty4E4wZ5uGqVD
nHENO62/TSnuWa9UwHqfTZ/tAJ4YO5w6TYc63x/Ag/ydnR8um4ePGa0F/AJ6PspKLcP1nQfbyEyr
Sp949dPS4T/PIFHSZUxzNj5Ig0Qr7lqxQUNVHvni2V2UAnRSkBaMMSnT6HQl/gw3VpTgGJTlG5mt
RQETxrOAE8czNSPTotnu36Dkr2OGoy+lwg3cJpxejfAgvcGe5h/gBSlOE63J6Sbep12R/2dJr9h8
xgrzFDKDAzw3Ue2nQ5Gq01WwJi5Igbk8vgUhQr1CN3Ffr9/DBQYLTs2QpyLMxhGv44mfhJyPUKhz
MVGubeDjx+7QKfMYqjxZ4i35KBwo3a/k42MvMG2v07JWuHuCq/A/tP1c9gnggIAIuvCFTDgCXaFP
3cFYD+3xnDDxZ+/8RtA1cI+u8fQxk12quHJ+1/CLhTE4DUyi3fzorzH+g7qmC6KMD+ekNvl+YzXI
OG0SpyHxi5k7bXpuKdI8rlxSG7GKdlKUzIsq4+gb4J1nE+fBAYHY2RkmC+ooUgDNG2VAnVLR0C09
I5NRkudYXcN6yRPw1pRDNaeV7MIzSeb2cOdxawc4zbhkDDPnlOC8bYy1B6uceuXaPUgN91AI0hld
TCFEKf1ECLTsykY9lzHfUuksV6A/Hvd617Es72s+N2xlQceGbDKeq56N+2gbFQw8fRFoiCSQ0lcz
mMtzDi9Km8O4jqyQoah1ir/UPEkZ2sbOsPx3HuyVV+OwFHDPGVvNHKBrHHGI2nnIcKrJLkpb4oEi
iM6zdGFDJM+kwNa+Z7jmuxRKjJ8qITjdnVDWC7T5zPbtoatvXpWsagrkx5xy9yk+zFs0Qu7iqUt0
2EsGVXWbvHQFM/2PbxGmQBXaeiwA91Awyuwt3h2lg7yZrr4x6bZ9R+T5k/qrIiwFj5kKAmjzgt5C
MObb4HnEqck8i81y1j/3lL75B2ZaG2RzLQiXif7Sr3c3eAxK9E7LVQmTscZDLDZvtDQ2+HBeRc07
oM3F/MBEuBypIZLpTlPvokhQGOMVTK4C5S4zF5vSpaSX7IV6kPDNa2aHF/hNubO8UA6ffflgS8Mh
U0xIbGbUjEKKtM2VDepHUU9XG7I2FU+H7mWdAz2KnH2kUQbXlHPd517PWAGixRG9L+mkKUast0So
hXYW0e5zzyaF5DZRfaTnytHTV1VsimKE4WVbXiK8mhNA9PEVBDcNrXdd7QGqbGSj+dzWbhtH5U+k
QY7hJ4w9f8tcU15D16TuRpB0n9e/kdYaf80r1pH9/HeyPpRF8xVVZVxQLurSgy+PjJfiK0c4TaPN
jc2xUDYOWJ9HMQiork4h/lFYYxU9W/DeJWEQJ6pJyEP586GiHnE9lo6f3A5+/Mz/Vry2hO6dWwvK
6tetYXohohM5LlMiLRuMkuXVGVzrjQYSLgPu+h+I9fPhgBJmTUaC/UpaMbdxo2tYe+D/Icq1Ek7h
d4d6GH3gZFk5mreqGIv8XlBhypwHdGTwBspXlHvEhjyQtebtwBhiBYt5kM0s78mnC5QFFfUK6Mkl
Gi0ceAgd+KnDPNPZ+iXxjRk6cBaHZ6USOUVhHF1FqJNULW8foshjYGoMBQB1HZAz41RuH00j8D6S
TkcgCUUC3X497ruAksESUMv+n6AbRW9LSrGW0XOTeSPyhsTawFOFvV2x664kvsMSR03H0xhUHpxu
kUHmTNg3ZPnhgM6vDd5Awn/7zUAwipix3E+neNcgRxwQhgYUrb7nLS384nC4s/d7gA6M3X9fPXQC
/ehYMkd80tgu3AdGmJ0NyBGK6JMRcMUEyIq+4mg0l4Sohyh/TESCOeC04dlMvEVvin4s1qpvCbvO
3A3csW/Q15pyegKR51Qzz8NcbiOAs9k1a0Hjqx5viKhh7iqJ4Fbkgrrgqm22SDqYmJr6BJs3y3JP
P6fmo1NJVpiNLx1Qhwr5FT+k8elnzlZ4eNAKsnPXYaVF32hv+ehzmvDNx+Rkijxvaw1pZ+ZlFzqQ
DDhOvULYxaILGj5x8q0BV+GABia2SDoUrCFjePaQTu/nn7TtD4lQVwIKImfkrdD6fZs9kj8uF2f4
+MZ48K72AKv6bF3Mh+MD3oFMA2KHCSQ4CLyKcw/OvhlKqxx308VOSDpFD4qpDZOGwwhE1sOkFvk3
4GI8jfkYpOTQoVB9VKXaGr0rAAqJBvIieOmHzGdLSbfFP8WFpgALS+CQHUSfVtGaZuQiXuzcCR32
XFyJc2u20Qyq1FOkX951IR273LKynVpTy49PaR0I9qzHe+3DsXY/eoE++RHML1KrMzJnQfwEKzH4
rngkZ1ca8zbOhF1aqJpob2a6vh0armjB+thLDnXAgE8IlMw7QMyfGtfuIY9fM7aqgFzBNa/ModoA
fVrZvi1r7aodnmeDsj6bQx1CvJUj1H6Slm6GLoy/ypfB/LWkHpIt57qUmISNWaBvFZ5v3bwOBn8x
q36FrY/23COjbRDz7HdSFHP8NWrZ2Gt7GI92NZVkLy+gHw3LWipSAw0odhmcy9/iUT1q4ERy7FFf
zCarg+2YpAPLHCnVeNBdvn3js9GgHFwBweAlZPGwEqdQ/uRrqUXJ9Tp/kD/bdzzAPCZy9IWgVpZx
kmeQUkFpqheZn0aOGufnzgAyeEpNUJar23Ken8sKfPuDvhkWBMFeqfhfOz1V7cEt6NLrzpZEjOrB
Mq2mKoS2boyCvC0L/F2ngE4vX6P4lowgweJ7SCj3iLbgeCAAv4lD0kqTAxV2YxMFzfwai/YdTL4s
/rTY2ktOQ6C8CHBXQGjyZJ3FfzU/uSB1yFUW+Wxfj+Jld1uCNZKE1+lFWs+WdJDeb0wGR50OrkLZ
XhermhCjXoxWW+E4VICv2KimWMhNaHUXxJk8v9bwX3E6QAM/OFkXr2aacxqg+JPKL45vF6WYt+0V
Eg93XDPhaTc9H5qr3Ct4iKg4/PEWe0uvHCocK8JQV+c9+gN60p9paSixrCLWgLHirrY8HRGi3ZjL
BON3nhe12Re+dmYA0IBznVOlXkqN2eeF+nF6tz8V77IuD4+IuRuOKFU4DNrRpRg+7FOg9KhP1BJ0
ddv5EU5oObH9Z4eHJiwz0RK0NY4WxIJ3bJvDD5f4zbQoX0F42EogjJqwfL21FQQzRXSMXg46PtBD
lattxhECNXtYim9G7ytQkfJ5g3Q9Xl3Q8SUxEaKzrOE1Zv+Uwzv7afFBQBpyAv4hQj+1KNaSu3oT
kEIQuGPRbpIbm9SzRYNIdsu5SgbJC3TGiOFy0rkyq1uiXzEBxEbt7JFCTDWIqXD/jsY5eux1QTIX
al47SFT4N8OqF4WN0oq+W/mEP3OldkY5j7swMz715WAwVvZkhOWqy642tp5aEpNR9nnLfwqodnFX
lL4wPuN4rGYbc2Aj08lVWm5jwfgGcoBWMOpnMItk8uU0r6KPo2uDyyKmrG45eLhuMS2YGftFiPdB
Gm/9v5xIfB+Ms/KH39V2p89mEyFnyYIt61WNZJctV7QYJU3cZDao+Lv6QqIE+RaNXlFPwU5YYphS
7yAnXoZmq4oXrXPZMua1JQE7Vq0Suh8twloCgck+2JGZAmVzkgfnNOfd+6Iyds6RGZENz+9B9fAb
Z3+uyDycbDys9yr89/1WpsdCzvKZEUpMyYDye01DcrS3bRS/WMTBBp3Zy8HuA2WdoqqDNoDR2aJV
WaQieoQEzDkWnejrR04cPjFDuI4TC58kP4sGLkJyZZINJwz3ONfivWhaigEvgTstfT4c+gEVDr5y
HXp40AJp5b9Up/ouehhE8mHzDxv9ixUYstMNtfDVdLwhhd210AAaCZVwrdv+7U9fhKsh5lwQpEf8
A3+3fPNucQkjLpZsKUqjlcLd4PzhNVNoYslH0msN+gQ8ikpeaniLQyzUlx9Lg2OQWmAT2H/R0AHh
28Tnn2SFpKVv7yfFQfWdpnhO5SrvgvaIjRjT9mNBOVttME1Hvo9rIuBXkn9KjEjRgBYfJXWodWn8
8ii8/77UqrdXWepA9u7udw0cS33SiYi+2UHsf38RQqqs7wREmpPpDb7+1iPZSoa12+0dUpclu/TO
293i4J7xET5ZwQ9DOXt1gFSoCeVGyuwbssWK+kNsj6f84prDApU/5Z2dNOqElmzhmMEOCjIsYIee
T3cBQXPubeRsbhELQ/m9ZpMiF8DkKJpzrUluPu4O9b436UV7ESBrisOZFsqbPB8PBJKhHNfNA8S1
RO5+tepoRaxeeF5zns8UmfB/3VSZdDCQ9pHrl8jhhu/a0qEXFnNP+O9KOrxMVq4rNvk6HsYWIdbW
MufS+jGsmMu3AhjcBgMinyOX9F3uW0scw8v/n3MfOt8Plh0AAV1RrgfcqDLh6IDyGcqesbtTgbla
YUsuzN6+phGjIPn91TbaPG+U8mbP2sqWIavmeHKKHcDfj23loeQqpItIOOYKAUkVJNPTrhXKHg1F
91+KBRtI8kkMRuHkhJiZHqDqIAktD5U37CopdN4a8XoSVFZdTsyAckf7MFt2ED2/MDxe+Q4B343R
IdfbCofpCm9iu0sn2SxfOYrfYtJUCqgPEMbBwB0A9LmmLcNFtKwVKu4FF9TQ3DZjMlsr2+hu8YHU
4ySGqcIHVYaOLUN68qTTQGS/iModRYf0v2bZBqWhNs+LvVXFsIcNVozHblpuaHG5vVrSVehWIc0s
eLnCp8/+3zHqNgMmHJvA3qXX8AVmmoh3yXFAX6TNiFxIQlcvgfZRGAg5dv6IwZewWGMemzXfSq+H
qQlws49jQynwXmGB7bdfz/tBxbkI3xxkLni16/xXYC7zZ3AVNvqJP0J3BV4Twh2Oi79ETQuV1LSk
Fa430f+fIUOp61bhXMYP1xCbGClTowdElYFYJjNzRMXPMegkDhOGK8LxpsnZW+rFnCr8ZKicRIUk
RO1xqq9ZgTrWTw0A51XnDYqY/xEZMldbIuBETKVoN+GhZFeSrOqtXDMe4hBFCzieDDb6T2xBK7qt
d+/SlqJ7CNz9CSYlh9BL+Cw+Qtkmq+OWUvVgStEzv1nRMrIj2GTRhtyeEUsZQ/qKHi0XhfKbaqvJ
VhN6rQBBYqoppUzjU0FhjPbEQbajwu5RZ0dYBTywvuUobfAe4O9tzdIal6vJklnXTgxFKwkz8jyP
/mjXrssBxyAPMrEe8eDV4nCeuLnkG0jWkkwv9mqKTB0dq1iK5RIk6FmIQXE1M1Mqmoc9c700K5v5
GkjrC8rllNENtK+KR71kbHIdzILkoeilbAbRLjHZSKCfFrzoEirCEPW3Dl2rfagAs5McfIS2REpw
Gpq7P/U5GsBbDTfsd+pgbW8mnuKvTMAFUwPlAqzq16EXP4oc1BMtrI7YBKXtO33K3OFrsl9cb19W
ryMSg56oasUKO+fAdX3KUmxgj+KrPrdzSJf09GaVM5jEdkgdRqqMrnR0WOMlOeGdS8SUWWjld6fH
j3cp3jb7/Bfyk3hwTz858+SxphymLSrqr1r4yc03RLFLHvr2U1ceGuXpQj+zq7mU6SJ0j1yAmuLX
ezBKa46YYDSw9rq4/coQMeOoe0HprMyCAmhUiem0g+70VnRXcZfDce4QTDAjbNPH+Xzu/2o9k9NX
2gQF5jN9tLwu/kG7K8GhB0eVOto85rd6gNYx/1Eq0uHybxPcmjKQKf/uu3dRd0vES+cyAP5wEjzi
ETKIypvBPu3C0r5LxW72kNSlBKB49MPLr55euXhDxQcuX5S8JoyhLiUweUQ/Ej7/HAm+EUBAPit2
jj2xlo7Xe8YRtTWGem5Wo+UP4uFLQoDKXX4YcV6J84k5oGsW60q3kHYHFXtBES+4sLrHA+aK/D6Z
G8YZPt7NSxhgwISibqzXZpf1ClAmaEfrGtCWLSO4g0ADoKG8ReZWbgqhxdxdr3YwHUufzncUam+k
L3uPOD1BXd65J/rLLq3beIH7h2v00SQ/Rh5rF31WZgwhglPTcoq6Ym0TbsR6rCaAPFwWgoq+ov+V
j3UjekPAILG64GE2q+iSVd/UAJdbAwiXRQje6qSeLLa0Xl/EJBkCX0ANMtv4JM8RI3C547xzd2Av
1MyRkQXPkbr3WOcbvkFy6ueY9/8nOqGLofYqpax6rzlwBk8wsEA7Qj58I1uYEREEmsnCxY2K+lLZ
yyCHX7za7O6abjxjk6qXZT0byMGlFSBZk0DZ5wLmVGVJRxVAIhfnxDMUQ5KRXCSbuVQWHZlMFFZ+
oMxQn14I5As1gBMh2bhYHlF9tIfuXGOV02yRQOMmVX/eJ/HHg99Ul9FDVZ9ztsdXPFLkuVl8Gf06
GlnvdcOphh7A86TAKO/5s8qKl509F76Pqt+ef1vwgnEIHdE0Vc7uKgCPXjBpBCpyka/K1NdV3CYE
gXC3UmsUVCB3naWPO9RwMfBm3dQxRYY5Wv3wQrSMZCRPJpBnyHiuDbt/DsAQ5n/SfiWziZo7QVMI
zurRiJ6d1CB5OhPLmIrWSeceRn+Uo4L3Qehk63w+D8uOIn2x3cME93mBBruEVJrgohX0r67e2Vnt
XbI2lKl4rnRBYnasUlyGmHfz5eex06LweDEkqy8hJ4gLpfNrcnKyqKf5f1zf3KXvKEJAXuho8ZFU
M76jt5BN/fvMlzQTe/55JuD60M/mDbIbPS7XOVh0GYH6f1CzzYwvyeP6flp7KzfYVwQK80JUFCvu
UCjxXixrrCtGuwGeje3kFSwtHF5bFI3AApfgvbC/WLtSlXX1oF+290d/gSZjN5ZoHK6GZ+ewnOL9
T4/yTafm9SbPacNwZRWSVisIbZxQokEAU7NpMriG5AupdZRXuoVtbe8Y7x1Ipjie6atu8518R9rV
cuvSNopimdo5oTeASVHzS8vWt7zSKjnHkx3ZSK3Ka/FARsd4g3JQHus5NudX9knmz3gjT/04QuoW
eRb2cY2aTLbAkjClM1XDnOYPJTnvtN4muGYOsKbsxV/45JxPFm7HSwI/vlol8x3qNDEoZwkNF4Ns
Yu+vw9RdAnq11nmHaY9TEoSS7fjB8pBQ0cX134Fu+X/bZtQ+xW8DMmFQmeGndDICS2ry5ohWijFf
GBPKAufCipHb+mNZYi6yt7QEnPhKtyXj5Jox+jE/iDVJzFqTP3nHl5mPKsJw0TPqA+1HPkByRtPM
7kW4j2yRL+IOIkNS/LVSxf7v40sUqmWkhsdRc76HUrsJNalLBa9xXZ5Xnb78ARfwboH92g5LpR1O
FwyskJiukP3wRTYmIwbVt1V4c6GHeef8CO2zmGXoFpihEHwXvGoddour6n37TomBrhhtY5RUJGYI
qr9TbXPYK4vO0RJElmFY0egbPx5NAFU6DXxTLam7mfsSxhpCfsQZ8wpbcdQfMSL8U21oHOO7RjRP
MkIGr/K7i8wQ8Dp9MXw7kwIEBf46hPQsUhdlm/jlOEKR7AieM/v7oYrk3i/vUWh0O0hDgECjtsOe
gDotahM2KpJ1Zptg4yD690uSoEe0T389VhBKyTXczo7CBTzXPnnuDXpFJs8ltiz0SR/12zS7e7J4
LiN5ESU4D98DrCpg7SevMrReXk+XIsBp2kwWdYzo4aU0I60HX4bGhj6M9n1SbcZ8e7ZtMzhw++dP
LvpXAAxM/9g4sYMAiTrv9p6DY5dxX9hjEyl/2vtD4VLmn0My5NVwYFwp61uRzE0+JW+0l29HP9L/
PoJ7gSAEvGfkXllV0XUc+uQiH0VWCKagtS9iWBwI2zukSK9BuLBK7L024C4X7MFC4vSgzcbZRJUT
IHL3hR4vbzyH60iNdPC9QFW2kOF7M7+CNVePv1DxRUJyn5Z5pvIjWknU399xH9rFr09PNVqsdUL4
Yq7V2rrTmUyJ2WMaJOUfzUMjHcR6bulEI9Lb62CxLIJV1fkeH49PdfUn/zZ3CDJ0OjwrMgcBo3TI
5Ii9ATAuyVQXcAU7NXc+zNx2YnOTckKZLbqVRkDmYqNWdmUuiBImq8vKrq56oUfxX/Pgn+gSSAzW
SP0k+mhsxZDhWcqLCr87VIYBrGk5larfCWUb+BPJILLomqLo2krx84jdhgymG54pUB+nhS3QnKgk
zp8ION1hzHL2Mez7g+69xq5yQI9Qw4QEd8JRuYxPsnSt7Uw4KaFdQlJiTBWFvCz3sJOjpbW5n+AB
QMm75d2Wdm2CH5k0Y8P7UzI4ALO0vDP0aGjQuFE8hrsWcA7Xk5PkKsDV3FNkfHK/6JWGp2TyObgB
3wnv5OWhgimGLvQGppDijAE4IYs7qV1RDrsI3m/T5ElyLdSQN6JRXaQymWeUVG3nhHTMI3r37Xyt
owz3kCnFblTX5ZtvD6z/dJ7Xf6qlVFoMLpByLyQh+ZzYeePL58H5cOnmIc3CFcLqcVpW2D7IjV3/
VzO1IFcXrNvMgC+x6mh5Y/vze29wNo1XmOr1SMKRpP/mUoBobgo9v1afWQc/8Yp42iLrOHVnXMmQ
qXvPC4jw3rV3fgxTxnBpsuvGYb/uxRa+aJ5y9DrhjYIuof/7ZRHoef0gZbvY7HtFUoScGmOYKg4L
V1pMwEZGKxIWvy/aP15nyC2eH3ylLG0gtyRJjkNcUv3SwDmbOL7L4gedBZRmVyE/a4tbOBUWgZPm
Z0tij4YUjiIrne4EVRF64W1Q0/kAyt18Wnj281NLWOGOELQRS1LXYodi9FIPOrVQv4UnjeaF4lJd
kgsT98GGj9kSNrchCh5oHT48Y1ndm/Jxdc6ZNiADL5EHul+Xtysz6LA2d1mSAxIx6eAVU2RZkebr
bv72YPnAb3/B6pWV1Rxg+hleRFM99zn7OYW8kHyzh+qblIVMWCsRISvtgy+6hiwVEW4MeYHLrVdF
g2bTQgSfIkrVYecBk0PYh17jcVAHWsaT7dLyn4+FWgJbxNSCVQEuEyk0XXB0SejdMgQOXib8CpE6
5yJOuLYuaIijGcZ+gfHYCzAHT8HkyulY/KG9wmT91AlisewV9KQY4OT0L5l3wu2iM48wzw50NAMZ
dSx/mN1A4S2l4KTaYYaAZQixfOrSUVDkxSdrE6PZaWIKqrug7b4385mKVtVAdV179yibQHi5JZN3
ahK9MERdWmzs6uHW0phvOnmhObroHQXw+u6OiTChsfvz+BZrg617UWp21yOREVh+glqsPSFlnvF+
+T3OKYXD7jK/IWG/gPu0aJrwuqTmwMEBrKU9nTxM9cfAxHsoNvY0s1ODCEXXdQz5v+o7p337PIRF
xbhIB6QB8NMIBRXGQcJ4aBBmlMpz1GWHfVPbZ3W1/4QP9r2tQyiv1uVENlC5QJqrRIJs3Ni7KC9B
jYGFXn6ov/IQLw967mej6NKIMWAy89Smq+1WF0u7T/u86hBT2OMsteIrPJ9vUSdtL0Lb432hebSi
NK1g+c6W1ZI9UikuMd42lvodCkTuJOCMojQeoW5nX08vcLfQaEYYFj50Qa7xMsApdl8PCk93AbRR
9eAbfHzof7wPDnyWEhH+n56MXPajqZ4nZW3h7nHOOc3n+Pc8zF2Ku18Tu2Qyz0qrMXxEW1MZYuWe
pOFyC/pZkjuIWxtIwHTlwoPou81HlkYCgV0ZbY7PO9e8yH+k49Ed2k/OJMM4Y4c/I1l2hyRUEY6g
5g3q4p80e3vMwATHe4Wg7pXYz+g30EtTKX0IeQbhCglejzN2cm1aSXmMET/Mn69Hh2Z5iRQP69CY
Xo6Dym0DyIRRd02z5urXmPIa66qZ+JrWSwMAB68eEfPNAoH9NdoDv+Wm3Q62NXpPLPCzxIXlEUYP
qdJETTSbMo9zYnQ4tLc11qtrwFWTYVGgV023jYgd1NWOdQYYoV1zSQ6BGpHtbui38r3pxQK+Hsof
LIyBAyN8YZD62h8ERyksoAqJi+5w8VI9t6aaySeSe7F23/Nlz8PEOtHSWZWo5aayyq/uXnifB0IX
AjgxN7eiui3YmMmdws4gYYI6rQ5C2xdSHuvI760X1VH8oewpoJ6gdsaQIQw6RCEaM80cYrWb2WiL
cq4X7q6IhEbu5+GtwlyXPqPEReZLH4zINFo1CIl6CS0CPJfiDqb16546XRJexxjXAJzG35cZcZvT
T8PqWH7GrfcxtJrPxqnsQHpJymAypklL7OBYHgj8+E4tLHurQbbpmpDbZTDYVZM3CFTJ+YOr8O7T
PoVm16uIR7/1eQZL7UncIxQUcADy8/8aC0Sh4zmjuLxc/MbnRefV2KB2E5rkqUkaICtexjfwZSvA
EA7GnvCff7X6k+r2069kZruwoc0E2UlBR+Yr5yI0hzYznR5g4vGKyH4EIyggfjqOjpGuUpLZCFty
fvLsQEDOmd+EcdNFi/nnApLyLTON1weWx7naFIM4Wbj8gnncyFbyghvm5c5YNCvfyGFeS6kSlwN1
e8Kg7RRnr7Z7Vob29TG0zU+CrAUrFvap21GtUhbIt/UTDykjcr5JZDRmEYrQDFw1HAc9fAK3BvxG
x9/vpDmTyBOgu3l8x5nZXunZwkAAR8SM8a2xBaq28adubhanu2Z+jB3qK9AmllsTNY4VVi864Wf/
Auxy1/q11gDyfsi9KCzi2aC6P0vqrP+ew1r5VW8A/zW4J/SWEbNh17oLBC333hAAl/cZRvCjCztg
qhnbORU5EQvesWdlWiv4GP8FOPpLpd3L84cjxyF8+5HRoUy3jiGHS5LHMDYDdYBzfIZILAgvin62
yUOiqc05+xKreMhaWQG0fscK4LU6NpcX7n7YJZwLNY12cW4c1ekQYsAb4GDPwEl5wvTiqeDBvese
zOF7E1Z642jZCptF/cMowvZrlId4fpW8fVWFA2jHwgwSekgM1gr5JOOMHaoO421CqJPAm5y4UdeP
Zyvw/ZsyPSSKWrJMkbIfrBwHucQZ4mjFwLx9uldIELb39Sc0Guxj5PDc6LgonS2zJpF/Dd5Cgjav
XlMGk4js1jxGCppf92dDx+5J9Ew2kbnQBFrGPD9qzP0lp3P2GOftSQZXDIF9sn7+kvAHUyX2zSYk
RQcqCboNgZS0LzUsA4s7asWkrc7Z9cr+tk7tNJfYRfFvljKOxpUnZCY+evoW4F/58RBxfRR821z/
cRtUdnxjmQCvaUj1Pg11dWKMGYADt7xCBouuFcY730+4OGNanWenUU9rGXOS6WF+Mx6ufHJxWpR7
sH1PCKviKSBMCguX7A9rb2efNvHUNZnApYkJ0rumMDZriVe6XJdgR5WUBNqm4o8vJx+YzG93T3I4
9Da0KUw9yedLPTUJyQI/8PTTuV4Fl9d0oUxtnugBpdKivW3jNJrqbvZBYE2lGeLPMLd8URW7leMc
KAxo0ED5XZQAc8zYxnz1QU8WI3mik+hXDz3RE9hFRuTKSGTTHsAwCnaYN2P0/Rjaxqb0XIrNUJHx
7cOGvjjlPKFIRFwTdA7Y/42FFmWgJKD1+/y6N1Q/1aldY9p/DN+NibkuoRnYqCUTDVso23/s42mw
axOBY18dBZ976x0o3aVmgAJ0ztTxWbelbTrdJdpRQIdxL3uq/br6heHLuIsMp+b3gfHOKRmVuKGK
lsNDL9ITFiHbIvzHZMt08gVeFyte1rTYeIw5KKF75L5aGY2Rnp9jf7ODqIaD5hdftBiioYcy23Lm
reNaASilqvhQ1g7LvrleH3vbcF3ke2z13F8GDKPtb1WtZVHTgYNW7zsiW6Z2BBw2EMDckvsPpfmo
an/X058/cHjCkivqKBRZ12zMoBaMYiFutH9HJZfeWtS3qtA9oBI9fEFyzJXUUk9IQ3XqIDso8l15
LEsDWAEmECjPJvfbnO+vwU4y5TCHdcNWPEEVrz9+T/CO4BVe0w583+HTsNKITyZb+AEHVtHFUdyy
aVAUeS7/tDoafOpCYnJxHQe8iKer9Fqz0vyHBZNnrKOUQAmLCJQiHWpb+w5Pq+rUsbBcM+WgSREX
ImTZuhT0WsPAQ7eQ4eUljvnnQ4vFYGFVbBkfjLapkfW98s8buXEszX3Wqhj03bIkIPCDtX9AzBnK
hOm4L96VVvZ/jV3JkWUrbo7Yh1i6EwNlzsGlQF9NMyx0jU94lsMtW4vU5PK0iBi8h34vF9TWbbp4
CR/baOh1Am5vtkKVNGl2RX+9dQw5VGp79z7Z1zox8rBrSq+44KpbO/EMxe9LjNDyEUzSFlfdlUif
eb5utTcq3FodZPZXuF78eMPscJHd/YLP578rQxjtOc0KlJv54o4c93dzWTL2w4WgS5iY2VXO8Og6
3rV14LL1M0xhD37OeMCCyzcrst06jRsAFWieZcjIMDMtBQEEjJTwDesxZHL1W2riPWglN5DdcCsF
9HCCc2AI7ZtnNi+s8wS7xvTXYuCfD7iKH5/e6y+oZHUo+lz+xxhABFXsOoaVP9Vycn3KBSI3+Ej5
Sc2TX8CJCWjZUKPY2jp0VpMJXyW4vw9J7axaDLNBBhiKeFG+eAq8JALQVuhwp6T2a6KETH3gvLFI
5LhIGpPbZMEqizAflHsLLp1Z5TcNRT8FdBZEsN+dtEdL5YY4/ge+abOWcHlZA6wgQAZVDTzGC1Wi
5Y6waAThir5E/Eaxvo9hUm3O1NhCGZyI9/l9FTnwmI9s1XILw6vH0ehXGLFPrO6e5YcZ6tU67hQY
mojR4j+EYwpICIAotZ6OmabQ/19z2eu9u8TxIfntfq0LDD2F6KIVOERIKSRLWhdacfBK9w4hFkQp
0g3HJt1Ls/Dg2UCDXyh4iddWDR0xWugYot31u8y7CGhzPvqNLscdbOCq35X9X9HUcvL9MD81Hqxi
+JvLU77GCXuD8WGQKQfc8IwAX0nfh30xtxOjDefVQ0VMAEAoQ0rjFXuPv6Eq2m+B4S9tfEBlEDqg
06h9n8NfNiK5tXRWMUQklYzLiDLjvSDwl/0m0UaW+Wz2tAWWrsxsxDzNAzL4qGpxQemU2Pw4De0r
lVWIn53t9EbSsJ7wfnQlnRQoIy/XNGmtllcmgdVioNFaxRC4vcg4FxdHUsLm6VaKsKyTJKyeFBpr
r4ZwpUtOQ3IxQLWzEug97JgC2/UQyT2D/C+irQQTBO7y/K6J0lHPuzZiR2JBB+Z8NCCb9nw0aDqq
D6v2OQDNmL/0p4O9BY1Ug3fL7kD2AxE0lenGs2iZ+845BP363X8kYGhzRnBwVKem5nARA1HkNMkn
cP98ideDn07CheMKLFjPikVAJe1gSWgKVlSgszC6dz8zuETg4gWO6LEQQXXw7k2Xq4AX3EqW6GKx
uJwfSYpjm60NRhglnl8GD8zWdnOlINwSwBhNxEQLdWqHR4DLnIX5LZZ1CwmsITWqJ2EErGIDyjb4
9Nx6zdwIda2crZqN74whR5H6vmYFrMl75UMw+tUOSW5uHI4SnwezLODNSgrYIKzHSzVFxWRj7qMH
RmQUg8D1fCGKVQjdCsi61NApYrJacgi+za5CRcLKv4COQmC1PnsMuOUwL6PKDwafvYgdX+86KwRp
tBhfcBFR9CmJwntBx5uEYHZDqJ4McQi2vH/knf9uAlmaD3+5d1o6tNMG6yn7sYG0zl1hKu94ZviF
NFt75lb6aZEFxorJClPtITGXqlBvajPW2b5gvddQ1IhhNG6McZfSmGjEHZMQraWVS67jrULgMDHu
I2ptmWJlUFGyiXLaOStKlsMkSiZW4rWM+cinpqP9SdMs1otxi9oQi6/xPkbkHcj4tmUdaEH24oRj
wvi+VWts3+JotaVsna3Nw5dkKoZafgHd68Wm+5LSF7GjAtE3029/kh6wU9lHCVRAbQapkXhb4/uc
5gUu55D/MFFFL0gDIUVz6NnAoYsdB+rvnLDgMMhxDX1O6wmBvOEKi7JrRo/j3uWFvhXfPhFnSQsm
H4tUfAyYRHPUWJotVEl2MS51VMQYQKreYyQ+bd5CE1BbYJcRpIGY14lZXNSear4u0RQVgSWLmTbG
addFYSQuqg2KAN96ab1n+qZvZXAWOCkiW9UPlrvFn1G+lNuhKi3UyhZ+inaG3TFuHxKI+BRQFzWR
kAznzsjCJxzXDhVq4kKPomMXUkGwhY+NjNAeOSYqUrYZ7MEX8I0RNnTt9QEM8Cmx6taoF7sarDB/
Ezhmk6vTH0yxTmZDWfCI/dlPjPiGLft99PYfqujiQ+sVUO+Tpk/7pCTDiIAXT+/veAG1997RdeFG
xqfliaWM03ywV/tCwBY0q8s7LV7mOgZPLc7j0RKeZ4vtoLMQIAEqmpmtVhCtTpsPmXYSthup/1GC
B8KdC56wPufrNb4SP3RGG74KEgrgnXs1jKkNy3DIOtHeRAoL2f1YzRpFKjiKCnAfa4DxC3zVlIfM
frhhyJ9jVYjo3kLYhzwS17dXy4tTMvTnilCRx2PekcltkQ5ggN/fjH+iLhsB6z7EIToLuHKoZYhK
Y6tNpkqc5HYf0Zbcs0R6dUwEPO9tNSJIuwGa95aPino+uZwKNBYJfG4mNKAMwfv62FjhBcOIhWBE
/vs7Wavnw+85Xekl72bdhjUqParK7ufR5kaWUCM2F6WAxiKeEqJQHGX/fa2kCFSrx3MQG/mtG3Vy
DPUqWPq/KWJEp/4nj+jqlIN/2VFqkofVaSZG4zD1Dk0TD8RLtQ4us2323ssjrZMumnY3OBagNyqd
tcKDn4IVmPBNE9NKkAg/Dxd0rycPmFXlZJcez4HAjOoRnGr8cL0FZNrDGTbAhfxo8B0xtl0OmDmf
ndsnIqelKr2jd2PpKrm1+w/70DlVp64Ay8nrU3mZ+krmkZryaVtisMJkN/0c7MxfO+q5GX0VNpaW
9WrJED53SXRs187dwCpsON5ISi+heY4QliXb2iXvLdiMIYMV6/DtbnTdJ+hY4UIhjCQ3k/fxOI1q
CbuJvfBmw4OF4YLYAPDkw9WeL4oEnT2pdWAX2RSNDeuEIYC53DPVoSjLFBwmngI+yJXl0j04eXM9
LGg/eHwsoOGipc2Fn5H6ilbms2Iog6OK0gZ+RhIRxaiKLJky3eS0LzeKkUeR7qiNhybs5nj6phEJ
qVZtGsRKUJYlCSA5IbRj3++ofKdykyUghpfrHJQ9rlzcfLV29wiZjjhT99dhJfWNYmrO7uClyovA
rF9I5aXNB3qoNmcXmIZN3cYoZHHdvAP7oZfn3GzIJ8Mgt9ou5Ob/uy9hz5IPpRh1sXMa/8b38ilj
eC63VSDvYRIgCfygMzejj5rORmUgfjS+jG0yAIgGzdU+0dFPtTMdaVvSBdwWLS22IFfSaVlc7sMq
WA1r2Hi21dPavQbkFCMi9+KrKWcQWTOLivwZIHta3MOD4dPNemid+JJMHeNdCEYPzuSZHwsMU/uH
g/GQWFKcyEeaQB3rcx0CfO+VltfamlpopgqypbLHbPrHwRANemau7tlBaEa0DJ/ibWFo+pD9VmdI
YEQZWFnN3m9EaikCTlKSu37vb5r+X8VU3WfKqEyDHnjxnR9xJT1wcELZkuTSFteoRHRYaS169iNf
Vjipt6kEBtSaynKcpNIoeUErQLy4uZIOgPAUf6yiplVrkeyYWNaAVu5piZjuNuamF+cba8g3opjf
GovB7LYq++Qba7IUuauNRP/HlzBeOutiogJtueMOY50gGo7Z2GybzfdjVpGrweihvXPsrSRawjUZ
kVJgMY6ZH/4b431nDXeultCUHXPRcJqwoYJsqp0iqxAKTFvIpciW/Pv6wpAOwpIO60ZhHpVx6BhC
C90R8DyGBbNgh8xl6aLI9rx3uDvgmC0rw29psYVjMpwOBMyNZBjHYMdD+c42cz5wnOGcwmd8iK9o
SsT3BFAaLr4sLnu/dpQFGNg+fJwiaQHQQOzaGGlHo1kkf7YvRJ1ow5nQGVZspSqH6Q28bf5zZhP4
W2R/MAqAIFykvAX8wCArBTk7BaH7+rYnjkwApG+8lH3G/Lz9ohuGH//Ggtp0/Qbb642/LS9Npcse
teuxp7F3RoGVzF2BFfc0GWiHZzikml29onSnD1jYwSzSY2mJiQ58p9t5w61aobSP0+jyE7vRAv0D
D5tRGo7rrOmM3ypWhjQ75x0sqnRosqZ7G28ZhKrsoKqSv2ywtvaiMdxAxgAPqwyLBDlHTNrD33NH
Legwi4/qx/2XqC4xilDV5eOXQhM8kFPibEfUqHCdJ+n4ywWgrAJl+Ah+gBLiLygQaDrhzXRLyoUP
6pq3i7YEXJzbWtRflS09Ml72qztpV5YLnzuQaalQUFDVNSQCPFNN0sFUQQmgDjgaKg6ZUI7kXb9V
QQDSq0h5IAG1wQopfPsEHWojbSGAvCbhZL/vXe9oaP+nJATYUWMhFBFrBd0gfeYq/spiTLK/KEj1
Cp0Bjz8yj14lKikRlLXqBxSohqI9zKrT52qhBCjZHQZs3EEklYTH/dzN+Q0EpdeEQSTaZyviZeCv
6A/HskH2BHxx8ajVwIb85644KajEgHg8lVGFm2DLjRLX//sOENjcOddDANtthFwnigi6DzOZPyN1
BNYogFK86tCRGsx9mV+RABhkFoznfYwa89d3aeHXlVtMpGLNYMYmEor9Z8aRId9wjZXnylVbn4Kw
8G/lAafGLJsH3QGYjMupf2prpa+baE+S1LkwZ4A8XDWKiMUZlKyOwxNxS09k5Cro+BrUiZC2FijG
wJqMGo3yif6YW1/pRBTcx2Q34bQQOdgRtGHqacbHijPoNOTKFowavLlP6/4BTIzgFi8O1nKbBkKU
opJU5g8QGDfDrfVsqY1Go8zlWCf0PY0gKvrXDjHYjweDMA/TJXC0wdNF6pmExmCGmGeYg9F/nRt8
iAk6e8pHdM8GBg3eabs0C7h/o+/wOUzsVxQBAF4aO/j8uwjD/C0QV8IsRv/nT9Qg3CNCk+5rrpq2
vp7yu7uOIxpX4PHQWbRf+3S1F1reV8mucRA7jpxZrdke/VCkIqmLlI7DateS9pHHab1O1NNsztZZ
MjU+p71VeIzk0H+xgSw8S6ZOJEmIS8Hc0HuT5gdGv+Sb/2RdFHCUM12IcqOoi8tzvk/gIPUH+bDs
6J0eo7q64FibuknuFBm36LWdlU96YKBc+cnsL7DxGSJMHjmc2666E3FGOnzcLWqCPsscMOEy3hXe
5LK9AT0tVhJPGVXrzDS0d6wOw48cEnxaskcIZQrfvz4oMF4mfOGBkfzXcYvU74szetIkhtwVZD5W
XuoVC9PeC2mSCWeEd9vXbBgJPNWUkSdD4JZjow5TqVO0/JucXPfixymVExg4GRQKBGM/BV8wagGY
+qEPb+U5XidIgTj/VSa2HYpfoddiFA52JDgKbpul2gWd5ucXruV7TyvLE2kCwpLsUYV87CH6PAym
kI5xYSbmzQIZ6iZiLspy+usXZJC0+WhHVMxA5dPxjdnl9Nt37Ec+jY/1mxTq29LGxmj2em+KYkX1
jJxozzyJQHL+HuuRQ0YFDbMx/KoGkKdGPIoul+mBTXkqvUzTnpENr9sU+ULzqfcaxKuE19HWnZ/L
STIK1IUfA248ey05lMG45T1cUzlfjTuzK4NPdZ+JqqL7kFNOZNPnb8Bzu4oebjVg3BsI0ktHUUEy
fjsNF+qk2kAGLd3mrtXd+HJiqF4wbOUQZlO74ocxIpq7mcuZBMwgGVEChbvusFsuX4nBs4TFNShs
VEFj3bbw9dQtyhz2+w4nucHWoP3WKyc3kzpLLUEGzD/HVDmcJbiJWaShbIYxXLyNR9kXd7pMPU9q
QpwF28owUd/RZcIsZvXN3rmgmuHcygkKTyTsBjQ/LCtbrEKZyzGT3IQ/Mk7lbksEkkwwR0UoUB4P
d6/B+tZ6/QupbJ4QAqci1JADRgH+Dzf/S34wX9WDKM/0GBA3om+RiB5fvE50X/se2YWHtl1pfgec
SUyXoEICw3k+Dl9OnfzDd8bP64v8gc2CrVrhkSa+6FtWCXRN44RiGg/47c5GMsCURiiqD5nTe1KQ
2BDaqqva3u2xrptU9MvJ275auR5NH5EcAjdDhCn6bwIFb4gWRqAYwDVs5zuCOHQ0i2H5SOzW66vU
D7uo9Sk8aQBgyMxSztgoVAPSwCPnMLC6aCiZsGRjh8l/Aq4K883M+jiaalbztYhfH2wQYEqCsDly
SbIme8b7oH+trddxMxWc5yKJdxMi63FY5gRNZohoNNtpmdz6wSOqszZwpOgct0bUE/AhwsFdWCwG
hsQlyo652RNJaGep93rc/3iL0AroqXJEiYq3DiD1EcT3vbpL8WBYF77ZcuDdQsN8Vy8M92BJ/T58
M3p4xKEJCFzwIE4gADY7MhEZ7h4MJhho67g1xRxOx5RPJi9Gv03b837EJwXbVqgI/xMVv0n6o7o3
eKLFnYXlKrp+1xpOwkJJYRMc8gLBnP43RsIL7p8DxZsZigriJY018s7jN1GdZ1WdJF6lom2NFPQQ
eB7DJjzw7Gm1HD2TiGQkMkBeQTbnLMzL+qx2lDsx8h54pXbFVCnIfWhSzE1b46WQGk+k2GxBfouW
dNFSjibOEU+Zodfo1rzAxuhfIywlvN9aAJyyU/IDg3gIEdXcSlGRUbPPgfqSX4Yb3Z4T1UGJjLzb
K5JfTTQmplEiBYE4EuAew7atm2EYTcCBIUga5BunHU1xWHksPUV+4kC9U8fYRBjWrwuawBSZgiN1
iSk5cgaN+SltQ6MKg5+zUrZIywxL57noRtBXPswD1O4pyv+33kxMRZEL4gE7kH93q2YOMmZV1nXX
j8yG/NrsFS6zUB13Rf2gMKsZPANsWCNK5Z4y5JbPIOMLsTAbfNpYASrIE0oAUnM7Jezzeviu8/tV
BY+1U9FQk3+9SwCkIQ8MM0F2z+/oPLwBQ60Wug4WPQQH0Ao55pOn62MAITXuuDQF4nl6tPa6jSSw
BVGfftGcW5/+bvKxMlW3A8AAlHQPm2fWsWFLHt1FEQL36kwS4viveJ9vkcrrygAV3s5ADgrFZC+4
EKTMFnOIe6z/tsdd8gRXmoutkXpBjWzKsdJQ7XguIGIrUAXfSWvgDnNFCmRpSXVcMuv3A/FlF15u
jW/lZWJKjK+7GtzHM74x+hz8g0qXfvmFUyTofSHLKE5fqGQhg6x87JlSU+G1de9kVlWyEU8s+jsg
wrR6Hor1g9Y2LYg5hTUs5Ufe65yENWNGAWoib2/gO32XXEtdb8lqkpTxGSkYrDKIr0cVMt6zBR17
7Bu0b7OJYxMZcwhK/b5cgJVnFSDGsyE8H3DSXl9Ab+1YuXQogCM6kk+pHwKmxqMbAo39PxNzvioz
su2+obyj1cFxEHmQkSmHDm0LqRt88FisPuPVG0dOAIlgGq0qhQ3u/7AEsH2oKFq+L5MFjnAcqs2R
HDkDgpJk+7RXXxSx3RZr7/9mibmdAw4Z3kl/p6dAglej2+kgIDpntlayaZR/Uyn203Q1xUOQNzEp
eyv4v8sR8RTovJal3e26qXOCP9X8Wd1UlT9h5h3LB7rKhO7SQ8RSat/OoMxRf+izFUrh+lwARU8A
WS6QwXk8kANRrk9ufzxx2hRsBX63HNIkFpbv+2zKpQ41PAJErAmIRlV+E0uJeJ41skdygehT57Tl
XeL1L+CI30JlBlvbTN/bdZUePNaUqqU+WPByTKObxtnHv8v2PYUYWefAIxDz5okGRupSDt7O1R4n
TH1rW0KUEwIY1INmy5mVgY99iceFDjvZQ72+eZcdKeDew1cXzG6voKkcMhK7bIs8swH4Ob+i9L7L
X7gJTOzuR0n2nZ645rA6jn4Mmp2VZYDbibPHI9WC1jJ1G+PaN85dme/XgvxQnWNy0Lg0yPnxZ/H4
iUmp9CHA6uQnUrZQgml4m+/kpcbd9fI7W4KimBle+hrYgCM9Vw3HIR93YBIagei2ihVZ8x0hVH78
MLgFaMp9p6bWsWW5kjiVOsVq2YYWMOIs3h9J0AX1V3gfX1Nvl0fCT7tLc1XqMwWJAgLDq/qsvFZ6
YgFibiBfB9KAGu9uDxfH5trZ6uTZa+fkv1Tg6ec/wE180h2PrfMNS26Rjnt8Qu3GFF3obZYotj7e
+yHtyE15rPbmsqJDN1GKnx/JKgXItPIV0oHcuaKPHnYTD8u1UXwwdnX1JAeq4LcLRZ0hve2sWMTW
Cy7/z8vDnltGou+tigIjkX/5zXhozsg3ELBBb1H1GY0VpKOhv6fiRE0Fjk4s3YxPcJSIkY7hThoe
hyqRPSJxMxgwXwwauzC8Og/qScDJy+qvslM/fTVofxXZ8kWX5mlgcvcvVEymzSU7DUg4pglh+CTU
z0iAF0s2xGDWFiZ/h00Wfj2aQ7CoIw4k5MEXbm7y+oaPkKyfHgiToTaue8BWC1sSB2yN89FGhm5V
vJMUh5kNuL/eDpXEwYQ/4KWXzjK+KfVqTmqjY1TIH/Iwdqemj1HkLZt/Vk6Fhj7rOxdDKl1Jeguq
1YoxOKjuP/G+rtBM+yOzVWS1GkTry8rYr9BxVE3xpj2G3sBxdMaGx3dzpIbB80iM2+sdwsaaQz6v
3oTB9tmzjeTn08/y/k8iZKnyBk3k0UfCtx1jhgt3sWet5afydbfo2K2XC7qAJedYrxQCQnY/WPsS
4h2/lNQVBiVwCP6xDuH/QwMtd2DSopuOp9gIAw38m4lFgUBB2zUgXE24nZYCxXj6Bk2P279PkZsp
qOACT1Cakg2qWzlMDN9kofWsSgVvcLiecqNNwvzsxuLA0GahJTK9f3WRWxir4e7f4q8k7knShtUw
o7Jc2Cj8lPF8kmzpowNISJ+HvaHAnDWBT07Up2ZSSmvZFCBqnUCRXQ7tovz+Xvc4TH54Zs2jmLcY
waDYL/i8QW/tbMfhmhBjpukKcYLK72GpA/PDltifxwwj6YGNg98k6sRyEQdrCkaLQQaom3WkE7nO
OrK4HhPrnLmgnq4NfSHs5WfWSQK7Ddj2rwApnSPIfF9L1z1f2fdC+MFmMOm9JcdG5IS5J7cMMxVT
UtvHCebLPPRAoVstW4Jm6fNnBZM738JNyDeMc9OvErruRdhT+bkWitd44GWj4mUK4TbPvZ8ElntU
LHs5vzCZAKASuhW/4Q+VUVX1EmrkhLkTnMcOjX1XwXb2wNdvc5PsY+jGYPlwuORcQ3ZTSQsygWzW
ZQK+6L2sYSdfN/C8NhrcZJDsKvJsC8t6j/HeQskO4XGOcwlPeYVn/vIVCAx5tPZxfH5Bz++qfKm+
1WLnyoL0/4Yqz8V79qgX6VxS08mKaPkxcAnb7EM7OuR7EUkTQ3fr8tQ+C3aIXxed90qMiEP6bCC2
loweRBovzVw+r/PScZN+sG3E070qoDv0GvdLHagOt97fFxPFa9Mug6qDhDqkfE5WmYrQNzbWThrC
Rh6iCWHxDQeIohTkgjx37LO6aC86lfcAjfLE+DSXLSBQJRfx6NAU601uKCizftil2HUkTWNg8fCy
KqFX9tn4HNH/c0+xog9J6s0PLCpHyuc0NRGa6uGGBHWY4ctJAr3aZlOCarVGjTjYgjNoH9dtspNA
vt3pMSWq63t22TlP69kpJ6368aVr/DEDVkR02hDDPUcOAAzy/ttzKG4NpTdpRbq/VGCCFg+FH8jv
DlNVLdTLuDBpPR5VMc0A669560ioWmx8YOgZtrtgGWtaB2vPnmUUW8dRl66DHmisqTApmmaPbi4e
GueTlmdW/Hs99nXhRJ0bsVQGV+c70W0FNSyzDNzbbv3oGti/YJXx/dKZBPI0uJOJIrGGuAqqnbMQ
bozuqz7I8c/sQYT1EmWzxtT8qVNr/HK3/sFu0c9CA/9rUk9a+FL1qGcnPPUeRQuvyMS3Tx4xcHrK
pI6DOEaa3r2sPVn76tefgI9+11C2nd+yTANy3tlN8ydGCBqCUdHNRLZaE+F3moAG8mgA248UQSR2
tBEjMGuJQmFjD+tFzv5ofJs1jKecwE0ZRuG7PRo0ApgKw/bY7vknR9wgSkZnKVlXp6kgEgUkfVpq
S1DVzVMIt4rs9bwOGALXAL44N+s7lgwganpH8wQKPTwSyBD25EoQdavAxhYYYazUBJrDd/T4a5SB
fVnIXkQOLBDFlbeQGSPQXe9l9QSl9ORyBmFmYd3jOCilD3WzCqvRHvnDVfR+OgDt96E3bmRfwfm9
04DQjzK84tXSoZsAZNKPrIIxlIKk3L0WItdh2ZYwV0/4hkZwd3PpAwOACnezfJD/1m5V5gBc5EoN
hMY1gChRl1I072Wb0IorfYupJGW9Dh7j3RtBN9yIEtE2dMQF8WnVBMQSxoulG45Da5ViJ5gJ6Tvt
L/YAFPzMUS1sgM22WFEvsPiHeAawpeQ4wWSS/rj76mtk6BMToUpWAIfP+3Sef3cDj7VYB3dqZAPQ
Bj26kG2HoCctlsa1LYPGYYPut1Bmkv7d0yWLqCb9k42ZD+JqNqy9JJHKIMYqPwC3LnFA2GZ6PbT/
NNkBs36TPH+DMYm2RqppV9kmox9AyVQwmhdRDYSKgqEC1SwzTp875m0fzpaL8hlbOyDgUJHCTpBz
GsYwYMJxvhURFSwBMeDq8NAsQ1pP/jVlDZk86aoAqrKu2zqhYvd29ed1AbKhMJ5RH0WxxZGc5Bly
x9R18hgwShx+9nirgn+salkJZf4NHYDKLUuDnWnfGOjlsoaQkB9/x/SOUxsaezgZw/noFaUYzGfU
Cd9cq2kwOf21KCHOgYfPF82Rjcve0F5ZiQZkQCgLt9M3O8SClVNGKg3rk2kcsWBBYJ9uDUBozC1q
kSCtpvgHnOPSjETHsnWnfjJVcuwyn27W/+ekrGuMtK1GcHnHUcr6YMTonK9eNoIBam8zBJU8dTiC
BJ0sKRNzaomWHSlZGklqqaCIlnc9uddxclkBBMO6E7vqWjzVeeEiKovs0LzVvd2HQJKyv52oVm0w
NvbratCrJELNmXjum0+n/M5PHd567gDWqQmfX+8/ugjZqQ3Smzr2l5EtoA/3ziH9mCcvsqLVaskI
U9e24/K0xID6EQQBoSwSOmRvZOVYKXwqA0hdlb9hhEyk7HK27ZhWkm8E/SKKQAIONlU73aEEl3l4
ysHNPnW6KNIHAbbNxvs3IA+f/WaCx1R+GklQQAT37omkp57jE0XM3qaqTvJ38Ts7tr+/2LV6T80w
508Qe/0Ty6u2TMlFYGAvb7PT0IMGJEumLz5KlDwHWvjtLk3Om8wPbFE312aN0blL4EPwItHnYIuO
US5cgL4rOHaX44tzzTDl8lWzjNcrJpbrS1Jz9fqQhIFvm+0GpMHWmyeohE/fWVdFeJNUoYRGGyTl
uh8xciu2uyYZPFcgYqe03LIclkKfeyi6rFmv3SeDwXlyoEGtz91r+foR6LLipAJ6nLe8F3DMD39Y
bBfjbBJ6SoXCfjH2eHQMtKFvS0E9VGcmZQjvFbeo5v26okZHhTJwaRmVf/r02ZcSrnM2srmR5f0X
+TiPjdm6CpHc3d23hR1l9YSKiNGNYdWY0AxrDhLFYICa7QYGekXFTwsEwPNYFxpiI4+QRRhniVol
jnxX2JXcMhYeCS0SiVlqrFpQ+jHjOmsgycS8ox3kVrILNr3Z/r+SeJ+d0wDOf2ZKDOLolhzeGEaM
r8AzeTAvAVjSKsToLl72aWX0eOxuQoD5dkv/zjkA2BcgCwnW5rIStlpcOkSJKoJfG/YnV6iQQKYa
O+RDKD5yor583qjyAVSNNQylm9tYBUJQKxEfHWYzfc/TPWMXc6VlGbE7ySqresCHwNGMdkO8I/np
nxTw3mtgWmDkG5ZhtAEGJwgs6Qf9jYDLvvHhkz6cqlhLgVOZoT3A3NhcRa3KiqqtGA8/N/7sruhS
9kVy0Kvb1v8rIVjeI75UPKyAe/At+n62pxADFCrNONKrNqtwnrKKk8yJpJf0XZGtC/fW8vt3qISj
GTdK6RVaroC/WTWcSaxOhM7DdaHBccUHhcrTQ5gWk26mj4u9LitRZ1/iMYdXbLS/L78Ftkaj4Zbd
4DLXGV8WK1OK5S+FvJclf+f++hN9OTsh+MCmKi72Y6Mz5v5A+YXIn0c+IqfBGZHd4yngfLn85Cym
Bf3FUzcx5CSs4T35uOEOzHcILwXbTe/wXFeH5C5RzwFlc2moxgU5NY72kA/4O2p4Pf/q/OsSC/Eg
zt8vZ5//95JaimMoJW9XEye3ZwduuHOn9we9ym390NBsLEB7KAerHuOUGimZcgfx6QzUf+GZFKX2
c/Wk95qOldmq8aRDxt7HH4CGIHsTU3tdI18C7TvTLvAb2fNXy9I4LDxcelwoLr3mHfLy08EvHqYS
f3oR7BG3iT5f2k0hWZjc3efP4q5bWHlJ4k8xAgc7emv7j990nPx4LLXHKC2Mu65pNlcQnj4wYlcb
K1v8FwcH/xfuHJbTg1qMT3ykOf2z9/KYarfByS1PxjvVfmFzcAJ8WcFFnnW1PaAJXOkOnPfBYAjK
sdiHtMVf4e4bZ6EXsUwToKLmkHI+mmEWuGuEGhwVi6JmhSwuoHDyF6GN5HGsQ2SbbliFSga5/9Ix
JH9I1U/vaS7opwAqOVAEV7U2cVIwNjF7C5XCS3hbYen5aJyXnQp87sLb6TmN1AQn0Que+mL1OSkX
OIRVZzy7TweSVTSoDBLdxtUWX7JEi14HhU54RXEowm//FxucBqPLiYbCgna+3Px2x7FCRMdSZppE
eo20NGGWtRB20icQ1jrecfQojt96kXJxlVXbzDIEAZcTES6OmCW7j3GrJ0Blij1qUPtWc93Ltl+U
ZwxIVhfd6C9Z3o+ma/emmbGsfhMIyY/OuXH3Y3dPSMCrWEpaTK+N0Sw3eL4dtH4dy+HzB8ryF/E/
75BzGJ9acInVWR73z2G05hmpZo4RngNraSpZksdV2JYjIYr8rS7yiGEzLP7CBXMgvy0xWYvev+z/
RscGdTzPqVam4V8zbOQZs6lfUSbP3W7JIeAnEDBbONAJeikNCmWMQMnyadrX1pxlveR0L5eEwE1F
LczKPs3h5VgsJ9KOxG6E/bcNeLU1FJcsRAJo8DfiQa5SOG6eyXgifYIHCG0qgow2c9i7stUt9biE
bIyQcvk2848e/i9WI+XaadgbHrRI6bBc9vOhlCgj/d2IcAkLOLmgtZQH6UhpriALCsYSROralkMJ
IyfPb5rlFWKQFoez2XjCZr22KchQKZBiuhr6BPyDOa+sWqAmvk+8ZEqVHYoSJigUegudqH40ig7W
40DG5sp/9EVHHAmaTp9Zb5jyKGPLyx45KAzCT8VZP4zaLYt+EzI2rqY2AoSjjUgGFfPHwg0eefPn
B9IwjFkigE8+5D5a2eUzYh1kJfW6mPbiEC6QEVvXxE4LlFWYmLZGizje9yqOKy94coIH4GwbH1QX
ur5zpaTV2lmo5a+oRWDhqj9sRowDxVTopzoEPQnpDakaRGh4POY/Gy9kxo7Aftf/YoxXGWP/Z07V
VJCuPUayDpgBRBqrYRrJGycae7mZIdDdT2pnQ/WVsWNJAmsImb+/YOYKiyA0oe2akIODhMlBKd+h
mXihh9vtLCZctTr1XBoN8VFQYz6nQdJB6wigiwqsE54BDuMbQAs1kgmtWNpHoPMbx0vX1HJ57KO9
KZqqeYAkPdH/HOeXnrvI/VvCjCLp1t4AuAIJPEOaqCUoWwSl81V93+fXqKxl6rQFjzYVq6DsqGoR
aomv4rIEgSaRPx0mBAmGAD4CGIyZOhPo/RwL9+KgwQHL6YWVYFLV8gEVG31x9pZlLlZ3kcz2SgzX
ETPNQBdiYJGvs9C9zcCVzVIlyNKPv9+3PADsuwumlx9RBJvDhPdSPItwNDaevyxS5PRhxCQiJAzb
NO2xOkmh4CCzcChmIhrraXEn+vnHOhGoimXzcbs2JWpmpGc3zinpOO5vA7rIMHqoDlxPcpVKHzSr
yC13A3yvGtJljZM/3VnefIF55hv5QtuYf6rT83ALXZnUD2g0zx/4K0BUhJp0dFp4y8WCHW+EMPuI
tKI82ufzT8B6M+1LcvHEu905RsTRFueEeA4ifjmqj7+7bWVU1W2t5bQhmc4tt27t7jffmkc08is/
7slEmcqJ/AR/zrre3gVwLGzkotoNFBbEvVNDc8ulUNA+hZHPuBSgTdco6C0N7pUbhAsp2dD3Ll43
CZH8DbdRdsNVtDAcbk+DtTJH1MOkFrazbjAipFrXOBvkW9FZNaptSiLp9+KWZ+Wgaph7PjcfYXoC
vs7pQhMcb+VrzfW4wE/c7k4UP/fXn9+9XhdEbZRqsyuYt9WzHn+P5ecSUEKXwa418c8SLQqxmg4f
/E3pfwe8X7DO/b/nGJKVCpq9ZfPnjCmxLYXKpEBODB2v3OsddxNNYPy9tBXVYFPI36/kguFT4n8A
Iz34UgCz28cxr6nB+5MvxbGvy1ewLkGF24ICsIrnxXdJeInQBCKE6YzXfb01TByig6/GKfE7gUcs
5YrxmrP0vj8VQlcs749/SY2QBEcNAl/NnhSYOKDVHg5cB/HdAQMaF+Q0ozfG/SJL5KMe11ghB93a
wxCN9P18bJI6HUcynoKh3HSdonXDfGeKHO6LllxaJJeAYndF4vyZdmjr2RxOHhh/bKBl675/kYF2
65XdQ6KE7Vhu4HxeBGTrqp26ZdM4+AQmidY8wU37FGQHQ81f0eK4geZvhx+lCSTw1xT8Tr3CH6v7
JQzPYBnNWANTDZ3/0nXgxObPTjPWL/6W8lNzMTtfb+2SRNjM5ivhPPf3dAVkatQoT5TSJirNlcJS
MSca2/1ovLwRieZK+UmZj4QuyjI9kn4qyxaAlkL6YF9Vg0KoQe1RWIEC4vHBd5YgFIs95mFURsrh
FRaWG/f6oRRGKgZJhQPfvIgbUA9+inXsA8kPAJv/nphVyzYoZLtLf8b4DVOO7DwLPNHsvL7pb2Ra
tSLB/P01uxRkfJRJI5rDNlrMyYSWmo4tYoh2jz6Y0je+YbtlUf9mjcEZ1RWlJ8AB7DYFLDQyRpfV
RsTuSj6gnhbPgwC1sbZmmO17BxfrTHJw8XoV1Tkv+DawLYlzDbD1OyJ0/XpAFS8cncfV1Jrd2N7t
cMhKhhjTmbMxfwCtmVuEoOn1vzviwwXb1/JJxnsywS/ElYTH16Dq7r6Ks3/KPMqa6B/6oj5yOBpY
YVgnth39gon2v1u70+BdgGBN2sEwKKmmmp0e4cCOeCeRLDuqaf1O4Vg8NlX6rnlpaoaonrdFX9wf
3ZklIGFizkVn/dub3yVzoWEOfc89EEk6+5DLDqrQoAglmLaWDwNnxPmcco8spSACBs8R9gN52WkE
+GPFHDo6dPYKIC+zVU+lZpleKETXowSuX9b6F4CJzC2nXFT28XQ5zGIc1qYBf39lxV5qARlymP9D
s3MeDKqVUapc2bL3prcPnhR+89c28gik9/zrGwbrj0rKkLwhqV85vuTkyQNnfEZ7YCr4lKHzbYwE
gxGb5mhgs96eC7SR2nwR73cDd1imMKbqiy6ZeKkcU/3/s35jE+mO/r6DjEf/Y6tfCulwjIYzWxaT
l84zxHvyoxeEZNvCWezB+Xj8jsBPKOjqy6HVss5wTnxR1QFr4gNutj3/2oCleIN+NWXGn5PkIN1S
Y+hgVo1IuTCUhr+l79DHEDPjQEnU5H+izab5vzjeXjv3j0sn/J70Wdf9njtFuy5avA2nDGb2fUs9
VJXNjOTrdAjM0N8EEh7jzXsKOsX7Uv5G/mHjB3SNcVQrBugaaVo0m22uQQHcDznmdQrQ4YHaI2by
CTI0hldV7e+gZ/2oPVB8Hgp9KeHe9+Dy5vudVBnHk93lZ1CGznsPkoKrvGadFfX2isk/4gifqrf5
M2a73gT5g32WNtyeO28LR1z4HvjaoUWQjN5ruMY6IpOuKljg+varBgiTwTRmJ4BtWto5go9fyi9d
Gt+yv8bsrEA3NPwMo6z7iW2ickCGQeNE568iNwW3mmkN4rzzuPI9WKn8yYVW9DGC7vsHaMfgOSdV
MNZEueNjSZUN7spBXrfOwFlTfSTbRRvTQ0sPPQTJp8rGmES5eZnapAv/nW3fFaDSmA1rx4p7N0bq
7C2ZzMGyXvOHDVqLkx8eN1V69xCvwNm7JaK6POdvgGOGK4LtXsBEcaAmrIoAyI8sUDDmN9lTUOCx
Vnh5Xg362k/Uk7oKSoKYc1Xuo6xQ393qxBHgTRG6VFQAk+KPq0h7N+X59wgzhlZdpxtFvO1uq9La
f5YBN1cSiUmWD/1KeDuOk1xvUxeI/9Zs/YTM7FiMNWW9wOwiyu27iFUNHMTcymAxKsxP/FGvYCSo
r69b7QgEKDm0CFFswW4ezbWXr41Xug94SSPabdD82i298NgKj6UsAJgmjsjtvUmwQIyuvRxY/TtG
PoR6sRA50lFs2qdkESuo2dKit/v89aQDvAQUOeFqAZkrKzbJxrokuSScvnqpPpWGz442QPLzynm+
+NZbxV69FMDkPOofpgcrut6l8oDkDnmoRirO6e0i/6jGN86nl9/kRwUEFCiO0zVmc4muR0u39K/u
BoXq/eaWv86IPfXmTmjS+2rD1uo8fKqyepWkjdUu/36S+wuvxIa/3+ARXcL2wHVTYdgVps2psrkA
zap4Boy0NDYSB87EYbfwKT5KSeqsneIFbvqDcW3f3hDMNKig5fk2o7zRtxl73WWcBEQ1nkTZSYLb
34pqBtJyAzIJfv9d00WIyBALtrYLcwCXnK2TnFt5SSar8XDi0BNmQbaN7Uebfm3e93SLFoDhAq7y
EXpj4XQmL/CzMKXzL0yvw6uxSbBZscPyfSdA5S9hLqEI16VoTHt8S/pn5KQ1gYzj31+xALoCOyY1
qDsVEoPRWu9T/+/FRTds7YCV+2FV9k6Y0XsvIC8ScCRd1hMULOodGs6OvoWnX6a3svt6v5PuWkJ6
h4+cEL2CsqNrgoUgsxbf5Zg0ZYK4BINafORtB6gCt9pVSlps8wjBriAso2buRJz9bCG2nEn2VcyD
BqqerzkvgqhOf+5DCTdjSgThq7Cw8d2P5/wu2M/m3P3gDjJ3Gr8LyH3JdjG6ODaW0+NfhsxBTalj
zObobPkkxDWK7C5VboDwM1wy/cAHdpmeDi+EznnwZ+aH8sbcyfsd24bgpamMzYWt8lYW1ngg2Yyq
AX6nKaKj8Iv7SKvqrN2AAOXbkZfGEvXwMj5ayZ342pQKRlFCGOATNybCItY5UJ4yqvjhTA2yqxS8
4OEqaMdU5DMw8KOtCgpiYulZpzbyAqMOwAv+fFzf35NKhd78APB+XZrsEGPrNpenABdWvSWTA4iy
klrI24Kom3rfMskFdYj6JVsdOVSTUHi9WmgWYu1wBmfJ03KKN07U6iylnpdXwf1gRIVb3l3NoMpf
mmRrNEbwHi8v4CxxPGSl+iC1Rm7eNxQrgS86iEgNleM2Lv7dL1FEDigK+z0M7paT3/pKjqspktKm
ctjPT3cioG4+9mrb9/CcDzODe38H5fEnsklMDxfOpr97TVk9BjYoN9YffBrZAwi8dAG6YJewIOiO
U0p7P6xc9JExwTq9FS8DIe6St9/T3fXXygk5KkKRFKI0EPQkLAH5LfspMq3eH/Fi1gN0cUdznF3l
no9mWuX6rZ6Sb3/kxEUTYE7dzn32+L1NAoNPHO+KTI1gGjT1w2UX0ptZu6MOgWdXrqrLqNLFi4tl
KKhkClGaEffVFw0JMAdJQbhF5FJrHa52Y8yWxpWrNV6+3Me+eK+PFoysWaA991kSM+F0yxhDtYDD
HDovILytK6UEzO/x6aO+A0D54GoyaJHVyuJiJPZt++x+AFqDknG+Fs66oAeRjuBGIsEzCjWOHSQ6
OhFfROxNV27HVGo3vRyuN/RrIam0iqt1ZLKznUVGaelPCPcjbDv3VAt5g0n/1McCXeg/jhWnCzXt
P62CpiFn8LIsmDhS+uM6IE+bYR85g6xbZ+D35xj4ksiopODb8UIWjeModQ25Ed8jfGXGqKs5qm0v
Zx/BIh0A/PVuubcbFL7IGL3HQPBGpqvi7StYqwkP7k6Y6LubN32rGbC9jf4rRwuFEYlXRzkQdgq4
QRsq9kYiZEPBOPlu3VcAXIidQqyCBrKUekAm3ohhpmqwiVOFx4JjSM8mrtv+SCQYTHuNR+bfL7ma
zDGUY7lfV3VfGDu7NnZkohUF/ArZiU5Rp2syN60jAFyNGXgUN0Chfj9CLaAleUf2NVFAwlMSHB3B
s+0YLqoDxzZHkVaGibIUKqOY9HakDcSz5RejVvT7wujAiayoqF4jomYjiH1kyB5NXTRizdh+MKog
1Eutv3J71E4x1GriUXKTMKqAY/K/M7dKMPMnEOZ3jLGMUNmFZBGEjoNH2umEItQPA2jIACmiz00c
SqcaHxD0ery3Xvth5KLX3VDy52P7AdIMUI51nf5mqD6wYX4S+dAd5klBvBqIpHAwItZx9ZEVSP+p
y2wvNyURZ0hnTPAOD9jEZPuVQuNmCRS5xxP/nRnd7dIDyYObGF9Dj/juBU/tTwtxSLl7CGpZVUJ/
u34TEa00RZellR5fSrlZhR9QyXv0LueSjoMiSN4Y/9kFS1zP2+58LiZtFUrTfwQHP5nXbSviE21M
HkXFmXmtCzIEQo7AyI+nMTNofmHyd0ZhpEaeawcHhaU6SFKPxaWY0N37lolJZUhDiaCKjl1Wep/+
i6ibY7XgK2dzyGVvyF7xlZykMYSlxaOEMgjPn4nzj6pMun1aEje85v2t+TqJS//M3cqjVQZi7K4z
tkXaROsHtnhkPN4ktlf+TgUQVzFtfGGZ16wKjydugduwu173+GIoJbTOKeVX+WkB6UJ5ALT9VO4u
iFZLGJNJCglBoCp5alXaUqBb9kgMijJURmb1G8BwDCDT4ltxm6j5AY7wWwXPIMXBTr9+NacjShO1
3osUt6FbyLdHeN39z9gVe1HebOnaIzGLBazqr74CqcBqlvF2GhGiQ//0oNiiv1TZuvFSaQh3aXhf
FVsl1do0Swrb/FrcqBupKBRGqR1QUoc+GdpFlXkDmGCu1Pt8yhX+YhwwK029VQ+SWxLRyXYAg5ld
YmWNyYceScx4Ft4trzLC+SboKEtHQJmbx/pxeqoNd/3tBFQa+FhHnpLhyXzlgajXoLbL005eTjc4
g3qHBiTv9BngoRV0Xyykny/7et6Pa1cL+gRskN9xB3JyTeA/2puL3uV44iCPvcwfYkx5E/t3lDa5
cuQbSVXlfocTp9Kp1r86iZPJFhJulTK4Kmk+XEK+1RUaYGnbOBZVFyD/vqNJxtnofNGrfPSs6LUQ
1FcGDchBG2twmDEHFrGF+mgHNcm36rGuvdGM/Ri/sGapAV20UIe9A1LF4CeKXd2uxar8Ut86KHRe
cdM4wLJFhuMEtgfvSsErG9l882hdVi7sClaZwKaAC+CZweDt1mjXU+33r2zRRj0OqmimFbRGzlub
ZBjFsizpVQNNWFvt11sn0/CscCn7/HYDFRkp38runhRiO04Q6iYpJx3rc45U3Q+00xG4lpPXZC3/
e9mOvX47P6RqPkYciqne6Mlge8I4rF3kRR2Qna3POW6i9GnHA0678Kd2XHbcp7/i8bjiOq5T7OXQ
Ru72qHFiEzJ8F32JEYgjJe9iEDZ9m6ed7iaxlp0aiHzV9emr2tieytspcoRFjuyunWBBwCGW51/6
Vse54R7GpLIU988NZ6n6Xh2tLNFvHz2nldrat5Tb1tH8mkbzjRS4zK/R6D34XjsXq9ZSgAMKqFVA
RtY5CEDaRuxBS7TgkVIMvZ3cQBwCYgGQAa5nppIE/kAO8U4IS3F2Ral63Wk8Zi/SofMugqvYfq9y
nQ1s5JfblPhv23y+QaGeyAfJ1/27N9E57Ky9sGPHGZ+5pTiY2tSS878FoO4n4Ov2XDy+eWdoPyZi
UL73PI7kJanm8batPw1azAZTNiluR/knlCbibCfjLSMdCeq7W03liKObNjb8AChyfp7AmtWS9Nqg
lG1C0Mk/3kbYwR1zZT05GmOHSlXm5i3LjZe7odpkPtvK8l1yZhEs5tBFuIiDP1ZHT4NGzOVBBGe/
WIzhCYbKpgXTxyjHQhGr88kAt7QKBUpCRq8vNgRw5v1Zu0EEvlSUxs0Bx5GH80MWpiZ50CFyBtml
gd0L0i/IezJ0kETZHh1odAdeoMMOW6ME8QHoSYUg7HVJDvM1I+n+SN+nb6EGtnyHyZywJBHvKA0p
TiopddfO9ufieYdaNGLCe//N81IvkdAWL99tU1foMfPSD+0AuAR8py7lJNvA4yhfFBO7CemkTRuv
kMCAgrJj99jkGvVvRxyx1OYurbVWzBMn5VCi5FGaImP3bm87gxYkgEaztr0U1wUxk0ihNVy9LzC5
Dvh3JnNp49rJ+STaHbI0gxlpZ+DK0glkzBzTpvp269nI5Q/eexPYQ0o8rktAfXa31S+TLntRDe8s
iLgE6MdCzP03xt769CX9x7aQChbkACr8XaKMU2dj4O3KLBFYndPXIQ6QcyQU0hVdlu3ZfP1lJl1n
apAcRCJP2Kl5Exbf4ePXNYgZl4w97rR1l5ehWyHl57lqfH9qqpy2j+SHPzNJ4ZuRe5yfu7MKQgKw
I8MxQ/uLcX9OAPfIDr3FimiuaZsy1s9u60SVvxbxnGJoqlGWuKFr80iV0sh7ERqsxSfjX96MgEGP
6ayZrw+bjGhOUWx7PbqbO3Q+awNyVu4J/pAjaUOtmR3bX8tcg9cVEe8R8CcUAV3/DdI7NhlRMg23
VSqlqzr1qrak+L7WY2461zXPk9f7NTor6W+YeNm7k2hL8Qy9Rr6TnX4ZN/v0n8UXnHcMUAL8hVdY
XyJQx25DG24g6PLrxG59H9XVVzwRsRvVkWlNczUKut4J9QChe4FFhwb0rXCWqqd4u94H8iK0TpLy
fsP16vFQyQUTq9zGQeA6fJrZRR7WXimUWKZ3gZmj7ApGqKxAsuAbUzJxEln1MY1QyKq/jc8iFW1k
U6EnRUo6TE7+53tjC/m6Tt7QU3NC+SmGhOxaRrSaQLetDpQMnoIW9ZuDiP/o9JlznvYNWMYtFNdo
MyY9cbWnoPAgMR5QxJLSo2jK14BUVBKor4g7KXVh+xa3QtZsDxdNzeWe0WpmeUGCSuQEmTUln1UL
ezDuOr5YSyIE/ETRB9Q7/baX+P149Oa1jNFtIpbqrg/j0/f/uOozqQ6Dh+DJRmvZ/rPBwoDnmHdL
EUO/vw4cxLD3zLpgNd7fCXnm+BC7/aCi51PfzX9F730JI5krDPIgiq5QzU1CYwY/RDuYPDyStXV8
EcrcF5KHCyDFHkUEIAkPVdN8AZ5iDCAZpIAAgKGBtElg8oeOqGPf1LrvMU+EFHGRX8JZfmG7e+v6
CgQEii1SzQWvMCM2OywdttwlFVHPVmcpO9HnkPECh96zNtacwfZYuEY+r6XHLZZYRFv1Fkm5jHdv
AN7u/9d5YRdfwNPR27o7y5K4yKWbakA/fkQSVLXh/Mwf5uPexh0ITxCYiPkfyFrhilkDOPuV48US
Ukx50hyr3Eh+RvqgL1UOLOrCae6h07SQCiRx+v1GGj6GulTd4X7SV2p73Flc+ZqflOSyoIBjjeNc
t1BOaQXfgYlJMCSDyqbCM58DAdhpMog3qqXYiDOysW4eNVhVogEFtmdoOeg4ZdqJ+jF8DFhwS3+g
KjRxx756/yfDsoFvz77cgrAqpv4ZEHRr09sBY1bGG67Ts4u8qXTIr/VuSd0TWZOVQCfVJDP5ozl4
61/ALrk5BQeeAVBwWXve/6xO0+8UVfpIVuxPI3k31tA4J4ZBcirZU2vW/VIlX5f363130xyip7cZ
D/oVvxaqM9Yp72EVOpLwWi8pD++p77f6fBPUJTZcbip5nwA/A4QGqcZoWq35src36eeZJqrOIitt
BOZlTznmSC92F8b7SbkkFgM5bpowrG3d8onmvN6pb2sDI7NsvCShkwWjV1Jbhvawh3m9fkMBXmUY
ljhH6UrmgEFLPnAuLhHSPVPwpyIlwZ9wtDXGu713ewrlmipKI5t13vQvff1nOsB2OMMbcX1HreaK
CFlDAD53ZxxS0400YDnvpupOgT2maNMIZysRuFibzIxu+0sk11ehKIOh1VofEZn5zKJ0XWTg5lFV
HBY3Z2msrRYC1Vt7bcxHK8yVK+RaHGWX308R6Vpamj+ratxTRrojKdTP5nGfwJsZHG2Y9DUnchGH
IroMzrlZ9ERdqreAycenbyCpvpyDGXV3mRiuOkPSc94TXl42iScg0vGKNddl8AD1CQA3HlyIrxmn
R0v7ZDlENy/yUu7cIB88RU9CJCQ9CPXNXfU70XSVCpzPsDmJHACIpG0Gt+gHvDHYSmvM5fMBYMm3
Mr+All5UO8DrVXRW3jVxfcG+fjrVW407SuVEKV4nJ293jZti6K6H1bRIKjq5+MW9lj1tO02/JhKF
41oL+Y4z2z+rDYtB2wAXzSMnJp35RlBK40u6Nq6lIPf+QdbOf/mMxO6gFY2Z108LKrOvyZmysIdA
lCRIOf32y0Q7+2UVc+UGTLiS9vDdhth5DxyRt5z/BcLkex/0oqycYDyHVtPg/Lba80Rw34K2Yepr
t4sIPKvlPkwLDVlhj3JduzRL7f8KColBoHRnCXVWFAKY6CwCK1xjlQa45cw3HksGzY5w9tyVm3Tw
SyV3SfSWeYnXgEObnP0lwM6KCYtxDhxJeAyIncYflt+TJQlK9ec2RqiVheHQPNOdTpGyjd6fXjTW
7Pw7HlBXtmAiIZMso2H9DC2KI/a7J5QSKzixmW2xkVMiHfYW9KHdBarKEMlGA0+xqtqNLAQGYMAk
+3JeW0GWqIDObFp6uD2UCCaiWmMsgIaVmXoQqrN04vHtNn+wstibzyDQsoC9vYymMqCeMihqR/A0
p+PziRt4nBfZFteswnz/TfGRoGMSNB87cmURORRMhsJ62ZEoCZt16Cgb6NEE6Q3SZEUgTS/RQkPh
aEv7kMKEu9sE9+qV4QAHJhfNh0TEmkQEMZbMb1ZnKLjfos7nDSBUaNjsgHpf4pUIeuOV1vFZyTkp
jR+aBHKdLZuktsHqvXLFUVmpa0N6tEsjbmZYTX60LOAIm4vX6a7jzP8qLVQ4YeOK63U+djv+65Wn
ldUJDNx/hoBxSWUpmk40UvPt/bBPhlu2t7s51uo/mnIJ5t65oq3f9m+O6G3YAIiqLFIvDVjkiCiS
nTg++KR6qDJI3jFkZ5GehYUGCkdu6W5LC4D2FZGV19tQz6u0XIRF1e7AR2ddIyP27gnxoKGUtfDM
enuA70YaWEpwyXn5yzoqSK6lJf+T2Q11EQinXGib3M6T6vBtQeZHaV3HpUtnjxOFdpP9O2CD6fpN
3Mnfk/x39NToUJRxiFcka5oxMiUpzAiyWGXftsXttwU9jnMI/Z5yw+VWRzQWy7YM1Ukww4ayurse
rQPGql4MRD1PkFRvaamR13cWN0rp2xqAvCFo1N7Nm8F4KPH3Y1cU/h+hUCDK00jUuMI4mA4HFQNM
/s4y+LMw9SAKzZPUvWCcSkuUljMGlWXHKdE3Fx+uO2Dheu6Qd4gNj5ZMGKPafuDOix1wGx1kStOw
p89SH1A5ahI99Nijd4mMSDncI6kPTtXN8Rt0G5iP2QAEv1/33nWpp2EjQNw6Ptxy8A6ALzPogfDA
PkAc8KB5zGkCfrCfRRqBkCrBYJ5ngtYX2Ay+NaiVw6pes8uiCHg86I+NAGY2ksFW83M679M+BLfH
OVkMCwsuWg50BbtzaEoTisKl4Yyuzk8cIMTAVG3ptBo1RBQp/ccp7nBYuR8AycyEIsrTtDYlLdKY
oHngvn6xXl+8PWmdttyWrUFJcj4cK5fheLH5eWD3DeO7QUB5HsFlbzvVIiA60mLTFnbEex/PsWPA
Gumi4jqYhMns7FwxdzILS/c3w57QWSqSMBofp2gOhtn6V68mr36HnVmoIJVtkVcX/BDRBuf9gV68
9k2WpU1fh1uxVM6DauwGBpKUCqAlw7xb2dLZo9NlKQpl/1eaOgaprbVcYz54SdC5zZ2WuABfO2Bn
OpyzeszpPSIz+bdKP5jvYh0hEkBlqSI09mW7nhdrmYHGk8pW08SckXtLUxLqP4HLvivRVssebU5Z
quryYqXxtDtX1kv+bAPN/Onvf7xMaut+Tm+ceMD8GNM10fKbFmjeLMq4YdTG+QJQt1SYzOXuqwZN
GaOhrdEj9Kn1s1wrgk0fafUSmw/Wdv/YxfCEKwiS6cinTwBP1KUAeTPIR+bcwZCjyGU56tAoGAKn
j2ZUjCvWK50Pjb/VHgTocN3ltRspRWr9Wi8KxpH4oEnU0cRakvlE9MYna4uvjCq2hMb7/srJR3Wc
s49ptaPK3gIFTwON7HVGQe+/TZMhtySL+GpbWQxzkCX3zlpiyRBJy8R/4SyMdN9QwdvEZlibau2C
nZO54pyO3eAxFKsRL/S64/kNn9yDorJH9VstRfi9QzTvo9qDCjXGcSzWWbDM+kHyUcEnRqxQ+s02
UwsLskmpOLA+zKXGMBJPGWApwywf4dFy2l1J9Ef1KEBPnjS8nN4/87QZPD8FXqP4xyR22MQVlV06
NUlIkbKqahw/h+ymFCrbUHSHsFJ6fqUKyhz12MfVJHhm5jR/qwCd1rLqF2c4dbcJOjm2oeU0lZMi
gwGZstFjvTdsts4cxYz53HtRtLk/lL21BIBI6tYSbUmooHVZaF/2wQwahzY7/KZxnvtBHIff66tH
tXcxKd/7y8qJoru5IyiL6eXX9fd0W1kCdG9seDJZbuK+/9srD4gK/suVq/80h8OIt3GBwBwca9nv
VoxiUDiMIW2SMCHEWs2aQ/W0DKgVJRWGFXhYI1/ZtFJw7cvPyQKi3EexeET9GlHv6MQEKYKj6uhT
nVrhUGpdm7SgWRkvYynobuvGhBS3xp3S0sHX1OykeiowWyLncO9IcdjWLq5/ukciv3l360FHcka6
Sn/6+40HgLSjIQlvMVYhA54FdeBSK6wFBGCg0KYIO6fDtupTHAQ/xSHmbZateqmh39geccbYB1Ta
fhPhbKvGr774yXkJW2vl4iydxdyvTro40iWvOwsLSlhGXCAA5nuvxjz/ZISEIzILb+pCfX7BKcgG
QMW8r7aBXFhG0yixwlDtQfYVsnm6+3zrsSIIN3r0FdFqj2aKN7ZqOLAAV2plIQz1K6MODhQ2E/s1
stSPFqBPmRtYIuXcNy/kXMc79BuRi09DwPd9KG3hOzC/yTlWim/VaPCGldcp/M2o8MtKig+mxyp9
O5X37AeobvLT61QGuljRMzO1e1BZm0uOhU0/xf689LzQuTUj3QHt6caXDDaWNm33Q390gAiuCyr6
R37254B2OXFJfcjK2Gx91Xtb6ExF5Lq4pKQd77Jjh8GsPXGKOGMMrw+Pn9HMIUrUGcitWBIKOQqH
B4cxsOkZzCLOf7LF4DhrIaFqfmXMyTyEp5syKd6m4aqQTQXAbA+K0HC40T3K9rANuO6MkjY0FYpE
d/ZeMoPkS+3daDAegXoiKBVSboV9iG+r9oypxJEz44J8q/7kJJNcQ+SSpJuaZqvkLo0l/6vv5kPz
hjN7VyuKjUoWuBA7Fd88xWuhMqzw3Du724O4nnnAZUY0qWSi/Ebp7ZUhnolKDzUb25ET3Rr8E1yD
E4YgaMcuuKuD4zvGFZz8NWldXRyy5ahVcm/tTdvUKmHawaaqXL2SXK3iDR5F/hwm4ob2NzvaZjxP
1XlW+LK/QHrvVOXM0UUgVB90jSnq7NeSSVvGIAxqHWTjNHQZPIhtvlPsJxjUJuoW3X8I388DnjL+
02gWDDa6f/4Q4nMNj/67ujpphDLX43ImrshxzB7MUHVFhhqrgwEdlAZVTtTe4Edi2Wl7Yi1BY4Fk
Trjk/Nu5abAsH7SLpo0COwym+iIh4WkbEcojN7jo8LjsPxNeAWbUNYMdGRkCmB4sR9w4YnzvWDAy
KtyvEM4F3aiUK0SJmtyjMVU279sR3pkaHteJ0cZvcGrLsV3XfuJjS7LIDE9HMkGTioYURwfp6+9q
DYKk3owiAbhzaA5tM1JZuvZhrggHhTpAHd02HAreaIxJm47WcWS0yG890GT3oIjA1Fe80nQlIDC2
xpzOyMKNpqz608mPiouwtM4OCn1FpsoDegUrMNlaRu2iZfdKZ+GbsJSZL2AjhkzasCy0xcg+ztmP
RzuB2zUYFjA/myBEzzR9r8Hx1ptgSaA/+Rk0pydGV9caOTsR5eQ6KV1dfapgibJRUqZ2c1VN0KA9
TE2QQzJH+WRA9CUcIVtgXHPlqaIGRuggTaxT99QZ0ds+c3aFj9vpUm3t+kyGT7+0Wj1sVXBhU0dI
3vqv14ImNM3Yuw76UqfJSidHyhgDhSWPd7LzO3i9+oTV2LCoikYX+MVMoBBJmmOlJNrvql6Rj6rS
/5JGhYrGb+CdBvqSwwTCSipI0k7hdlxODawGxFVE8r9ZSpV5pvUyaygFEj17Cdl/AABVTW7ff1G3
bemetMyDYPCNY6a8wvNunURXTUV/PkzCi5CIE0TbckjMFpzIERRBBMAwgDjaEG00PHpCcSD9NudA
gzVCFjZZf6C28G5eK9BrHEoPpNciAM5EPMEBZzIGLV/SflYs3CygzWsVYtyePp/6RZ4vLROxoLCk
3VerxXIZzMqNxLgLOc2pOGq4rv4L/WiJ1ot6x88iIZgde5SQ0tkLQlZUwSRgE7FRKKTvA8uYv970
65RkCzy3ULhR6z5PADp0qh92BR1AH1prqeVdYCCF5mU1qhiqtN5pyfu1YNXrCWmUY3Z1hRVohSQ2
B9LPpgXIs98vNK0uM4eAY+IWrRg9oiiAAE+OWz18Y7Ez0BKcYjhIgg/t8iFredUF/7FFF+kA8TxN
p5sKIOfo8L+Abkur8EgQowtTzmAkjWmtTamq9IrwUgGQ2wxoWseuZblGEv3DWVOVU0Ns5fxOk+PB
eqFApbbtX8s+5EC3N2h0upOufn97/Ao4suZ8G6atfd5EFDIzXu480cQfsybbWhTR9/SOUfrjn0MY
RvZwrCCSGuEuU1rSJKfR0rS3dF/Y3/+wHtQMF66ZhJyK95mQv08LQkeeAFK80tfxKvVWTbqn08r+
PfVhOrQFl3x8dhMbfrDrwwtUkr3AG0/BCX9Xfp1EY3KDlUzDagrex1tO0SvWGaMBGe2zKrfEO/hw
e9ucU8u5Zw/0SaxRPqlUrrBUx1JAFa0cyHgMowXq0JfUa5SRYYFwNMdtquGVMgqq+IOw6EErmLQA
kqqs8f7lNwiQsXRZMjFWoa1fWfqan7S8hixuiVt4XhdAXUceKPHNrXe7CgwKJdop3aEdTFFiMO+R
mes+VWw0r6YbpFG4+YWeVTIik/q3F/rCbQwenSqBRpjPjALVKi4mUE+2Dd+cp5RuaxnePRdMciV6
AZuaPFKekvm3sZqCdkrHJ+q9kcMqbezEvmgAwWItP87+jI7gaf2+Te9bdMlJPfDJLEgHG1DOfsse
hhgExRogsk4hOyxrr6gT1HOiCb1RojgcaE7eFktI8yC5toCCWmtgKF8iBRaX0vAlPjh59lYN3PXk
Z8ew5zxTP9J4tfemoz9mI5ORqbMoh88jrx2S157JgobMD6QnWEZ6ItfPetsnWz18cM3p4I58mzcj
d9WRqE0BDk5x5gpmPlWcmdzlyWe2H6L1cTl5CnpRezH80Tyfo0G+NpV03WwrkipuBGXUiGI9uk/T
t9KGWgVS9k4LtOeDS1JAOwYdhY0Jq7udJHGn6mjipj1Fm8mk9+Jsc8CTnjzt8vFlyU8yYr3xSwuV
/tNr8KzPIkQV7E2/rSJppF4eqApLVd3hGz2xS9IZ7Ja6/+zSvX9MalTBZxnuzrtzUIVIjO87Y8c1
9RqUDWRBGtaIH6cOuCeO7SLYmCO1Lce0RO+6dIXBi2Z5wJ6G+o/jqZ4kk72Ma7b6c9Vhcw1YrVnS
6xvw3Sn+3kTQ8L6g2Yfj789qG/owsHMf3PsErSy/LMD87MtRaJGrmlArXWv62Y7a6oUrcK3Ql7RE
Uwqg4ZxAQgb4ULAcDLJFa9SRUbS58bxUlRlLO8xWrE2Gd1N77cAI50fPs3mu9lCqpkQzJlOmRpH8
lPJP3EWkaGBxAF8ZEBD0KbjDL8LKOD1BOzS9l7xWhM10SwQqN4a9IrqUinoOsWMDtCCsNihw4/TO
+RQTc9t/hnQSClP5Tnv9FEuUHS0l03Z7W2grHv5mIYRrhKfXt5cPMTjSD+tXxHvbkj5D39F6+VWF
9ymWQE48gX8QzcK8I/fVjvId8x0VFS4R8thskehyWPNdvzhtTm8FDAvMOCjKBkaqKLlDODVB3j56
kquXhAFzC4UWYgi59K4LS2KCRRF9khcZi3tC/Zkpo/xe3Y2GeFj5Bhqa7RIWcYIOQm/aIW8CB9YJ
Vph4hi7o5eff/5kexkagXAKLsirJnYHikwx1kxTu/dnriP92x+zXD1hgtZuMbP3W9lGrf+wcYzRS
/ilvnY917EKrqt2h8qi7+FR7dlnliiPR3E3CHMB+UKW7LzyRI9yUcO42158bUcjMgHQGqocibP6s
TOzKQbHutuWjT55U81oZGHpRUsV2k5s6XYj749ja422wSxalDAnEbN7t5HFdCVMyE+GEo5IXUG94
SZjNFfo9O1eAdz16dJOJCF5fjjD8dUPmvAJUfdN+inVvZJXy2mg9ftSoxmv+yljmR/UCR+2TXvjy
qD77Nqz32kP+h9s3fOHRjEtjxfiGpJSz8WR+uP+8Ezt3EhBn3//lySZPDhgw7Oru29r+SMMmTYFF
O6gNFi15RUUXSFvvTxYz/FsUyEF402NokOsVYl1YOCuNbZ5/0U56sljqTbcZc5rZlPEPPqEnOEPC
IfS9fvxqCXQhKfE+vFZRgb/HHFkL3Poe2oRrdam9LXEFqzPE7M9kCnTvTdCqNJqmoLweOCoNUp4s
C1O58r1eYfMyxKFiR0Bt+kC900ejhYJ622y+FsKNS80IjnFr8N/UlWmGXsSWhyssQjg+3CBKs0I4
UA88f0TMgcerNScRceAUDgwJA266xpfc8lTYkRM0RMrh8LQXTFXEm9HS8tfOcrlh58ae5LTqRCa5
1/dzQLVjkYIi7TqnwiP7gxbWRx1M1MEhBOxwRk900INC0d8lcAk6wLF/w5e5JoLg91sWPMuXyNXF
3iPbYoTF4/TkeQGceM/d75sFNLRL+JkoVIMJc5SUgO2meHHvFW3t1rkpYEzPnKYxLHPomaIy13eX
xTKRa2zpNMoaZOZuGjSywpOY6cgFdAYTFBXZ8wWduusYKWGShlCtKPyD6HT8CFzHnI816l/fdJcZ
MrqqfXdqeqNY55nvf4bXDY6QAM69Im6qtrr5y/L7lI3SyDLIIMRvmrkKrSmPnss4qQhHd6U7CDLw
WQWftDN9eIqw8Ax18JYVXXWPI+K3fTalza3u7VQ+1TZAgNTekOh6hGVpv/VMs1DYBzR316x96Pj3
QD9XUDVni/yw4o3+RlT/ziT+T01J1m7hkTRg8PdUNMYREKjDM25WvxkwCjqxQbpFCCOIybPjVSa5
e/NKlY3OgDoflqyabZqDsb/iZTDBgsXuM0Z7YJv1/poyURf481sxRyfjfpqVCVCwYrbtxNdoP057
bZ5/exBV9W0+W1i6XiC/ftdAIyESgYJpXWcY8XvfuRz5QRhH/WA9M2DRoyy/xS7cToTmEod1fY+M
TI5eZdAO2zQOxpO/CBVUmI3LYRJiU2GKX4V8RS4gUvLm9mthREM+eP4bzqucwdsbqrRLAx2bQleA
sAo5KAkyhqYYMTthVXl7n0W6j2ybEuCE/0ajnrgzWzmPxi/BtfAUaWWiiub+Qv0ucz1HgnW9t3UH
Bdsmr3QPYK+0Wm/g7JCU3ygycJmGexu2TVG/x1q1StiwZxgPa/VcMd+IAUGblGtEGFvJb2WDyked
xBnqEF8UcfjiXHo8Am+lMpDCq2ngJ0FXlUsQXEzpccIXztWwZNYmlyKYfXzB4ZPysD2qp+LMtWgm
fAp2HCgJ92grLddWbCCgWTv6Gw4vnOxJTBywusFhg+CdORcg3u1gwMVEcprzbTZBklTX7vuaOLk/
ZAS5zyX5b+n0ik9/3HoyHj+YstViYjIUJRez3P9aYiRXjdoz8OwA0wJudEXWUkO4Fz2/Pa8ftjOb
iOkWHmf+onEnX+f7RELYlSGWzHnWSbMx3CHWFmWTnWQNA3I2nObTPPU7mAJOYILDPHEtkWyiTUMn
BE+3ofqrqNqFfEHSjNINzkIA3mRsumbn93GPAfIiKcJirzfu9A3QOBTJUPXHRHk30rCcieoeEaH5
i6LT/M92QO+dOoHG6DhUejRF5M4ZFrjrpBNEYnc2pXmiraK+qfit/KJGJizyF7whH6827HYnqweN
bUKTA2ufLFRl3EzfwwR3uHd2SB3vJSZFXqtbGdLoXO4raDt1NBPAsEwoJ5A84RxlTLBjCBJJDJkk
50fdRrg+JZPTcPjzkN2bVRToum8hP3j7V3c9xKPBt7eoz4K255bn1HtuyPqGY30F9U9ZqdNXU3x3
+BmDWK2RqDKL3ffKZXFw46CzUjw3Cm5BhyLTYiso8mboJRbPmDmtmPxPumPPiQgg3vWDlr/5RtZR
wt5d907suAY8ievYJAstM/Uhqodb4A5W/s1ynaef5wOimSxGp7B5tfp9eVi4+b8SwGiNOhy90Q+j
/9huJKoWKrnr2E7G5oKX1rnbxwyj4q7pQFX9KqpMQTEb6VAFyoVi32tAgJg9+r5bInTV3+Zyzq7v
YcvyCb+ntzXDRaXNTSeu6cbDBP33Hol/g4yHnPm+fsIC3AYw1ekyt5VEIu4lq3itjI8LRMdbDoLP
qvdSNDgOwHLO0aYyjGdvzDkeZM4xkVs2SVIlEZqQ2NmlcNmur/hq/NfOhxaIlOofUmBalkj3o5Dr
3uNabxS9YGyF6Yb7qADEJxluS2KFTbkD642VTezzH4TPlsYP1g2FRcmfxcGjDKVpbP2gkktAopJ6
L1+vmacvuxXGLT5DyOZwoYLA2DTqWmWRpQP4sNRjIbXHA8JqL9doMsXropPHJfufCifvcBH0Ry/d
YOy8uEOAPRNJzvgke/BqBbmcnDrOvPMW08DfjgDm8vgirmRkP0UKhrWX/Qzqj2m/okIX60DsNir/
JmbVMpE6bXtACUuYxH8xZEWWv0lG9dBJlsvhfmsMJvwDhd/lYtXkZAJlWxN4WhCuDaP7xUMU5liK
ofdR7ZW7VXEwIv1kM1tihTHSgk9fm2pSSqHM3m6E7MmoNygGWhkdMirO03gCf8cRehZPH31cM3eq
3DcaPK/v/Yfm3X0XAmoRiP4+FeHWLDNPArx0EhWj3bu/sDPVaJZYyHkfQQBnixwgE32rvqxL7zHY
6YSnx5u1D8+qI0JbVBQwCdwS27S/Xe1M/94lnRebER+bzw109G2fg2h9mQkcSvpv6i4cj0WNtQdY
nz6BGU3WYgPJiXlVxkXJNwTCKdA57X908LNO/DDfEtGgwOmRXdViv2UJx/Hpsq1UkcDt4gJGO9Y9
cLsI0RWsNTHHEjgG8NsN3kSLkVr1EE4zkbXx0wPodVXrTYdMnz3ZYa1+tn3FV4PdiHx03e5Fnp+O
8+o7Q/oiLow0HxMLl3OJZpbEZ8zd1n0xGwQPICxhN2qDXxWgVKEy99yROifxtFosE2CZbJTIg+q8
huufu5qAW3ZeIT5xPvTzo+ksafWmC99DZ5Xw2b0vnpXDLWVgWiMNezwiIXAOQqCIU0hKYSDrONl+
+0dFnLTnrgCpv3AOUgQU5CvN59LCEta3gooMc6fgRl/oOiV3a4SAwQ4yZiNgC/a9DAu2hn5lMjEW
/Ioo09SRcVnUf+F9MFdKR8PpYYZElWnK8vg53GeqX40V96aXQN7CLMmcc1iIal58GBZ5xtR6YamU
ISzHwzAKWF/y5CbQlcTTKgrtGrk1dkBzKjJVR3iIO/PBycjRuYPy+CVF1kgwBOyXKvALbM8HzFxJ
ediGzMqSUCTCbiDnXjVna66Zwq+AozZBWZkIitoLVwimaOUnmhFieb+UxLdhF7sJwMkKy0Ni+iOl
8xhKTu563+swm5DApf+RyYcWXKA9F2gy9Lah7uiQEHYoVsyCD2nU2331ObwSsaAvZy934Xc/BX+G
x9Z1WyPAQSsvKzNr2Z4uoJrpANIMwlcuhCHghHHTELAGDI9hW7K7YwOiqfOHxXekSOI0lXM69pHq
9S71nORgf8+sJnxHmoXo9kIUoE4zaWCoVqWzxOUymy9igFy+z24SPdhPU7XukT7qI+u27ShOSLQm
mp66sH1K/BnokLouFjU0g9D9S9xgDYt/8BIb0W6OxN/xyugeMiqGioeGG2znGg7CXnJrSf3eYq7Y
1lImhH/vfbzx7kAZtS2XfGIyFCjrBjrbWuR3WkGsBpn4gtMQBaZVFol2VFLlJP882rSp1CT/F/k/
tm2F5zkOukvRTNboqSo6WlzaiSp4gpWu30aymFvfq9r/d2BTXww0obGs8H0aDN/xQ9xMmCcmPPNk
YrnpsmoIBuR6mJq476lVi3o0MfW1EdPydh5Z3X2z418yG6x+UtuqJgAmNGErvmDbkXbCTtYQ6M6K
B7Kl2DlogElorz8M1HGIxCr39dbJ1705p9DHS6UN9vq4bJ1A94iCsXOBV1csEscKOy9y2HF9AILT
w6+hmp7YnZEOKHr2cnMmk7dtqA1J1mAXI/h7RhLOF38Lap5gBP3EP1lPjtum64C9V6KRpWv6u6vf
cSq590NXLiY/ESsYq2VdvHiY7mVFeKA9NBPa9OxBKp+pc+r5XF0ToAWfwy8TsE1yeTKzz00zPqx/
DAbMLFQPJnWAMEnFn7tC95/xKQ8/cGDMGFewa1CD2xiBs7putVjRIv61mJUDjfS0RIREsMC1RCXX
wPx9L/1bWvDwdg+R/0Et6of6X1VGGB8iwzYdRhk2kXYsglbEGVc5MMgehNwPnVeNu/J/C94+XjjF
/tvHyY0OpFDYSkTlhCvvovUd5kQA3QbgzFpl38YIZ0ZK3xim+r415Gb374fsMv2GfcULnsNUAKyX
1kNuMZPj1InF1PjkzmMRXODIP6ff1gBwefjsCHp63amnqibuk1UcuZth7uq2i9jdk2BjgG+trsfp
CdJ+6sMx7f+e+AeLKffhiZC1YmLcF/gU8ivQQiYd7KrXOoaxO22LqL6Un76c9fYt2r7NKNyJbyo/
V8a8FTndhcKOZL8bDywGWEvE6mzYPXX8fy11v5ak4a1TF6B2TlGqOlVvJrVpOKsMwgYplVJJv+Ck
wyYpm6AnqwBKbNLUeFtReGtKSXtZ5N1QJvBhWJpdSgTDC/kMeYtgh5Jtl3NmAAaynoCE8EFb969z
OmqcQ3qqB6uf1eFvrjjGYIGSH922D68ayGD5oSoFkn4Kl0Qp/sZY9upGMeBtsC4Gh/LjhH2VZexe
gJmXc7W5EHGHdP8A/QqwPrYmM89zdDZ971NHiNEVpR6/ZYAlh1N6stmi780DdP2j89Dhr5ySgUMZ
SXFE4auPEagnnJ0DAh+DjCXNC2MyAkXi0f0pQ+4DSnlZm407xNAoEuJWSnRYs5qIRPvEKCxKEspX
RC/gUevpnsT/FN3s/EdkgTKdDzXJvih8uV8GM9xBKqWFAPmPQGjyl3lYM3xG+L7hoPjy1EuqDs4J
RENVhBuQBQmWfTfj0iPXIWUMuHtla2KfmRzHK3f9IuijE82qTDxxZWk+QIPPYE1dIj/LOUUSb6ye
Krdm7TfBclGLbcH6m+vEqdcX3rokKouA0vnzOmMeiGl/b2HvN3i6lNQXuLcBklZSmXcCaB3uErY6
iM9WxOySp5U0RJ/9XR2VQ97v5JWAeY2K37qKKvrfXYaxJzrhuFUUKJMhwiYmZwd3LxQo/CrM+JeH
OFULZ2Y7bzfqBXX8L+UD0FFA06WfHBMTDDdXVKmWyd1VnVotJDAfHYOvlnEv5Oqwv5DgII+0GgMV
rRtTnsor3y45XkvsXxUVm3YiRNhv85ZDx87UgHWs6mNicUhb25oA6rbA31v4mA8DypHCBiRw/sVM
K5t/JJIYAdF6iK7OIWQ1FpxpKGs//8JuzvYBiXHTJr63YoPU8IWcCa7nEqfxbaMckhR8UUj7CTDt
yr+ialH3okjFvyRJRFETTf584DSpb2V95xQGToTJDr2BmuSChHzPXVAF6dPuDQKwZSKNa7jOfrK6
X7fl6WfoKBdDLFmBAcOdvLlqvMcu6W4I6pLCCO6yB60tyPjJcJBm5aFNbiHGzsNgIe7I+mOZ1Khj
ttzKHmJfsqC6RbHQyoXeG15ervc/AlQatjfId7PaFUMyLjXPWtlIZqxhLKdb/UvFZ0kkho0V1WEQ
KarQcSso3QpiLHy2S610+XBTJr7aOvLuI/EwpiFvBGUYuXTxf8y2S7OgmJVzHlNthyEztdMbMBAj
CBMPqY4vtG3vFSqq0MVViSePVk5NML+GGf3Z+s+ddFK1GZ3PmtSPSTgPxz5ADtcipKpKfWeTAUzW
mR6B03vq+kHw0SD2nUGgPwRhzrxZQIOgyJ4SXU23KBnDkpXQYMIC49s8n1em1jBPau1LGXw+atLi
yGPhVmu57+8k7YfYQbAKUxGY2l20xSdLRAFawg0j+rwphIGCJlGV0b5lLDMtJBkIHI0LYjZmH1S8
CJC5ttqdw1i27gUVm5AFrOkHvVu4b3O/BmxLRLI/+0F+jTfxFy4GctvxbbWV3AqZxw+U1HASWosE
QAHYWDKEfD8EafU7vzqb4g6d6ZHcZp8cPeY+H/8Q7wR23L01b6cOM4xKUW4at7lxXEk5nZp1103K
LmSKm93KxN3WISCri9sIBLsPm6ScsML/P0ixQ8yCJCDNg7mBxjEODzqRbZmSy5GNnNeGHLYZYUwR
G9QObTYulvJR2MV1wvtGtcb4cJ6Lgm0fAqEHu4f3iOHO/wxvei4/n2LQAIJUOHEwS+JDigIbWuNj
dE6omza9sqIsKjL3hXCMh25icQACcnjQx9JutkXSyQdH/bbHOAAPXuy8srzM0Zvb8CLQzgrKJRwh
XixP9iDD+LzkL+8S3wIlSFizrcW2dX582dm/zRfEBSrojtkHpXcKJdXjgaTc1he1gv+wjNxhxfhc
9dYDxx4qJfAgpX5ygMx48/BdiH3dW20edHb91NoJuVzaTyWOyTSq3Qw9SHNmy4QOP4u6SuPLHCEM
zDOLd6U7FMAJKpT1ZJ2yGuDt+kNENqUxW1G+rzao66q3Cj+yg/gWJJHkKgb4ECc6K5+SZiS4PeN0
shjgbNE5j5ElDmVwMI3Lxgod9Db1vytP8aKEk5/YTcv891lJ9xZh9t+Ryer439yJ/Mv99nth/LVB
y/Y/+fP/2JnBq9JW03Zsys/g99OO1ArP28or3ZVR4OctcG9YgUKf8pFmvVraObDgtnN3oQwNXywq
rAKVNsnv8VhSPf7GYJQo4Bi0v1fhVF5CnnIph5+0y2rdsr7hK07etFKkHiAJeKSXRVU1YzORwK2L
Y86S7tVegpQ5EM7htdJ9Zx1rQpNtYdDu72Ix83GGxqhXtXn24tEQYpN9a9pLTqH+bKpQ34zqvSfy
ee9l/PkgVBdxjHf4VpXytBaWSQBuCAEDO2sanUUAUTA+6pnuXJDn8UHehjP8Se/pdadYaeZP9HMi
cBzlbRTeao++vQGT9IIa010IGgDdJgY9MA5iRPIyuZGB3QtlWo8STGMYhvReJlGxUCpsw8Dn3Nzs
Cv6IzCF3uVf9jHu5lXvX603GUkTMl9ldptYsdxdalt27QhtuZ/KK3SBoKctGq1ynGEzHLDJ+50+h
75ZUACigw8BQ27cElx8QCCDhxgkK3lnAiR/KESnEAVJKf5CE4Ey9zRiUMMOFSbrQb8Rht+PjBKt8
UHINEKZDWwRSb4KRJYilBh2S5jIgSEmOAk0Mggqs+NTCAA0NAQAtiUOSDQSlDN5O5dgxuhVsa2dG
KqxZXEwyHCZj7zcLwC+g7pXbGPafVt7x/hQqUihMXkcZs4nrJHjFGaVQXdPsZ9R5uFEaOtBVPwfq
ziMtoCVstZO/+PmpjKBfAIjMThx353KhEXoGDW8qXTs9Ah8pzLwlaOWv3UE4Hzsmgc4DoonBX8QW
+Wez1Mk07OnN2vQ9zTuPudX1GAd82IoHyevfsG+HnrOXaX6DCyZBZcSL7fhego7i5oop8CR5RXln
PRdCKL9mzZK+WSyRxrBTCThi7yqyFCEziuYW2jSscU0PzuIu8rlr7WR1QeF9LUVg291r7DSrDdmt
b01ZLkJn9bs/ttTgk3sc5NZZdhkQXtfNIM+IcVrMmvi3tRD6qOB6zfbPKvGrljwYz8OPsOmn9gtU
tzxiZrm8YVOkpxxIz4Wt8VPImKuC29EDWFbewYSzcj1RAn4ZnHJ8nVCfxd2kSWZkWtMwvkUuZ2OA
NTSVXEpn03Uv0COo7DzRFPb6lpMdLMLgrEwpzkTMy7+APq70C55rRmuW53NWTWXKuuQUOpncxeKK
ZGrx07jg0VeJJOrXhqekrhFxFKxbd/36L0a0gADDkFCK6X6AvCTLxkG2mzpvG9eSttJJOwctHj+s
i2gFWcSeZWo8DSGC6qwcyu5/OBCfR4NiV0BDDv+SUKUKe3DI3Ooqb02X/t3f8NJeAzUZAoaKTixj
tsZ3jff4bbClspmyttBDATq+01XxUghLj/o15hBVMCKIqrLmaNinqQnW+Ps5WbXIauSuCmyOtXOA
DjhJNIGM7iNLt1oXwS1fRnJiXNOCALwOsl9FUsHJy6ijJzw+uhimBsGgqJBcq/PgpIm2Akwy90kE
yiYyVTbP8LGX6yqQtvXTtnKpCQxLlEGuyin8tyvNmW2/Q7RGGBXfuCAQyxnDrtwEMD6jBgAK4xm6
o/z9rDEqKBygUCMOeQmj6xgD/BlCB62iHQ0yABBzphVKvA4I3TSDSk1DdD005Zh5wOj0+ixERUAJ
TMcliwDOM4DnCr9bDIH8ry4IaJREQB9cfwWskZU28jSyAGy6jdU+DlvUI8ft5oDO0PrbElsZ88hS
cZs7N8yUE4FKXSFIqv81OhJwYWy4RjEc1zJj51yzirg6ty7YHThO4/krptJHgZVYSL248Z7o3UEb
J8UHKEluot2GE/KQjkXYdz3wmJIKU7+7vJ+fgDRb71ayhSBSIZzJXlWeGs7s8mBf5O/r+J5Dnal9
+ZlOEk95MXHqe0w7ljIAc91NvMCpV1GaQTGAzyXjRrrps2JfHRzHJhIc+GLMFuBBcUr7PC7u5WfV
xnEZ6JdUAAVyctGiH6IlFYqA6j0UsXw+TcEkbqrtw2ypZW7JxQD/c5ZFnzsODhJNDzDy58lj7K2c
RAv7lBJQYRH1dZxwPIeEELfWQK6sPtXtIQax8mh3tgtykYAM/gdlthZa2sBeKEEM6w9bPTdWql//
EIlU1amVPS5rdlTLRAbyGGJyf8cAXJP8reJta3t8sgLtZ4m02AD7SdqAsrbq/YTvajIduj9XPvIS
pPmm1JAtiLyrbU24vWVLyYKSqaQ4ETODHnNPUQqdRV7KHbxYVeyi1nY1GwsN1/OgRqVAXzuO3AXO
AHR8gsGqIQGXS1ptvMjp5+ttDe5K1qqV2YSgziqFJvOKvUi5FCh7foVqhngTe1tfHdkoT5hHPqsM
Y0bWzKDCc4o+VPdO/NPOxRoQjL8zmdq/dUshm1BwY2ORtd45x9RcOOtnBEcipovdpU/+P26K1a7U
ubfHfwpZ6urPHgfg+MMyyOHizE8wbe8i/Dbq1PGsbIR+ddnMBpS0FHKalo9PBLNqTlU9dRRP7EEs
+M7jT/6adTCdD9Z06cEw7Avb5vsZeg8Gv+UTGrDnESL9TI1wnikd5PkY4828GabIrS8bnY2Ax/IZ
wR4J1vWhh8kbhuZh4wuM+NM9LGofXXvzmu8Qqx7LP0YZBimX/rr/dnP+6Kz6XnNQigdZb51sGiyz
VrIyQjHKhLe69cMGulqAO2TgxTa0+eABY/p1pj2BrpJ5iwCjEtxHjyj37wX/f1827ByFB60t9Z9h
6tyAQtUzfpP1f0jJifVbkHdSLzXL+z6pan5t0I9X0APp7Q6ijrTRtXaOU5tJLvfkirK8WsYzds6i
W1eJ6rh5SDegIOS4ra0SUZhxrqn/fF+rKTWgo+Kbs2iKkFQ9X47o7dsSTSNUrhi+P4ldNh4OZ5R9
P7AYsGV4y3JLXo0gD4IjIBYj+Erf6OBSAdANOgfFvb0V3Sjk6e/EmiQi+CxqDB949ZMDHZwGO78L
QCXEKWA+Ya1A8/VTpzdyhi4JKJilvZmIlSe5E2/JPX5PN4W+3BKz0h3XtJozRF49FPw+uPL7xdKk
Az4wdMwHTPAhCXBob6CSajaUSftOMdmMBLDZSp/F7zVfguPWJ1kwkrskKPOlRF7IQBXi69762urc
U6/TiV34aJSq/xPd71jnxyYQYI7N+AeCrx196GMI2Hc6E936t1nXyNSkxHTJ5NaasKTSgdQLxOuC
LP53MPwnFB34Uihj26G3J5alG8++CNVT7gNFPW+DruN/Oma+1RO0gCF+ylsq0rFSshvXIu30TgT6
zwbr3iPhPVWbNotwSk8DClxJ80qFEX8seyD/51gHEJXY+PAKXs2MUfdk75z6IJMmK03KlxDZk4Sl
ulHNhdCQH6qHJTwiW35vg5OMnz5EYB8adWHtrikiAZquwufYayMjK2d2Lol/4W6ivhA10bI6kTIw
8ehvffDyLEMljI3vRXWiMQxS3VYE90r0mh+Mx37WZ9kHTgl2ZBq7V25xnW4NZ8ponpPFAjZKOSiw
ZSGJR+v9LUqAjcLC2ksJXYo5Zsil7E6pMhpZh8jHQcljremEUZLEsb4vCLMy7wjGp07g3JjnfiRk
f7+dzcYvDMtWM0B864Z7wzMfp9+eq1/vC3rgW8QCUPrLAm0NPFUYkcXCYn+MPZ0JwpCaAC2lSrAa
BYFiaDop1OwmYWLSUp4iYfIbH44l/QSDSY7edUIQOThUlEAcO0+ZJQw3CmobUwQZW5R/y1+qH3dJ
F5BQsKYslSIxYRRofQX/K+0beepR9sdaNg07ilM4hFPtzaHpXLoJjjh8aMfpALiJTCfUPqXm5N+N
vS5M8SFSVoQ4Oiyt6LZkawTKz0BvSgNkyp7Fts/aoXLScbzolTf7Xba9VcKOCNJI98BFvQA04Wz8
7JvgBDTkbflzugNsZOeNnnExOTwQxvtwedl+jQ3HvJcZUtNw3mtg8P9ibslq+o7GTKj0OGtSMQFd
NWSz/tlYZqLozCA5s/gHmU6JaB9rzSQKVola2MU9Xjp8vIDz9CAPLqMfvZQwdR+siKZ/vv0rETLd
vRwMzAbSghEu4wQmqMMEfMABBomFxKd0bviuEvPe9Kg0k4PwP+Ik9hWrUqOJPYV9GZgIuxF1wxgX
UWpuvq0FZFB8iMiP0kU9UWxA5N+ZvHraSDGSO9stqh45lH8Y4dZmTGZtxVGeqkgUmURUki2JlxNQ
P7EMKr1F7xaEejdTvQAXeDzEL00eTQ4whRiP9e2DfKpJmDkORDZALIu58DXKsYUgoGZbWVAq9bjY
ki9mtqJ3st8+AJKDKQItrYRyLKKuYC4D1H+K1mPu2eBM2wXxOfVW110oXG+R+kepeC1jGBXYrovG
OoJvLo2na1qmxu/9rxYYt4hbV8aozVhdeL6E0TAuml0qDTPA3I3UkCubT7t+2ZyfcuSRxl+01F2s
Cq0aoBoHCy8ARbqmMmsuQaOhrolW9Y/D6SedjNORqdwZkcSaStxOPa8ooLBMJY36ToGjwzcPt9/I
D/ZGUIofEx0cu7xklT7FqEyiP33M9Yb86Sf7tlh22aCvwV4zrxsYsQu/He+kWzfEpW0KRh/0o/zy
s3sIfP9Jf/3Z+MUi6Lo8Ggm6vqUXHULCLmvtVODYfsrpuULKUF9A7G2Rj/Y623xGnfZcaQOsKI+T
1/0ydxlFPRZzf5oBpBfEiFqM5iG+MumvRjcT8WSwogexSM1uCQ0fHAPomy9ScLy0gpREn7Sv1SP+
9ZRpRjElWBJk/5tGHfgCF2WQOzfXOHdK9phXR9kb3OeJlPJFb+r6+UXO+hVnbQfxpKMl7qfQMKGD
6jGWPptVVJDo9QnpIg+06XvTNP1q+WARHyVuoUHfqE49Rlu1RuL1qOUqra+0nRJKe3ue7IWV/xSW
6hqjREXwA4z3n+J0+gSDH9qRPbNIQ0B95xj+dVbso1zURDo6oQUEGKprDuOEQwVNX2xB7qovisVy
WtUoJs7H4sZ3DU/IHXGYv0KcM2TAbmLYciuOzBUgMXu9CZSrn775AXyTcZoQ3FiGRvJ0kZ7NSJG9
a6CKv9z4IsmIr2cTx9ZljeBj3hePnMJI7645GvgWg9yJOmGPAyeWsdir9naDcnF9u+VEJuFGkxee
EXnBkpGgQXS1nW8INfZGX7MP0JrQSxXxvpEY7Ap02kFPmgEIm58zZoj6ffY6N19T9PgOmB+/Clt6
k8ZF+SmKFrou6cr+ql7I1V/Qzaw53ZhdznE6HVpF6RiLoOBqgV9hY4ad8NNdE+LU7x05+Q20z9la
Nv9Txav3VVFSYaVQCO661RWlI0MVWGmt7eWFZ/OviqFF70FNfdoQ4jhIrPselcdpWWjH54dVWSGR
1YbPyTkni5XkiOD28LmEv4c24RQzh1KfZqRG556p795PK5bKb0uNL6KeX/Id8SntI5dpK990A4+Q
XudlK4heXeJiDbSZ1Lhg9boRh/SesMWMG2x0F3SMhloqUVMKkMdD1+o6aErxX7gvUajp3QkxrsX3
Z2JLJg50N/AbmEGt9XipRmSbfrVIDAcDxSEpVeznqI7wolTBPqGj4uPEAAyp83wPjh8RJOQ1yonS
bxUYZcki2eFLvVl1X60sDBmwnyrfl1B3S/sr43aEUJ3reiPfrLX1SZGOkaB+BwD0i+TeUQXYGsSB
lLE+QRUb6TIuOm9TvwLRpcYTBdNTqbLGeGtkBnREkgckVGwS8HLNWuuzCdoGZ1YjftpHbbhOIOmH
/fxfzugXOXXq6hQo07ksk/llcemaA44KGZqWSN1sO5hb5VaOEpHCz8K1kKbLrS2dnd/nHYSSLNy+
V6PFNArmSdkwi2vtc9aWCSO66YCDD17BTF6Ma0PRnh14aDPA2v7Ac75E/wGa0Qq4bcZ9GcZ4gJu4
cdaI4eugho1nKSXJf4P1dU+0TtJH5SMYTNPXnwUwKrR4GCQ+pVqDLMMJXkOfa+kdTNoEU26jt9jv
YtRxTvLlJSCNto4vIwrvbutTSRggruLP/2oVz4d77JaIdkKsz23V/tGjgsb4f067P3CWrEXzP69x
87y4lX6UbyoxRC32siJnKJpBfGLx4yKiFFScQsrkHHNEn19oN4hAGO05kfbiwnzg2hqHrl0Fbgs5
ZQq2i1D/jNvBgIYbLIsnIgK2bsYDTpHYUGYZyDDtlix6QI9Jexjtt3Km0AFC4+ko2wCe11eIdybk
e3RUKFjNUsWUDF2hg6hf5bcst3qp2EXQYmaIMhDpDYYdDfCRdqM4qAJx/j2yUwG65XtKu8PbKLqg
oTQs51XLhojiTqCciq3snNc8Oelj5S5/feRP2+2y6hFSZs6h+7To0CzfowwiLP5FwJdsmQD2hlaM
8inEfGpIfP39h/M78CBjfGUN8TR8J6P0XZgoiZtM3K2GAFWAdEs5s8ep/hxDrRPe5UdPmrCOWLuu
UdwH6XuCI7Xy1r3fwiM1f8KH+m2waaXSnfFRTPWn2EhCVzhlV2/yVMwKHHvzOYyAQ2jIeB0+2h0X
m782SnFA3KBkIaxlecxcbBZzzMc2dW0RSMhSYL/7XQ2TirT1SinIKVmNpsMlYQloYT+cANJC51Y4
LbEpRFPLxJFq9Yl/1ZZBvN2rEcKsOZKjTb57D7mQZ1dSGCAHNqbaXUURylwxYjG8bGmK4DcDWAH7
7vZTPGVOocKQTDbk+lwK1E3GOePLHnK68pLM7TgYYiWqnDZ9sWbO5XCH/HzKrBgMkz4+vPi6IUdA
xVZcWAmF7LIxiedaOdx23+JWbyvJE1OnFNf0HQX4lZLzfne94TFoUlPrJ1EwgGsYF0h+3NFWeOwP
fO5knrpZBU+RLPp7xsdgXjSxXbYT4hqHbtg+q2Vy4F6/Rc3q8iqDIIZAQNrxSvEpuKdYXdlaZP8z
EuWwp/Lux8O8VwejWN+lJSj3nSwgt8OP+6X+WD+slItM0OELfrutN+7VAC8t5QbayXNj0+nS/sh8
paGIBrd6rDBP+JRr4EozgYRc/xL5RwSceghOoJmHnno+13C2EM/m8z96xnlfHlSZ/cE+ZpfSs7R0
Q+UvAdA3UiGC+XiBt/hogpzpIwGMuADOjn9YhmWmXBGuPtAljZVHEM0+3CtTVxp9xvop3FD5YicM
ilapaq492CO7TieG52vJ7/HBWI1SgmHoQUqXdMSTBwwNQbuwQjkXDwhs0BuHRTQd9t+PvNUrHWxp
q/UBNBrmeOZ5i6D8CbL/rrslAiIboZWbkPicxNn5iTpzRso8RH1WEG/Ew9r3wvKZpAwOaz+pn5iN
JWwyH4BNk6S+EYYuaZplr7O/dWGFsg3UjPRpwVifp0hBz0XRL0llXxzm5oM556t8+gtnLGiUYcS9
C4jk3paPJL7c0a4IuyhiGG2HgVWA0kV7qkUiWREoo2Mpfo7+dC4P+LspbuufJcN6qOeGfFMKr9P3
vJnwO4P+taFjhAsGP1RlDz+g+TWesMbmrHCFtr1s8eadcfg+FM20K7mks8k43P/fIyrxrou+V8IW
Z7qe1Q6PsT/YpA9s1jzrctDN1nCOxxX395Is9RTPXKgh+AnjLEjW0N2urJ/bbnK2G27ru9qTankE
NraFrVWQvA8Ev6iz8OI1oSHOj0glYpv1zdMP/dgzIvhMRv9T8r9iz+y5nJghby3d96r+gQUGc/vK
34vTBVLcfjWlmaBAg/hgoDh/H+9WIbYCkG8fjL/2CtdYprYjG3o//a3vTRyVXdQJelvyIru1S9M+
gADdm5v4DLy38TycHkkAb767MgcMm6W58HT6vRqB/4RMn42XGw9EYAVxCkGeTT8cHbch8FODTICj
X5MzCJWZ0Ur2JgoSFNlYDKr+hHMt7kx2EySIyZ2VzZpWNMDcb3xHu4y0wuJYfA0Hj1w+UwHHbRSD
o/KQXzmW0ySHWEaBsxEgKCNvjDJB7EJ0mVnmVc9l7BFtSkXPd66xsqu3h195QA8wqOX1WV7noTMT
dW5KAhdQ27p9E/hkDOpOiUmCy6qglXztp4mukIh8diVLGYaT8fbeDNgPBzw8+VQqY9LcT1uEzSrD
C6PXVQi5ZxxIkXqR6v61kGC/GY9Y5PDDw2Pygs6V2XdVcAx9RDUE3r+mXaY8OVlntMulXn8WSHrp
ixVwPJhUIJV+RPf9J0LqmndKSxHfzhu9hJUALMNuvmd6+xlSF3jF6CNae/eGGTmuMKXhPypDC2kb
GsBpirhJgbPoZyyY9uUqTmRuC7YGRokbLk083MuFiQ9LjQjbRogHDCHvze0hO2yBAO5oDAzlEwz+
Sv/sTv2DfgeohbU8o7UwNoPNXlpL/Zo1JUTytQbaWDh9Cse8JMHxY+DWxyBIFSg9BCpTEhuh4/AA
OTZvMYik5rIUulo05F6v0YYtEFpOOCBjEh6VPdUn6xebx5Sj6X2C/ez7H0+P4orwcIuS7nz9qseX
F5kMYyhawMYX87IARfnamnwK94TUhSqJHG55nCeVYLbFjcf3LVaUUpicmJg/eSY507loEWkaOP5F
KEPN6B+zuQrGIwej9PA8x8GVZ+nqKL/9Ir17lQ9XXQuotfjwGcY8Bb9qTusAJ/UJvLPp68pUAKQa
kQV6QZaizxS1RXYTXYEWqeYXDGxPIikDcUifLedJXS4OrO3QHS3WkHmYu1DmUXJja5vucSWpqiae
yXdvgaX1uu2gznS22Ctl8OeAS3SyaUnuhcIt1Aoje1pDpcvh+L4ZCkpjEjRKNTxZaju0HnQbaAvw
G0R8gRk4bXieF8yi0VY68F9ufJcE2zTfYXxNqTj+ZMgN2m/FjykRF2uH6AgbQOf3+OY3Wnd5Hmzs
FxSECyepitILo9o/uA9kOjXLIOxo9fh9aNjr0ORwoiBXu6/nSQbCTbr74Gl33dXCj/XJ+PxRYas7
CtWpEF0MwcnHRqdjcO+gzNyEenL0cRFcpYYKhG7l8jAWvOOIBRUEuwTj7FOJvZ8e1LQjglYQUpmA
2ctIOPmzOFJMefoaoj9BCElCPrqVrMu3aS/fT9jj9HNN5lXaHQtBePhrwz++lsGS1K+VZ1jB7aK1
Ia2/Qs4pSoUQBkw6t8dThkG0KPrdOewt+65ua7iHXVdoeB1yImfRvBb/BfqURf+1+fc7Kmmv1zJi
lvYjWp9M0ucAAQGrswQfn/hLUCK4KRzPBfOOJnDWj+xaNi1RcnhoAw14ijtLLZvXdel8uOYLTRA9
yaGcnE8n0rc7vxMbwycIBkM8d2LzqfMpwNn5ohvS7f7r8RG2I2h/nYCZNFS0lczhdaJNKXB7f9un
qL/Ek53j0jNQw+ir5bYcPHyw3Vv8oiJg2aOeyE7STUwfUW4TqJlls1Z98no3HuorIegYeI1q9Jl4
GEe9tiirYRen67Fnx8zq5vX8PUigm3/awS94afWRBPgkYiR5IMWkT7Kd5ff4WvMdExhp42GyI1dy
84n2sgO/qzLW24uQ2Rz7Wp4shzLEoyA5y7vx0hraRc8mH0FAxN7LyjpSnxdPEXiNZlOcwprvAnqg
R+MMhZ8Bwu4998T5K/hNsBUK6LsA8dtVyqSy0yub+E7OsD7Yz6IgqqigFSJAbJ6N81tzJTlFVSeX
Ive/31O2EhRg13OHfTfMsrDEgxv0CtlSNpRGUJT8YwsFFPqWzC2vpawMnA80cM0/2SBs24B+6N9t
Jr9mV4U3AJ/512P1uxTPF3th7aQMuhTqgWmkt2vcCkPdCjc6wg7Kb0tsAu4bSG8ZZQ11YfSUzAth
iJ/94SVMUsPgtc6NlJLmqkRXuCdNPYT8yhfdsK0xrPVHV6D/oXFwI0ueEmKwRLkj3TwVCvVmC0Mk
KDryygn95axDdGlI2jZbl3x7g1NUNOJZBxOHKjjEsH4a8LGj2Lu8iq/0dQC285fXl2rNQnkAl4ED
qlEyIa144rqBpF64+wVUtMzmtoz/8cPX728OWm02dhVlV8kni89XcraAmPqZ9vGPVaslym1U70Wd
CxKq53lWwawj93ambEUp7zmJEXD9ysynlajw9wflxUcdHwwc/tbnLyX8sz4abXuI5AFSO0Gzsi0e
cWk3E8zYWVo2CuQ3OFZLstl1PeE3InBj+rRLB8x0AWnTFssLLW9rJs3mFMZp7W3n45bSBj7b6sUo
AKYg7400rNJlgznQpzbwV7KWvEsu7OcnMohu/Aws6xAFXcaVEh3pOx0EbpS752eq9Pr8xZwbkzNv
pEqG4Ym2wb0N88un6OjFSaRMrDddtPyN1TjJWJjHV/CyN93nSbjHbyY4zm/fUjgSSuNfP79dzKEw
n/M5mI3vmqGRGdr0VtdEYTDOJxO4zDqxeg9YOt6Z8MO3qmYVvTVpXaPmFED/OTU/pWzqoAQTG2UH
cnz8qTKL3YO0jxCUvawTj6cD4bdbJHlZ8ok4xb+IzI36fz299ZSwEVQSH/1su6f2RUnmzlLXKLwH
5zN+opHXElyZ6ifaTyA8BOSdH1bUMOqmzw0em2qjrgfLIVWxj5GKWDAnO8gaG2M/3CCMsnmqbiwR
u5/gPHAuWBHqXH0BZ/XkIXhx20mtqNcSfV3drr8aBXPeQBUgEeJZ+7TIvLKZiXkLGOe3SH+JgtTt
RqUDb/YJwnFKqiOu3BghQ0Z9U3iICcEog6UZlw+G6TqUB+biAVVYBvMDC0u4iqAUtBZl4QioVF1F
v7s8As6tVjN2Ec4fWia51Cinsfjerozt3ImbZTE4l+rx7ZEOYhbtYfRmBGTk+5UnR44N6/HouSU+
TbesHH7KET3J69zSPXX3OTtqj6C8bn6NchAsKr6MKw2pZ+BtZCuUKhpGl7883KBNn45aUZo9f/WT
acumNkj5HvpJ/+GIXEYBZ68+HkyPC7GDVPsYWal2ZCfV/sxfU48vk5uoPKeOvX9dFLV5DKD6Vf4M
umHjIglNYwj6+F3qOe8pxDEU+6TXf3g1NJT7HGRWHtH2PBGA0SfZxTG9h/NQpxFCv7dp9Zu6RG3U
8yOZi7S/ZkZzZv5bKWhvm3JXMmzVpVNUxMpFQEgXRx0aEo951RS7RjeOa3dS5zetR/c03IoTQRT3
dcigasZd6cYQf82ISwN/cITc+ieQtQPiyGmV5AGPD87FTwKaGlEUd1aucA6bQEdq+mJMGQMIIOVb
jD/PzvIBAeSK6gnYF+PoDaYwfBvx7n4EqFu8dascmle0YTsxE2dyp8dcOpesl3DikKgmOBewIuFq
IlQjYKAOCHPy29/BHUvXyCRsgf0mxGkyawl25Lf5GnPdgFoOj7Y0ywhvZjHKDFNd/1ggrRL7Kd5d
8Y18le9gqRBP0svNUn+9lF/YdGK73PalCjQMzPNA0MErdEX/IO0Pcn2mt0OrbvGSpkQU6PR+WSX2
feNyD3TXHr8QdFkAUauOL7MpdZBfoStT9NuHSO45aNTXUjCxr3giooWBqUaNMZGIwVPyE5oRfedN
0aR3qEWHBEEnZ9Ft6wpOIMfq1t00fkN+ICsukqeUBqk5A7ljFvAv0S/+yXHzsJrLKjWhO4PTAW5A
nF/xuEeADqrjZCQPeWvUBbSDd4t4URXmG2L/JqB56Kq2i6RuXJ9d2UqiG1TdVq7mX1Jw+mfrwYDz
jzS0+Jpsb4LQPdt4uiuPzZNhdENxXzP2pOgZ7xXE3NM5NQ5BnM/enjwkaIwZNh7r8NLWtDCMSby3
HxhnkLKhjnNN08Vv9dMBCTOfFkJcrBeyDQ6+ZUf+tcwDJ6xz9B+gQKsmK4Hzqh1jb0Gg4rKqD/ni
PMh9pNr6aH/w0tUHLF6/9UyEglNGu9R4FZMpSDJGXZ2Sn4xDY4VIYr/BAFpoqjKWjcQkTftUS0od
UmU3o7f3HQ+XylYTR/UFI7gFDym9rF23yg5eFCYQW8qrsywgM+U2QxJlPk52L0r+2+MLI4Z7Rn6Y
mIo4DRQWJA/xb5wOconBheALUxovW5nY6JkE3/LK6+ury9a1Qi8NaPjZtVpkmmg/Wnl1gtWlP7xa
apHELtvKFx4gVUgDsfDofOo4pkFZws/umtyiiPCFzBnnUlt8jXxALjr808G7kR5Cd5j8261eKFiV
94Cd75tHEN0PtgI/qOx4LsEL1CWOJUoTfrzOmE6qsDp3xFHMNapfWsn+L/cRd5IpCiA8ckqvGibG
HxSwvFWB9YkV4Ic2UD2Hh71fN+9w7PjGZybJlWHpKmo63H9rLaoMyxgRcAbLXwfSSh3yeu4I7Rqm
DisRGviSJ6d+cwLKt2HJ4yVIAtKKnHsTH0thy53b7o9pRnRDFgTxJ4nQUuu6cibe1OEJ3yEg4O24
Inx4ItIUINvizXthDUft8AFlX5YALhBGqPQIP9YYe8565p6DLvDgVAshOYyfT85aAV99CmMnQxDe
LJpE6Yd0RjNvnofQnWTLobDGH3TOnumA7aQt4KVz3rvQcyGluHWNQlY1f+Mzbp8SgB+99eh47ViU
sFml2cog3o/8fetRV88qqxre5yS2LZTPlgVFY8JRbr0QFqFqkpdenBadI3bzmlmFy4nNpXNlNglp
tYCRaI13KhpoKZkC57zUW9hKxgjnljtidIL8Qv7VXcUZyk6oF6tK3nic9dRtD9h/Q08fwloARW1a
YvXcSbRK9ovdTI47W4Gin4crnGh0MaGCXF6sTJt1wUFjven07LQFsrWdrw9t4Rb6UztXp5oOvc+N
dIrhDjdFkmtL7c4D63DPWXK5pzLBjqHpnUyaTtW28GOJkpJOIPexi3Bq9p/KNNxv7hmNg3CAuJmD
Ay+lzpG+3ZQmyxDBWFC2cP+dVAFP6ZFkRN6l52rvqenBpowOwCcEz4Yo8a3hNzmMR0u4cDctc2jo
NZBCDjcDipLZZXwirC+lJPSy6LlAlovguUmFf0hX2jYUTJSp6anKYA8HsBahyofM+XO+dS4yhFL0
NILOKmm+oDOoTGU93zXh0i8wUDHhjhTkXkMSEVZqNBNyQk/BpCAGreDyUTrq8oLFabGIUqs1JA5t
KyelFHr4/8E37cdyB3kfP3kF0x1cdt1Nt+dcQOsSkohfEIS2YNANj0jeX2wBlwA2kbxKVWunHsWT
hi7jUP53xBielzd8dJcK1tL9+FaxEOwxnPCMnaqeVccMh1nQohhqMLbco07C9mPsD629v/dJam+n
nRGiFbAD67iMw3/hGdE1u1lzTf9/DNX/W/tj3Vjtg4szKzB71Gq8F56jf4A0lcoQuRtUZQNyy1Fz
QaoVxGyJhsH6j6nt8qMrfkNntd9cdyaz9ay8vDYf+nJSMgUjX8CSDxlNUbXFQ9fjEKp3DLG+Y6GA
DaNQBI7rs6aFl0wU9hCeCxcIayhbwXX4Egv1zxGdwkCsnehe4jwewNeD4pwnqY2URNo4nUMGFfdH
qDcsquiqeEfCNh0T4mDjmwAHH0N0A04wnlBUjjU/68GVSkCyCazIKF/TvKQGVWFqtgKXGMuXQnEF
4rqYti8yeQXI1gvtKPDA+w56gdMYq8XR21PcfRBaKw+IBY111Y3g8Rh52UV4mG9E4vUyRW3tWMJb
WKSNodxtvHfXIbthgil5RVDplhKZmMFreG+y9h/LnR4QYN3FbfQLDM2WXJPiqLqlOICxnHzFRzZx
pCzQD7id/uZVh3RAX1UjckSCdc6qITZ/jQdomb6tRNvUJdAr6sgIyBpvQo8Rr64Qkj6b9LGrGI+O
v9Y9EJb7XLoSF5Hwvw4NNCrWU6GjXFmxX5syvvYuazz3VAEmsJJlnSIr4QEyfGAPlD06/gqwqJlb
14vzHrXsDseEutVkwdatB/4zY/T4Ga2Ar6ZGKM2J83WPC7NW8nJm26CK5zNma33Pini1DhnX9d3m
/Io2EpgnyjY7TjXKfc54vMmnYEFVw4fnz8jOk3xQxF03sLb7EA2c2GSuaFziV8weqlZ56K9Z103n
JpMM/9pqfBRZSGfTmcKGWUiwlYW8qeqSdlvJGWd+ixtTtDQA09+a7i50sinS26S5k+1ymX6KOhwa
cjjmvKPNI2DfeLhMklBIC13bIcujz6WHz8icDDB65Fp4iGaXm57OjzP4JDYDHx1u7rFsD6iknIrK
xHnyQcH5MQAMbON+cY2FlObla9urIH1KvohnE0SYJwaakQTPTUk8U88jhZlqkDD7OEQ7c31oqOiE
oQ3F6FdLKBN3Rl5YHKUNxBGmBQe+623auHvTsC6gy0FKNA0T1R1HSf9zlOZmfiYyvVVaoiFz+hmL
M8N/+pw/VX/Zf8S2zRJWlh4g5dBMI2KGIc40pjC4GK/IGwyyULljlvROzhh6/PLOZuZEJp5v/qaw
ToG6bDQFaxdOyUMR1+6uW7UUJuVei61rMujWr46zuSXGM1ivzk5FgrpM/b6YahnTQYnwW4CstRyK
F5LJXIJDHKa9EGX6gOvLMQKy4ICcYABdjXtYleVJdU63gN/1YziyBzBzOs22susDE1yv5jAKFPuS
nuYtjP2kf0sREbTwysRcH5RM8mGEcho8tAwlXN2a6hpelaQtZiSz5IIOb9rYHjpLihKXuKW69VPK
v6uYtnPaXUMwgc93F8j03xU8hnvnyYI+gHzRFsC9dd353WO20twusS2VuRDB9muXHdgVbTlNt+Jd
XfJkYZdx6iwOYuqoHcybcu18x46u8wJo3n+QjxfSDvvwHdXQ1UitiniFFdMTOqccnXf77uiSFUhJ
bWoUleskC35X3lNG6AcyOKzmE3E6hf+oUXJxYiKQ0HOabekmdm3dFM2eDs7FSOkQl+Cq5gv0lDyN
8LtmYW6ejCR9Hm3MCrksJN/QwiMuA2A+/UwK/mgohC1VWUndqf7bX0VddOu7RHScJiGIgNI6BjXA
rgJrNoVqcXpx4CNJf44DpsF2u19V8Ccv5ozy1z/+oeGOhlNWEepr5b4UFz3/T+bXe5uqegzNF7PQ
qqU6tl/KK5npi9PacwGpf81Zf73zGXU6xQ0dJP17ytwMAbKzAVecDatLSJ7GF/XjrXCUb0QpzM8T
KDOSkospHSFxjX8AVab0nt5AMxGJI7JChtRuQBA6gTj863ItrCaGux/q3bEuaB1n4ahpwAnaQImN
p+2mYelKx8jXNwnTB6eM4z0m4a9ow6GoaFP3dcB0jL1oeVt6bqMbwrQmFWUenSZVun+q6S2tZd6t
ZLhF0rfTj/SJDPUdKXBvDvnqGhdRv1DS+HOCiSAqRMraxJmkX2C2FCV8cUIQRPjwT9r1bfB8Wv2m
EsNu35SbYj3kmjm843/SAAxXNXY5ydA4rEnEIzfpUx0LN+5DNSpv5dO5pqeAqbNAtfkl6jp8lVzm
CctFhi/8kcX+P4tZWszUwHs3BvDp1/ih2V/doZ26FOSE+kxVYqP5dciceLuxZh1uukdarH+JLnp0
LWTX5W5iWLBsesMiP+f9mdCns6rovy/PHlbu02OYSEClGTf+8bZD4UJQu6tL9QqXGoQBNOQnNaX0
MQy/GOcn4vqqfwyD8oVrijW8cNrL38VNMvdwmuAuy72qJWeBrFeVZf1uytr5BrVMVHqE5IR3qdI+
I1q3s5qG/NQf6x7kxv/rdb4I9wXVsukFLkPx/fQC17kpDqRZmuMVrTuuof1akXSy4X9dl+Zg6mqG
7LjaQ2wEkJIPEFUGgSnQy2PRWy6hzyN1y7xJQs6TOGGsAEQO3kAHp8lFAfRuTATC6LVODptNQo0Y
L5voQcZ1UTAX1Yxs9oh/yFrvCD3UiPlZHArnvbGNuJyyplVUvt/qrqBe5qgnWi53SfjygUdFbxb3
KxOyuo7FJHHnaRG4c94fASavlrt0HtpRPBPdpmlEbpTwpwR/f3T3mybwXru/vosS8jeyuMu7ELas
rTKC50wKlo4scEi5F0ZSMxhtv3C/14kdo0BPSbOM3HQ0XUK2jFsNoT4qWfxF76codvZgx/8ehNYQ
ESGOjaqUrBBt7AFfVtPl/EmxhbHKdGephZxd4WaDWW4zB1bCTCXP/8OUHrgckcE17Oy4LKIGE/iW
xY0HfpL0JB1UdEai6viPE0TJ1pGtdqCeOdxNF5R9er4YvENldi9Vkh8qflK1Oqs1XKk37Wd3Dgiy
zaimPEgu1w2mYkw9TedsKcSey9fvzvH2pybgMWQa78oiKSVKqiFwa9h7YlNjynABJ0VZm+3rhvLJ
06n3cad/JFWrhcHcnFC+TiE2NLXS6x6X5AMj1EppZH3TUSsEKJwxSCTXua9+Re+o1dmg9asQ791h
zMLcQFzqMPvIcbnhFq8aO7uqLsSpX3X7eFbPWuiHksET20bXAx7csoU7D1wWA96LxRqsuD72O+zW
TUc2neDXD7C6iRRfbTVEMH/2Q8p6K9GYcDE4Fbqkez+K/WoRLSw+5zBr97cRH0/wTzTrJNrHC+lK
a3lAGsmn1G0x8YzesOj+/x+9kmVmZC22QhCh7cTqOP1D4jbMAKx3haw1NEySvdNSK/rtDxwZ7mL5
2oh2RI3n9r1b2kSeiq8IKfZYfBMrUVyz6/TocmlI3tHcXKQqVwk8PmoGY/8BjIf4uG4PQDk2Bio5
D+0bptdd65pkE7AmFMrb11LxHDYGPEF7H3SvUeQD8p3bc6e0ZjveKjNyumkoB+UEPtwHnn6pt8wH
5kxddOeSs8YDVH3JiVnbazOFeoqwHFLjdVRS1wH89Gzxvp8uesATPcXJZDSick6zoMbC+PeXgTwK
jCq9nPqbkpGa4eCTTdwgHCYQpocWoMy8e8jmA1Nl+Xd72WX8Tr4Y0akoE68WYcPlkWqHg9h0aZOW
dvmPlrXZpPoWaCml8a1f2WCsZzEW4ng3joA8oaBuCHGFxIi5TOHQ+RVgEBYbijlqxo/YMoPQALPV
0vFckdhTBKvS8vJaVIboMxbQxUG+9Sv+sIaYG5VGwvQRHAjk5tyn8QqG19t3MzHqvFavZsRf+Xp+
ul9fYG6vFuAq4UQqDjwj7Zn9g59WlRPOIm62sKqsc/akXDqsiutlaCwvmDAVjrohqsCQBfi6KKL3
ayRTt1MNldZQAM3P8xQ2CvefDEjeBE+uIGc1PHc3pGs+BU4MzwufsWc0/DvtdEpcDkcs8nLjGaBu
KNcQP6Lgd04UslOnCQB4phAf9MGaffJJjf/ilVIhHGhutj9PQwo2l7CVj46vFQ4S5QIVqKJy0kFE
CP+UG42NrfEJ2iXXT+xFVOdKEpW2qIcTVdhN7hKtOWXJoHXh9NojN6hueYlaOfnN1YyEU+1IOWN9
gF+gBlb5cYAEAyugSzuRD6N7H3SHpgzpbLrDtLokK0kdPQcWqyYaQ5jxxxZxjrSHsNHXXylkHN7r
9VWBeQyGrGI0448wiQPdlO1RD29PmDHUm90Ar9/UZeu8PznytG5XwmFPfmDqXaXI/Xt7xfb1IOGT
+FmuT1j1MqKuPynNDxfw2jbWfucU2CJ86qOU6ExCXURx/2Wc7JGuTMYOyfNOHlD/mlCo8BG8GKfH
jaNtXtHzcyvOIvQCLOnvAtEYquYLHD2j14NMkcc3EGDO8EZJKn99wOsq/mqRPV+reCt8gssF6Tu7
xKkRSsWSR6oT20Exbe7L+RGXaZ6+M6Jwo03KTrKKk/8X9X2uK2386JMrmwuQP7fuLn+45KVs3v1E
eyuqAOHcOEkzv9lbWnXQlEuLCucDHla641ci6iLxBdyy2kCnUKJ1/TliSf7qR7bQmaXHMQrtKIfd
Uer9TtEqNK3y5TX/GI0ys8nsKQvi9OJFYeUssDm83LGGqabSComd9UKFYXMgj7UAGfc94sskXJ3T
EI9qqssJ3S/5YzuOfjE4V6N1sRuIDeQoj8A+VUPtny1DAWP9eahEvHLivXMPr8hQHuXaI4gFt/Q5
EtAiL0LYvM3el3h27wUezb7e6gRY313vqrEHMnywc+444gjB3ka5QCBpmxASbgcDSlVBkzvi7XJG
z4qd1ZhZl6RQLJji1fLPyg5OmKhhvUbjvoQhii5FedwE9ZRaTquM0HGLt1WK6jzhJFE1I/PEvtSn
n8RwQW8QTskb2/m6tDwS0rl3Uqd+mwgMCOdXUwXhsi53HHcEueH+Rme1BY/l6VuxXUVHHaYSCSRh
7huqLxUrb1rbKmJrm41b4nHxnUAwqSyIQMplNs3Sz5q2Yy0BSNTAWNKHc85kUsZueZ4uKbcijB0z
yN+OxcmvclfTEDaW7a9GNC7gwhXKT/dm1HnSJehuQVJOLQm+lTnzVsrNFW/v/G/GPipQ3DTrKVw4
Q78ERrNEJqaS7MP1R5Q4mHHmSj8wHhQOdVp7CK7JkQ1ToV4Owte+M9GHlhV1icQpL4lQUcxsUq3c
XIUTuepWu6lp7JWEJGt2p53ZT+8NMcSKztAUCAqdC7ZAMhqmgIqbYe/6ZZoitVBothNXG5tM4Ikj
GI+ibxceEr8XoDd5lJPGaWNrKCR99bMaDXvOnSSme9qZ2UejU60lNDHuFSEPR9Wtxgg6x8QrRB1P
crm4mVxfesth62frWA4sFhiyWtA4I1xbvM/FyUWCkKFqvowH7CCu/7CDpqvIyaHnJLdwVAJUKacm
8j3f8JBLwJBnXnody8HwRw7eOqrebcRARV+JW6209Gps0HUM9lkO3ujGc93YrkmBsp+TxMG2iTkN
hmcKZXncMxRJMLbdKwqxTe/vAy2IWL2IgQs8fdT11X2yOtE3RKCQdZmPQcFXGBOoL9AxUhSAppYi
JGqCaFwc8tNN1TdadDQNLwG0AJX//ETbe0XdAqVAByW0MwZpMyqkLZHSygNS9jleqyHZqs5uOeV+
dlVpmOgJOKWW7QfQV7dUZTl4iy7enr59/+VrOkegNu32xRloLUWagbXAbzXByIQoNiprqC7ejz4Q
djGvG70DmatHQGQ0RKxXCPG2nQXpKMdHYDvLqUxwgjPiTQ8wVCIH1nigR4oXTRZssn0RZ5yew4YI
sx5IiLQO8Y+I15QqpfNaPP9gtPkAAOJgQ8zECpWZ6KIDJ6T8TjTy1pgz7OusVHYecYddqbyl8+ZB
mQe5yhjm4e+qHixDpHw9tJck2Vj9PzVQ+UzGO3ly1JCHkbnzoC6ukA6xPrS1R8hc9+D7uYaxEz6D
ydkcxmO42+E2ytiZzMRgaAXIVbKSvV/UWJxBGTAXO0aX8EsRXpcdlJd7W5N/Mb7FUXjrx8fBPttl
SA9rCpmbcqnGmIbmX//kIkX90rUuB+vbyEdQMuXMOdqEbhhDQr8cz/Q45LgfQwVX0BeUvtfmUh4E
o4FtMm2cak7Mbde6GXcB9VJVcFANF0mvJRwoI2QVPtszXt/zeKH+mweWWH+iA6/KcCGj7N+B62+h
gqPutrNLdMNbMqh0YAITU/FYuHxVYl09xUxqxd6Ks8l2ZKetzZuEuMz5sjYeerUm5OPNdIhn/Qap
+8dxnoW0k8iOlmXNLZhYmc6TkHK5xndBADSD7DMJzokyhCa2ZT9Ap695pjWuuy3v8nl/Sg0TC4H/
zgz1eqb/ojiJ86/zL/vj3zpMtkDbwanN4vk66BRQnR9QX/dYp2i0d13Ah2VHsPMyBw3EPBbXXFXS
UlNS3K0X/wMOPPFtvwNxr9XC1SrM01bI36oSrLENocasPCGSDXFUdujTem3aao6RLkpgJoWfoXjm
4u9EjpsPR6lre8Re98fui9+bdqWVuFbiJ0QtlQ5zQB8/y4z9+vHOj4jFX+Sn8yxORoaZK55mnST+
CgrBx1QUTHNvXihlCrWXk4dzGHKYhesggBtSpEc+ztgEpIqJzi+gADPNvEn+t441yBkpmlMdYJVI
uNWHHo4TfVEbxBLvtJKFEOiZTM3brXsU7PtPJ9RrYVqtFFFIsdhsPeipwNhPqrKQ/D0kdAdrllPo
DUQX8LkBcHt5KzAa3gXv0238WMNpQTGh5pXHSde7M8zsXbUtgtevnvjVGnzcxX9Ruq5DQJg71bec
fnRtQcSEAg/EXNtlm+GtqZ5AkJuwpug/sPek/9hUwxugSEwTbpDKxYZOo7m80vbpiO2hCu9sSViL
VDG9SUvaRrAH3tUs8sfoGv+UQ057uUCxm7hmMdj/dgJmiyaSOOycb0MGSF3T8eTGPl+TJhbLy4cv
GKoouNs8hQfAa8XFtQKhCRk/4rxzxAPzPhAZI5qpDYjtAe57cSFvGrXvHYvRuJZ/7I9WFQV4Pubh
+S251RqqdqF3WxJ5M7rFGJueKqDkmOE2I/h8TbLYIwNGSfr+Ra/CBUyJTIA8BxeYugDXog3arbaD
d+CxBccfZVMoFKRo5aVXRD+aCnFKJG9UxeyX1QWlyPn3jpVBcUfGqLlxNJGZIYwQWFmh1tath7bF
ef+k+b/xtM9uwg6bBEcvmeLdursVwsswmWgwRjsWDGH4V0/wLESIvSnLwpSV6DXsA4aMOVewfhTF
eZuu88nq8Z13qmdcmIdMCzW7fdO9+frQPnrPHJekclwKQA0a5xaW60pR0eBKDEY5GLRZYkqfGGuO
dIK+kwsWaeehcEyYpviDFKsptx8dBS55NtCKiGN5ZFwJ4+a4RBH/eyKNPh3zRRcNmwx9Y+TyfPQm
uDSSqhnOhRyGv71uZqEecyusRt+zyvbV+wUaG204gswVcQdXOFkqZFEB0nQ+559ttbemmjwSEncb
epKK0xqxiOiusP4SZbDFkoD51s+hDSTIRofivUn4MXqKwANoRjsrCotThhprXuceRDbQIROTwjTo
nfXQ1GsQ0QSRSmwF2Zm4r4of+BDyWUnj8EUaV3pIHz1/MirsBEZtVTeNb2JlEgLduPdw1f8jf5t0
12rCox2yQdulSt2pYSJ2UrzOEj7FpUklWoaIOMAIpVmrZbENaBRu1eGMolGhs1Y5G6+3KyoHJoM5
wOfW8Z0TDNifJoBOgFyXLrA5SmtgdY0NPB461vDOATWe/yamA+ks/CM50YlqhnW0U0oxGGAX4hHy
SuDlXnh8IR8DYS+ZXtSSMPIpkTJDaK42hbiv/KQy1M3uVbAqsU1I0xRi2EgioFUqxC8H3pqwQuyv
2YBuru3o/C645ViGSS4JwpbxCSoH85snv0uVCaJpL7nrkMYrhQqAKG/mQljgQIJzlaEv09YdsVe8
RSa27lJGROmQ5mImFuOjyuC/r2dU76ZLzZRurZJuGXamknbQkfQk7bhEAmfrJ9N7xyPnRwQis2Sr
IpIJic/r4udLWorQhysRLf5SSfDCXGwEk7VlmPOtH1llMopxRyoY/Ia9TL99CQpKlEhPdIY2U954
LnbyH7Fqg6Ojr3E7s9ordPK2f60RliePyoijpbfaM8/mEFWLiM1LAW7qCsb7CKvbSxTF80Nob4jb
ZBI1u/Z/2vyFN5cPNm0K6hboYHndDJbvTmyPKecbfwEdeFkdjdI+IAid5mGP5av0HbTC7Sqn8nby
WpnhO2S56A8ssab6LHbZevRshXZ/m0270Jh1FHAyzXAVNmouJTZEvTvg7Fp2DOuCBjfLXmCHyZzB
/epQ9E6vLKMADXS81kSGBGW9R0BcYxsVZjHaafwITWPJOS6jpBYeZZjIgywR0bWbuBU4BUVM/yto
pMm+G8PxRlfDt92Ghx1C0Fqxx1FAimhkIKOyei03ovsaRLba6qlUsk/Tp8dE63G3GRkV9oWXIVdo
63lWy0+/syEPO0/ybJBTWbLRZ3M+DpWU0qpcyGtNbYFNodLH4qyUxZND5JT63qzOtVg8+uyjesuc
pcBt7AeGTOOa/A8P8I+H0Uh4l7bbTIoVUvJXbA/IR+VVvrZhqTjIUDXbChxNtO8B+rbVvAjCIMgg
mP11PQ4bZL2DCzfIjPw7dT6JMByScky5i2SGdy4xW83o7EJ6GvQT+FWx0tKcBQeYvdb8fhT5jFdS
0XO8JPuvJCwBnAUOfyRGEqyxb0ukFdHKnkbjNTJ3biHx2l0xD7QI7EfCYM55dxFj9DlLsclkSEy8
VhNqzkdY3Mp7Vq/UeWcDKA5jyrg87wPNGyH49cQjnd8NHow/a2kDnPIsOkRDWup516UJQ7MmOao2
jVAOp7pJIFziCN8kl9lC95D7vyRWKFu/67xFdItgi2VV0KF+apI5qx3Bq6Wu3aiPTaX+6JhmDWyA
VrFEwDHD1S17zKiWz2awLx68khk2i6QmHWkSbJJ3jt1mJxj3Yqs26BHZJr7mKjeDst3o0GyMtDVS
6NjZGhXTy+pJuyPjYc1acn1QU0C4YNmmCRLhGLYcV2tH+F9WMiV/uYGtRD/BkyQg+Dy3aVKvRu32
+gI6C4Q/3c2P6Qk3qv1kuAF2zFgWTayuTNJYTOLuXeBxRrMQ3gAllmO19rKtotz8DNEeTbbXTwOh
eSQWE/1ba5QdKif2XWau0Dl7T5PqEbLczpuljLDJs3yBDqfJLfS7F/wZliz7nmSVqFaBozZm+41h
+JhuT9SVNxBAJL2TeqN36D/qQ5+QTJSgNiKPojB090X+BqhjdBRXeMTkZn3xlDcUcs45Y4Nfil94
DihnYjDsIeJiLUFWiJQ92/V4vFH/cfP0gly7srzb44XkXZfKkWAWxN03YZBiWpGXtO5jvtRdv+LA
04gLotn1hP7Ld5dhZCqg86q6p4wvnL/U9DFPh95bFzLit94OmEU3ZVbjDFImjqDu7L1RmE/uhQRh
EUPnnNbGOPqEs/v15MYJF++xUl518Herw1pj9mfgaiUlQxRdAcnaurotX5nrvqrXdFPVTrdmfCfs
avo3UTXCcDWgY5GFnKbyqZSGHu9CQHHnBA7C3Q4z7zK1E1n3ZyE6XICbRY6YeNJOg2lHcZFO5LXh
OHmqjnZ7I3E5hIrI03bMmdroUwCndRFyhVOPorvsJeo9kPd8piN3xCCBbfkqPeWYg8xJTTYcNUw7
riiqKLOzIXICaf7geS0bRsGqNeraBMroPcUi+Vf3DYuLnoIFohnJFX2dFaa4ccDAdjUUtH5PpPrM
Wyz6bcoAnrJ3aaBf2wIZVRvdyx5V5dWq5FNqL3y/Lfz475VirGeSJeQlAhBKoDP13BocUGdBF/KN
uUfSCOlRs2SZoN0TYghw8tpfvUyK8zTscTauBUHfHtyWNDjwPtL3NtI0LfopgnIc0HCKqlz/jFVD
6d5qhq4dsnUzwb6VYQxdHP0Mm5mjUBPvgXDLUyQl56popm6+nCOsHAbHJVe4FK3s2Tkk/VdUaEm3
lcRHlPRVjznYNgavuLI8JUD/sioFAxO1qx1bfRgEBnwYLjCRs5tWOFsaatQAzDbS4hAZEb6ePT0g
qpPCi+Zc0LHjZ77XXxZrnwY2lcLtuJzYKZZlt+bGD+hLDYTqFefo6sbZZVTopxay72tVdZaX50Jg
CmqgluYhfL6TraqoaqzT/zVgs8cs/MgUHDxn1IKkPUhHFpaAMnmU7yGvWMDyAJ4vVNiAnSR1eoo+
CNly2UIuLOlDxaHUNysz9W2iZH3goL5tlk17uIKYf/ffqLrsuYPVwZcMrA5YqFyDhTMdtDq9I0lC
WF0QRNN0EQhJg0VXZP8N16qbJMDnRPYd1XyVzd+HB11ve4hpcTbEkdxItF8V/52aFJubcUON/12t
LAbBbV/dCbxyfiPl2sJgGez4ZF0DVv+f6//Zx0UYegA51LOHBkupn1wYKr1hggc1X+JXa4whddXi
NDXpDUAXkU8jyOC3OcJlh1lyuQrcbde9e3uFiQI40rsDqJhg3JueBguJ9GXABH9iOTILM10oe+Nv
YxSSajuV09SodtE86Anb0P/20lZ+PJ534cfiGsJVZpmOFXrB+hQrpDGxYnOrW0lN360xLLmJLRYt
THj6/wbYiRQq0YniGvd2XcptqYp8BhLRtoZORMcAj0CVvW0ibwRPASGsA/bwp3I9XIYWu6KlhYaZ
XmPKFMpq6L1t7+w3cMgCOmxlaGtQyppE2n5756GqimFQy8Hj/LgpHPa1yxmSMDJZ81anvdvG7uj6
L887Q1e/GYNMKXNAc23fQmwp6vrOphw0oyMJJntoy4fiG+9v8Yp0TLzAQBfVc0/Nh67dx83FWz7Q
pXT2wexqXdYy/wg8ckoZgrYPI2gZ+kFVf2X+biC8v9zqLm7/ISu9Y+I1z59ukuuoUK3musVzA4G/
jRvaN+k/iUuRnqbyBYXw7V32bJ+bI5GBbPwyXJURLcg2BWouEAYhzYdseTkBxemI0EFJkJcvbxJp
pjifp9ITEd8R15l9/1AKsAuQpaonyCqOEpX9oor1LBOrpwGLovtQne9JC7/c4ERpnNthH6sd7KM/
OUQp0SaOe8khVJsdY47317xNMlsCNaQKRdvB8V4H9cXivY3ybESEcjkMloBzgu+MMNdLQY6BbYZ/
ivtPrryPFIixmo3rfVL3NhF4kMtrGlPTxhPrNirC4dJ+ofTO4A56hdxvlYVB2ovM8HO75vZuu1rr
xSGmbzb7FAFOdB4EcsZq4hTHPqTFApQgbAVSnd3KR2fqlG3ewzh4nw9efSxjPKK0mZHBO/ZiPMBR
DivbHSOTPaJeuerDcC2M0JWngbw9FtCFpXI3tkdqSE5c8x0z27cJhTKHYGz1J5Fr9xl/SmTd9Hxy
pz27xsxDzYaNqLzzzbNMvCnh+VTyN+omFSjD7ijGwglOVpmTyGjhdbXSw+HfK8keZbsLOzJc/bl7
35ux5QhKWB8H8qWIuDaI61RxuQLhfSvHMXrN6pd4WsAXFOhKwhAkC32WG3POtcBeYNIW81SH2/8C
OtK5MbXdEBPB23+MXZsfQjWD4WK67qdBhxkcoSrmtp2IZSlYk4ba4vFqU/w74qv1EJASmcoendV2
UiiifJaKrznIW+VVbvrYiqsmBhmV0aZA6ZSM5QRNfLejyAQd+nmKoLjnpXEKmh3+DRPhmFmhW+Bp
t+Ft/xZwnuCrAt9+3YRNfalSjav2sxWEYXxvKOCrxRiickQm30q1oKIwVI0s6etDiLZeF6bV+bif
HxDCCTqz1wr/7KX3gqhE/7wYjR6sKSgdkTqP2dsdmcEEbzeZCnifrnyyZLsSwLYSuJ91jzyk5abQ
Ea/SqhPGEr5fOfs9Z/zluqdLBUZy7iJRiETNFAs7qS2GjjOBbMr3p/jPT2F1K1fCandK4XX+GVDr
WnsPlBE8x0MHulGvU2412ShFvryv0T/64w/qo5O+5hBopNXZdLeoGPgtqIb6NYySItNADAs1WvTp
W+i7xLPwWn96jdhO5I9ILDL/KXDu7ucRU5LtdampLKsX5bALkHaYdtw3JQpvHKNa8q+MktsL1alu
/U5OnstphxMV4VCOs6DHDyPwsmF7szFOIbKwdGHx23GHeel71RWKWUP70hl9yDJe3iWfKjLkR7A/
DsGlqXAHifP+ZdiDzjxclJMUY1i7WTOscuqTJL9DJxB7j7kQvS3G1QD8B1/rpGqJZTZ6cZGp/aGr
aHo5I109UyLX7Z4qsFfCr/lqLaroRJfjg1GhgpV7uLt3q7AacXjYJsXfCCPyGLXEbqtqJbse4B8e
uP6hUMUkgDP8ZleWoVV6ajy8K4jPgxiZyUiZYGzrvxWqjFnEkTosLmUbroHegNLaHt8z40h2e15K
3pVSzAH/S6QDR4qWnirxxhARWWEnJ4tSYzbNsI+gM8Rh//nAINFCS/QfZerLv5Esp/wTq7BI0nX2
pWW13hFeZTwYiq/Wk//BAJqIEIDzeDKF1Zka62U2J2pglTRk1FdI7apOhVWFx4bVyPHrmIp5LdZn
RM9eGZq45/NIt/6xYzp1tSgzOG8TXnu0A7bpsHiFHHVB+cXu2PkKEo1eqUIzDLydxNtC+ISNy7/0
ynH7JyPr3atalqJDxETaJ7fO+FA9zMCNhFpNyfu67KZvNauGJJ9mM8nsUhyRz8VJ2Dki5zbfMU0I
8AZviuQgHHS55kv3suIhrOGjv3grnA/c1kUyiPvjdNcs/Xs+wdtNYj7Iw0k95a5DPH/JgdacucOT
XJ1S2bXDMQyb6H5+8CzDggjtocrxBYKUzMSCYg95ucPKBtTCO3uK+ifJfSQsoo+gdoHnczwtC3W5
nVpROlDBh2s840MQUTAyyj8cMteVJVJqTFSbOka+bSydK0JqYeujcMGOf8QYvd6oPIMDCXYWcSEa
5QZmIqrcOQNQeUvjzROGMKJ41CdKyp5rs1dxVysvq/j2BrYKB+TAEI6K/P+2626jdnMFs+tVbJFP
gLymd7UL6QeChHqSLxTg+qEp/BLzbDAEzFFg8+GTnnZaWpJHla8XNeDRaH2SyS6bCtp1XZ2w7+qK
UjUjm+2XRNNd8hjRsRY+YaUZpvkEAHJ3OUSY4AuJtnWRlhFgqMEpAlmKpRP+JFeogzVjdod/NOsU
LyxABNX5L5T+xokYGs370xQ+PqLqefoJG5I0GIYxYvH3n9j3aJkjuHJ2iWJed9vE3952iBh/uWUQ
fEoOZKOfyQ6CL1xECM06KebMVRsoaIBijjILwl2FpvXZxPdVvv0cJf0vYnIFhX1ktOrU4r1QYcNb
XGTd0A5gj9RLD7uclQUUDIgvxRCiiXRELLsYcAG4ss0ss4s6XuwdLu5a+0Fm+Z1DvZrOJdWQMGLt
vXGjytjF9nzW9tsR8m99N/sOJ3GMYn2sGLLn7xCM1YObbPJ9kYsT/qGWFNx5PtCl2cuatM2Ahadh
hhNmpPUJmhxbu9ZOscMVjaSv+OR/iOPLc7hlN92TXTs2AZAwr+ZSUYS4EzXWQg9Upq/AxhID1yvy
O4vdQ5CUD3nksqMEpQJoB+wKguUgxktHCdcsyRIYT7scJRw8iK+9UT0mJmBpOMGxkK27Cbs+TSkl
q4SgC6nyZXy3U+hh80e5w8dyPzs8AULRjPV04DM6y0UjFiLE50xYc24JjNJTLqKv+xd8bU5TYznC
fpHmvkZwsQ4PhtQUcVN4aTic+GNq/Gw594Xtj1fEYyftNu49zRdINOQRJI2bMOd8T1LJmo168BZx
+lWMHxxPjYN74/GO3ze5DU5CNX6xnBO6+iY3/V9SSX/PLWlRtZrdibSODrcggvY6vRVlzogXRl1W
nBYlnb1R9LjZ5A1JL935RgjAxJtqiMbXxzy2mDVBTOGnQlltI7S/TrXUoz8b93QGIiHvxWKbnDDv
PEBjJSNyKoYLAftnm5rR95tadQ43S/y9V/eVdMhM4fFG2BqJaMDT1Mvv23/byly61QYS95BI8fvo
wSZ1qFgTE86toaC8Mtmg/gYGCDC1W68HO378hohCWoKP4CQ47zT94XSlWxpCjO1ck9i/C4zGN2rW
8CwF0wzYoXBjJXMkmFLe7SvtmGVa6qswgcdSy5vu9l+tf0hUZXT/M/SC5mOgLvVTqC+e7Dz1CxLm
M//SsV0GAbr/exYZlEnY0ElAPc1UHMSbJjQDEXjR5kjRXG/bWdxLF7G3vUHvJ/O6ZTRyEjdtRKdo
hOifLsFuGVb8NC6a1sUpomawCn3Su1xwurtCncCc7nQntwfiv8ZmpiauZX6vrqmp67aQx9ZPbjYp
mL7ceyM0OCvkxL5PpsAZbtXpPuuhtpKz9tU9VUFepL0Fqdxiwz0+e3AMJzq/Utv0o73Z10PWSIPP
L3RMNvIaevtjuVFS9oWhkQmDhIyZGMaCSuf5SboT/nRRfjN/bodPwZF3i4Cgy7MpRUXn//wk85hV
nLRzjtPINxURtahN2WOG578AxCPC2Y8tFJ1D+IcSAlI9M5mQwDQPCjGvOzVVRYI3zWai6LKnEc8o
WRtXEcyF8Dg/upPeCV2cI4v7MBBPrBzkW7SinytEmrIzf3gruK+QYApC26goC0xFn3K8lMMKprN7
GezJP6PkZy6eybdRLoXfCN6JlruRQZ8KQZ1srfMCgsoC0deC1DuLif6xBqf6suNoXoOXjfaJxrnO
CLM0XbaESjcKDqDyUgefouVuFiIa5E/TeRyc8Ix/5Y1mI5kK2whZSwS9tWeg98Ohzg6l0RYUOyWo
8wU8Y7gEa8ajNlre++mJ5mI3HjowA/DcK1oSou29+tcpegKFAIy9LlYXkhvDa94uBCdg96ZIWu2q
x9kyS76CnYXQN9uaLnTsiMZUtFHLaUOS7NIi/tLApSMh5fQAgOIhe3QGo2l4P11MLFu8fxSj5qKO
zKCT8RCmbGWUh1bTY1jO/fZKQlS4pvuAzRmxMxjTSU5Z8OwPPk31CsdiAy+E3eeWkvTAW3Wi88EH
rjZ+hlMLFB/1F0XketS7GLTLKRrNTQxcmn6l6jB8buWw4RjNEQX2J5jkc50wrGWKDKGmk+9Shm4P
Pc/M8IoJFDYpgl4I7APbZYCvdFYLOtjDD8SLpZxsdkgEh1gKogW6K+3xz9b2NAFNgLIRJiEngtqd
DPVPRl7uineg9lX+Q7KvBYZJMchUqhccz78wsJRNcKRIFJuXJqsHN2ICHAZ9YhuP34y1CTcd1Ez/
Vxpybl3av3HUYU2cwumCtSFTysQ6Hp2MYemkZ9SkZlB3xl/EQi38x34wntSm4+89NURRLl/ioh1S
hhYFHFZgFRK//Hi1NV2U75BbxEpH1578YNZ/y7QobdqgMgfbduuQ16lMNPUrXoro5dEONRef7QUm
0knv/RuNq3Lq3RmgU4x4i1u7WpxqUkJ3IWxFovWd7wA1B0w8S6xKTNLhNYzPZRQfuzegxAIkhu+8
ngsGnLUKd4oZaEJM+qELoKagvTOHygpJNbev6vffGxn7Fgjc+ymtCaQ11K2f34riEBx5HOO8fKTp
JW3Dye2RgfeU32rdYEM1+OoqR7uiW4z8haaonO+JxeHdbf+0iV09PIDnpWheMRg9qeEZWfuMoRNt
F+5LVusvNEWkalo+7rME6/mbVyaAebgjOmK2mSwKk5BBfvRLiVb0IxB7/1VSSWJ0exeNgt+9P2Dh
daJ3sHr7OohRc6ct7NjFoh2MiWaq2+N574JMZXl/zGhEiz3eWIPzyVatG1jlTMNyKVFFa0JOUIGw
Y9JdirZjoZmjwkbECna81ByVRuMPlILJq/esaTbi4+jn3aJKvkK3++n9r1HDpj8FENnwnuUY36cI
eg0B+SCMZGqZC8Fr3zkI2BYGGg5V379O/3P06KD9+aEI2zdPOKiz5LOJCgDQhvv/1rPn3tuW07XT
MeZrSvg08e1fuK9rnK3UF0X6RqK2dQHuQJ3ibgEDV1X/GOH45P5ayKLA62w6oLT+9o0XIlFZ0MNB
dsvU1lJQlDhvGwIi5OpCUpvSIYC1RFPSkc9LVYcKAB+yTrts/NW+vxMqpyL/lQqmQMXuLEI8dmCU
0Ew99zsNL99ooljZb1tVsZzI/dUkgSOahHai88JNRMSsizMRHLX7GOLdH7T4Hs7LJ+1uu/moNNH2
NEJX+XCf6bjHOcAU9pfuTJum9EGP8ENfFZv2hLDKj2TjHaGWi5I3tlpqRHMAq0PFvPjpfJ88voe2
G0Relim1BSwqn1EAUVd8T0/2t0MtrtnH5J6Wyuonf855kfeVonrpiNK5VWn7Gn6WfqIV6cpWC2Ra
vzRGiQSh9D7jIiq484v8DlnzXZomOyMBqGysOqDDvzk21j5zo6WdbpH5BGVpP8M9kwzAtZKr600B
DheoKWGHikLInC+y/bUZPtSOyKcUvjahIhsraCKFDsybK9r1HmGvZ3pZeqPqAg1AWfonMn+Fca5E
idyzwAmRkf42/NWwPOpWNYGKhwNOnhrnriciWDGm/BNS/T7Pr8T5V7VnCesnmDIJ4U8wjYz/nqk7
KI2BI3nekHZXGHyT5Tubns1dKwMJeb2w/gE8tqKhZYrhI8MurCvLR+nF8r7TqMHpspiF0Mzb4zFE
Xkd3jwgmUazw+k24lUM3W3fMqeeDc8j7RMZAEgRzwS6kN+K+F2tB0zuxQlX49kpj0d6xiaAcb4lt
U6emVo8u15qQLlTHuBwU9FP1tQu3hs/ZzqwUQPJ3/MKq63II0IP8dBnhorzheB67F35w2w74y3GO
tSm9P7jZkO4ouyQ2Pbubj1cL3xijJCkik+7ox4rZYzaWRusLqcESqQIrtzSd+WZ1tHnA/mRUpp4y
9eDbMrWysVdkZtY94yd2BkBeuIynh9Kxn9GpQaB9cAXMzqrBnanm1YH6zieTwhH3bxsASzQ3W0w8
5HjIEBRK88ox950p4qWta5qrdRoBbQnIa9G8g2hb27/+Mqwoy94byiKwoO71Y5LuzFY10jgud7UM
m/aRErQzpMFUilE3pduOQynu3sz2vlxffMSCmbxWOnZpMRUAvRfvI3z4VkW+uKcf5ZLeeReahThT
jvenjFBgAnBWFz/vZ2+kkN6a1rQUJabAFHYJXuiZNwlKKutNJFIcZMHN/E4fKeDnBfUKpchFU270
FiNOena0M74y/OVQ/IxvCC14lkQCAmsQb8P6vsAHQZgkOlPhPp6Iedu4yFztVoYAXF8K1OGQSIzO
w2KVGMvRu6KmjDayH3CCVthk05ICP+mxGxcoL9MVznWJSiqNJI5sPFNqlZ3yO7KgSezAxIg9g8ro
pHvyCzaLhpM42gNJDHy2hRH1GPpNeqGDtNGvnQGCEJs6PxI4iC+5Xw4AwJot9r/EHS0P3VzceKPl
ThSLpfG03VQzFEnODDUv4Lk9MgwcQVUFqa+iJndEfxZfEjlwyIhqcug0flq5awrDPevCUw9Q8k8q
lb4dY+ftwXx6h1enM3dtG3niRqENpjFDYrd2arZZ7e1999JB8TRf1iqMnKZVZ1uNFEupAotyL4dq
nz8PDDuJHrnAsHRNF7Li+RnYT8hINLa/DsZiTWcCZv6wHPrikr78qBjG+RLZiqrQSUFOvwBz/jOw
bwTcxF5dnmlF1Nv/WUFOsfqRtjqOIuVQIreEn3IV1J75Z11t0gDXfyy6m75dCi8s8TiwsfUNNH4P
/OsvChJ1OgCstppy8MHfuh/z4HrKT7+s2GxBdw2rxJf1C/F6mIMmici1usJPttkGKzXaDuFivZxr
f6ZpicDIT8nl2T4PZhwd8TWTmhMy22AnWLSZgQo7ZiAb1fm05Arp89tOxjlNHrI1bWnFyr+Cxv09
ie+o8WHjmCktnfd5Uu+kKavHtS/v5xLrfmsxDP5MPZzeLv29l3mKmOxQjgeDqhvWkjHkfdIBpddE
yPRUCE5SZvfynFxzk5WyabFADuJoCI/K8m5Rvmezj90368dTtxRoc+BbVXB3r3MPmjsY4/1NIhg3
0jNVzx5onVE77DmGINdYZz5JDin7CVMAKD/ulO7OQtDEPj+d2jNBnnpyRWz+/kNR3ndgE6hAlzwA
kA0JV0RNENKJafuNKe7OP23ozpnhrlJQYfEQ++4N/+XXmljp8iADGRxWmLqeGALrJJ1FrdM+aByM
crbG/IQm5niTmGypKw6iVLbOyaCye8UdDj1JxbY3BEHHIQjxf5MthGtywmrPYYAn8rHMIbPwqxky
mhFxw+htXXlsmzb8mfUG0ix0WQy+iAtNlV8/cV+s1V78RZHflifWmt2vZKOyrm+QhoJZ7reXIaEw
tIcVrqveN0LKuLWh1IFQw6UUvx3Lpe4ra5K6VKFXVCnhbVAjQuJfdOhhlmrw8djiecsGMpBpqdB7
tZmCtxLdK1PaUoi5BbobtkwPF8bhChmV7pfD6+i7O9xDUTW8AsKYGH2LaLiO9O98Jxw68Bqwj1cd
YaWD27eoyzWf8uk40AvsEpDXyIVO2vzgYCrfp1epFo7Td0Zw1+uz8v/fhgVbcu2PHOR0k+T/STxu
nTAW+muvYABrdwdaMPssKnkT932Dd+B2oBtzyEAgY/G4nQ4ICopHpDnNTQrb6fIEn2gcQtrDZD/M
h9UYPHpcMC2jhfOGPCfJC/fJdet5Gdnt5sAJ2wc0vSo4+Yvv7Ouks3doOg/k7B9Dpg8WeSe06j39
P+vFY9rYk04J8qs3wRq8Ph9+0BvEWTb8g7bpU/3Z7ztJqMkAq8cKGIy7aeGQVStPG5OiCzC4JpS1
9XSc9y37w+Am9V3PlS8DlAF7AoLepZSbBLdWCgivpYteULEkoehI3bUCKcYCUWcmnmfq0tADiUPS
a9dvfCa4L4b72vWoRpvdKcE9QPS8YofbpvDMU8A7u/bQQhTHMpR3h1x8p++z5Qzg4C2mQblGeZeu
2pE/eS3FLMtANwocRDDjzKvZPZvVwkzPRgvZ50H7fKARhbeP5poa5jjZIRaZa3USvG0lodJYb4G1
wApLXa70oCLEtGfYD3qb5DZAlmqab2Ad+x3ujDC8RinBo7DSj6r+ojvhLE07vsilZQyq4qJXsKpr
FpPjCWLV/DVhjUZwYRo2VBDuPPQRWF/vIJLVDhimoWvAumtZoaTFHQ19bfGjibtoiErEPNioz7eL
oAqdo+u/d2+kIqk7/ovLqKYg+Elcg9rS7b93rkvwXCJYCa40jZRn/bhgsdYDadq/KIo6GmL3AUca
q1GmbreMsiqphQa1xraaz09esW/malnGktNKwb/SVn/e0NLkOVt7vaJASCz2aEJTpe2CmhpAs4y1
saLk52YNnBm5vY8NCnOAU0zsTa0VMbFvBkv7Ka7FNLXVsCIcGF/hfh9fv63JQolGx3RItsixIxkq
Azu6LFK1Bymelie2jrIBf9ERnn4KQn54WSMlf0s9fGl1LPaXoQBYYmaPpmc0DJq0dxmTyBlyOSB0
Y8d1kO5CVm9N2eQFSG6sxVzp0m2LbXLPkbisNGhHbeFzuJP7iZp9GcaEx92n+f/8+M6hNnQDth3Y
cUeEkovyKofC1tAhQURdZYVdNQKtXhIPO7voW72m12VVLXiBV3N55CTTAuMB4elEyrvlcKvNEqK0
Yi+TxxxjCYbD5UBfl794yn4r1Mz8hnrKratwkgjamRPXbL9nXXUJYJ7QFEoayUxsgxwksmeMi0/6
n0Gc3KZIRbBJ3/vD8Ex4mg8ikNA+pzfkJ4607QtEZgSEXIH+pn7SHtOtmdKfkWbYfDJQ6S9vqzvQ
M4pWoriY7maCt1mydLCv6klC7iYdnhwdwruxL/vv9ZbrgM6ez2EyxKQCrkutsilMpKiu78VccMof
HbgTtDsW5i7IWUWxaxIALF+sY0pwbRvK+wUWC5iZeNTaYiMj0jPlWV7nI73EZnzOd+y5GD8s/sVX
u+eRfAmSICYhMdQx7t+loz9543IFAkELA8tfgy5CbfMWc0N6Kfut/jrc2qHJBEMSs7y1YurlGKQ6
taoWlkgG6YJstt/qFZLELa0R8tleZOy4EiRTk7bXjE8aVYK2N94s+z0tAYyZRDUf2F+rXtjz9eIs
8nvAPArQhhBuTgPvOfDTrffg3o+MF8avcMT4a5zltEThzH3QJRKMImwQFzBwGKjXN4E6D6u5eLHv
ySNu3nIIW6gg7vPThP3NPPdR/VrTmdhoIY0erNfLULRv6xcE9jn4h/n2nMFtNM1VttqTRclYoINN
z3UgveCQriVvE+nRlY5eh1xfwE9w46BCvqMGQ9Ssqyuz8UO+AUmb7hV8vxiEP330mqq0W9t4Z5uq
qdU1h3BlQLgfQn5MEXBx5McSMw+hSclr2GxZ59GNibBwcPY4x/IGPuVQKAHEuQYudNA0eqLDFuaS
1EOUX5CzEeqUYKzl/MussOwanuIchyrik5ukDGl6+DY+USQRvahuSrPlU85q794/93JD5n3/BQKz
moGFxh3vbYqZcE6FP3FIEsaP2EdxDalxHlD9xiG0vmRUPEHmgxcvcjIK4DI9Sw06ZZZ3wAy/SSuY
YTt+31glwdjcSV6/pSRyNkJV+ZPJOfZJBt4HXfMD32QYdwPfjhqJu/NUY1LQK1k2l5a3dqvT1Mov
Oko6bEzEcSZ0Oo+Of49MYZD8NMzxOL9Kq858SwPBCYdO4wIuc2PIHtIxfA3os+VIfaQvDKzcPdWb
X7hrf29YB4PYXat1H/lIEw/+9AiUC3I/9PXLNJ/tPoqUqQZ3jEZUjEz/vVnklnfjlyAeYq71/iU4
mrErffuICZ+rGfRlZLzE1Yq5M9ROVIQR3wf3dtKSrSacrmPua1gY5MdY/kaoYr/IXErvukJ4bKQH
80BL2qGogcT3x7ldsNY0gN2pKqxTZ2PUQjcCCTpoTkUYoZSYO0FUW4+cre5YPavCCs/mhU79eCqN
ow5nByyqhsawgpkxsQqOxdKMQLx+LuifXD+ABHxJHe9QQeCakxn8ZCM+RFfPfpWZtTS1Yv50GO1P
U3bq33U3tdwi82Di05mempFnLvONptvBjKDEP+1h18heSykIseA/VyDoZyEUR+rUNDcGwHg8JJ0l
/rhbJkIYhQxsaE/4YdI99bGZ5CH101fm3Ew3G9fbT9/rENbnHW4rvktK60DgI57AftS2qVUnk1C5
pJ106bTjqIuaL+Q/Xw3O22bxpNV3NzPWNIqR3OSTxIF/qxI1WgwtnYn1NactZ9YebP6GJ9fxSwhU
p1Is5QjPXBitvBkv6t0bwHxpGbajD2EUZWeiXkHfq/f1kYXRbCL7px5je6uEVfv2tT9ViHwiDnUA
3vRoFnXO//N/ao4rAWzA6/lgGcE0GdbYWymVFqSlH6ftSGKE9mToPVwz5TZvdhHmTTm3Io5FAYF8
IAbbp16vlURSlY7fFh48S8mWRDhKAliK4lLgI7Hwgf3EfSlCD5j6Q5LThr8bTBDkGpqA/6+SOaxT
howrXHXX0c0Lw7DGq0Z7YEA1K5YZ+YKSBfJ59ZUZUvfZR1hyW/eWmjoXIXQuqf4BiaMtOofnJSYb
9XBXLXvJB/7ENvdkKTDdtx2+71r9rs6Md9mJfbclgbVMY0KdkMuAyYYTvkxBHINf3Oq3m1qKs+o4
SeE7UFQoYVGtdk0lzJN7HYaM3KprwkNQXuNxyN8C990TklKhzevW9LFUy+cIHvA5fZ3WYtSXY8PE
Oh/qxzsa7Sx6tNdiEaCrduxhLpvKC0LKzO7FFxCIL3ooOY4xdVDDZRRCJ64iJJlp5xSQichJmHlr
In37yVjgWu7xc5JKo134mulL1p2+rpRL+EciFnYQxMVnx0pbuPKrr0AJo08245moZCwZRzpWyOuq
dAo1KbOOfUBnWro9gFV8pP0ftsAxws0jIfGDpkeDk4Pfs2degEJ2A7yAMTb8T3eKtf1ghj9bft9+
1AEo/m9qSAQAMsQEiUkrt07NwDD157LJcOVrf539TT/8RdDKTUjTSD9jQfPeOCfDnApiKcLDTR4s
e7UQm2MhxuueCkvOleV+2REkZZQYAxObNbRY7EJDEqDpgweOc4HqjYu26Zlf5ilFR5+R0UvHV1HE
sRhCDcossEIYM7wzLZjz8YGuWLUUZTZBQ7fpWokKtiBqPVQWrEc4Qz6ozpthahDC2sV3Sg+3wu/D
a8cp3TbyohjEeNbo4zN48+PvJHrmvZvu+wI+YH/SS73aSEjY6CN65RupWq50omXDs6Y6CshAM9LF
Rhz4L1Rc41qdkr4JEs/J8MY5Azv2uVmfpPVm9FpbTyPfy5BLWO3LSeNzU3WtsRRUwlbGIDuO5THX
AGXpQyxSwBi5Y3/CgV6Bm8lGQl0RiNhHPvXOmUjJnnk+ZJPoNKeY8sO+F9ONkc16VBkGXholSPXp
SNDGB7rMREnfbcYy2Blbl3jfJgqFY41Dzms9YdUb13q0znDEeSF3QqA/eZpMBZUAKAn5w4PGGruj
itiApI0cpa6lNv5nuYFOpr/YIDkAE6yaVQJ+rAJhiEpZ1S121IY2SzAfe3Ii/aLK3Hw7Bsn+cRaM
pF9Gho13hvwMF/Y5bS0eTo7ChvBsHe8XsdwXAFBPKA9J39hj+D473QRyy5YO6TH5sV8vLO8TwLWk
uMsGg0inrTj8O7T4b7pnBiA2e10iZekr04/S0HcdDbEI1FOViuKq2+rzoR0qTWFYcQipAxUOUkJ2
NBJS4diG1s8yPPMSXZYvU3uNHYwGDkzoOWvNa0cTF2r9d3d9gzQLazdIaS6KoOrjT/k7wQff8emd
4JrRbFmw7DiDIOthLX38vLJU7YtLwNBDHO3ExxvbAfnO3EA23zaG0VLhrMIKy5p0QENnKJdyWc9n
4RdSVB1Cq5CLV8KmxNdN7guU7OA4oMywvSH/JApHO9IAfPLogJFywq7a/vncw9MV2qQ230vcsKO9
SN9z5x5fF6AlRTR9Vw3yiNklko+BS4G/XFHOndRBGienpxFeldvcpP+hKb4cMNM4p2FBzbEJMabo
ZqgafcJnjdqSrRDcWOuxtOaqnKIMk1W5KG2w10JenSF3MBt2coOU9B5x7RMsTq5+5dV0otdiLaq4
eO+0RWPrLGrZZqfkwQTh2GuI6d/eG8N+M+s8+6efdyGr4K2Rd1BlRT8eGtXLtkpgjcLegTMf4jVK
2jS0y8KBY9b5Ne+RD46PR6gbvtFHs9PSiXYW0yJi7meIaBalrHrW1pGFXS+SFPHoWPk1i5VjVy8j
zK/Uku4eXWw4Psoa+dSJXBoaqytgoVxZofexJRanM3wTAXhV0uhxwKSlhMxeW661tAB4vNBXaGDm
1ri9j+osNFCI6lSr30x+vkzYtDkgOMhNnkcsH/IE8htPbLZcYu9PpqztS9lpkRCwkitgVvuarg67
6g78OiFXx9ke49PZRyQJlghVVrZQB4+e4ALxCos8wVKRyermWBRIVh0rfW1kjzw1Sa7Ekqz/s8sb
s8E3c/I+RoSnEh/ARSk+wxpAYI5hnMfsSUnQRWOkUskDMBXmSJTBAess6WHNMu4bdrEewGboiJuI
bjrDgWxOaL54I3y0Txk+r70mxFe6UcGMF/vZL+AZE41nhmQaQGyfPy7oFRjoniyoC9RMyEDyxZdU
1qEqLZLmNoSxc3GxLbaKUTfDwii6Aax32G+YuVYdOvz/7zz8vLP88buEQ4F3FulwbRSFiNogTjwl
z6lC7vaoX9dcH+WR+Kue/htNI2G/oLkPH86KqQlvW6reyZErIGVSSNJYPFsvGgkITqO6KCkYzIwZ
EE2CA4zHR81G+aPZyYcHTFV0OlXlbS4jB6mlq286eVii/a55cI2MDwxd4WA1vmJA8/dd9Ma9ZsJH
sW0FLOWZddVzlHcDU8UlwM3M4II1uYjEPcBKTJTcGJrbifYfbsanpispqmLC1/w/FeeWfxWErF/Z
pZzUCZ7k6jfWTI+krVHz6OV2vH+oGWMZchMGg9IuaVGjm/KWs5+FROhjeq0UNCZeE071H9tZW3lm
6GVu9lItyvukxj13eSzKENwZcAd/C/sRYqFIrwuJsLOvSQs/RXtTzBfemsQuysJLOobRm4thO1qY
OOJ4kUTU+OjLyvMjKpYt1WT96uT4Cx+larbzARkdr9UNF3QKyRRKtBjLsuMJ7FfZdWkuOdAwRpxC
3chkRpS0pExlf5UwrMOkTenEcOC5SKdVuYlZC0WDerUUMkZWM5J9/mbQlXonq/Y6iCf0nFWCF3WO
W68Auc4iqW4rRtMhic1fp6bZY4t7ZND+FefWs93I0wuCaaA/sgJlH2g7fr8MqfHaKD4FJh1pRLjM
xoEpbp6slKPYNh5b5wJPhmVsCuRVTadC1xDI9CrC2sNWJKL2QAI28p6PB7m9o4Rf0POtIiArBw8z
6KA/qX6Nb14WLy4yOz/7lX6lM3cpTUos0cfgv76O3r+j5jWZE4nzYsxx4mbdB/uJLrMl++AdGPOz
ckk3n7MrWlVG3kKYEwoKNmNHuheGPcLkqyl4q8RoafAFMeatHLAHmLOP7hHjhHisfmFiCuG9volw
Xj7u4EyAeYHAYaMglnR1E4dsmttgZXTS6RNn5kh4m6a+gueL3SH39yE53k4qpA9CoDy3lO+v/tF7
3LR8kPM/CH+A70YWgFJIbjp+ffsVoVAsY1l3878Uwxf5QFtWZcNYkSNNgMBqJMPeuc+ZqTKrKeA9
5v4MIftbaSRCCcBVRBg62ncuYodKgearxqs9WthZk2ds/T47rccQ0fYRKMhWQKqTSswn/QXBhUrQ
3JRhGMFtnx9crTR1RKCTqA/tAXZxbTw0RpPbIVaOjB5ea9jXN94BbyAlMFLxLn8BQuSSYHhmw159
k7kIBDDPDzrP8rOq4rLATBHZAJpj1d8Q3TYXPL3EtY3bCCFdu7RfRBluGtQVjE/ISCKLDkjOEJBg
WtLMxJeMprKuwQ2BIY5FCI17ekgLcD1II0pUYTuI+CoGMr4kNlVTEVtMRPtO0vCWzzdRWVfbrxo2
hIuEHqG1G+PAUqgYnRRHdcun9qCBgwv2PDaEExhKYlmBuIjxwVMI2pLJmuFbAFiG+vM26DL/+oo2
CUr5ZG+9tFJLustgEbArOuVhRrQrvZfbZdxgyl7/I+Uktmm2Baij+5BDIdl6SIn9faMhVqC2bpZo
QplNjrHCEUozXz+kOWCYShQxDZdVXeLzUb371DEE7KU4vsx5SuTyOaj4H+lM3wv8W9h2IYvSsO4e
Wg8K7sT3o2EwptK735PEtu7/hoHak4CZGZXSoAAnDP/xFsEXsnuW5I8+jGMwR304elbFmrp8i9F0
jecgRRFP6p2QIe+zkCnJn4iHFcKZvMcVVWmBrUxoZUasvON/L2Hzw+SZbGKdL9p5vRjIPEEwjvci
mDbAABYlvbWkoNP8AQyb6FtUGuA5QAv8qEvkAjFHM/7Src2KYht1h1J15SPWcjjiBDYzAkHaW6p0
8Rum67GSYGbzLh7MM5OvfP5Tf9JJtS1iltduPDC6FjgXKGDch7CQ1zwETnoQaoetf79sTnYRBKm1
IM+Px8xWtxDsmg3eGNrQSdtlg/w/3Mcx2qEl+KUOHZ6nrKKDoFXbD9XUQaLQLxmU+A+TUth9GGq6
71mYLI5qzRQeHKm6zkkdjhPzVUZ6nWr1KdefiVPFBV8zjvfsFGTgGqgGCdJ9rzzvsgzMDfjJAge0
VIiu2KuA1WkdrLRXwzKdv2GCGDzaG4BR+of5PZJYMKiHKVQPvgFP4dxSJ5XgVydz5w5WzULMpEpV
l1E/CELXCLUqlRYFJIUwF87yl8/mKDIxv1rcavjpB4OWDu9mCW9ouuyBwME/qRNYs8CTyZUKuHTA
svZr7Ia2MBlknJtbrbl2bi1Vm8+8ofPo1ud3KH5JVF99uz8gtCfALfoLZ30KJLtTi12suvH8LpJH
gJ9iqmoi+2uu/w7bmoP3clU8p1YfdsYxyQwz9BPwMIySbvBBfnawArv16Y3c/Z3tEhqLvV2qswDQ
dFuplV8JDl3rv9nXDO+iBuuP4qDGXK82UK6pOMzuqKaNKONFX6h6Jq7hUpH9S9ikM05Q728SNtBd
yjZrR9/Rfl1PfzV8jgukHB8BvxokdC7+HtRGftQwFPl6pSQdSxJ+H1+MfFTVcrbRdKFCZUTkjRVJ
UW+ogek64kgYAg13eaJHYJ3MbB0gD9PLTyB63fFr4ap08uWVHJyPk76NqNBplzM77Pu09cA+Rby9
3M2eZZS9IMDETUZ0ZiqftgJeCCsRgvSn600H0nr7le7B8ZWHu55gE7wxZiJVBV+z2PB6u0SIujYT
aqPqjfFgD2UvzBjUS0cytWXvZHcZuioAxTVUNexwSq/eo8EqylUpP5H1FPmaQWkLxOkit6lrpGTu
n4ck9gucexzYj4Lk7j22wRejpvI8XT671wC+F2Awpf2/hXD41BLqfA9DdRBne9qKk3dZ8wmmDgxN
02TCjwHbaE4gfRveIGiHJjuNl6oEIiDjFNqehTtLfq2R4wdnOR/1iuVB9GOLOy0goYQDnRU/NkOM
vuH8dwZxbodhsGUCyP0spfQCbknRaJSjT9xkkx5dKYvBWqBX5e2xYZE4neMnpLZt91axvhAXgvbp
h1GRtTifyGWKBVl7AGgZJCBlouuIPwgFXpeS5EHRRNXzF9c4UONYIXxZyI7nodgQiOh6S284B+jW
wVWqSrG22Zpuq0cpdn8wOGzYY/6iEiG3gXQr4I0FIzk3GaxemgKWRROliS81S+KH0OTBYxDlKzKP
yjkOH4Oi5389hMPl9Q8ayOvYOR7MTDXPMgYbM8J4qDrKFg9TBOrIHaS4EPLYY00tI9rtbfxE089t
1X6HWFBaedToFIsb51z9n5QrEF0mFXSKCei610NblEzYDYJhGmhcHxhe0Ph9s1aF/JV1/yY82JkB
MGAO1a4SaVIqfJLUDSOQY3yVHhYTLiflzcQbI/C4qFyc+lmWCy0+FQuD7y9rQiQXhyERApAW2KwP
36EdikxLqlzXkKDJv9WRCepIVo00v8GdltymAA3+1bYqTs89iXuvHtQFa0dxOZVApuVV9ZldfEQj
wfHzpYKD9KF2W00cFiV12g443mQDBKbOOt82yi5UrX74h7IN8FMIwCmpi8xT0Mdq0r99muXEnpq8
yMuFEHLKRpjYYnHccHhQ8tNVG9JtrugsQNTlarEYndZKmjxP6U/LbVl8er11YxGmK2GJvU+f2DyO
UCMCBwhUF8nIf4kqEO95SNiauLp0lvqGHxE4f4z2v5Gryy6LjR86YRbizSBBRMHHfES5OT2Oq3n2
LEadL+qpjZYsVGS9DHzrg+qnR+oc9TCTULGB34i9MMOBKW7kqsqBPx8sSHTNAdmRhvIPMbbkMUKw
MAnD0XPTweasTPiupJEXDc9nTG7DK3oedvfaFfG0s9ouU0LWoMYt0B/CPjh46u1c6AQibaHMzjAo
4DUxvFMzr07pEOyIjXvh+cNZIM1NJbMeGl+Bpz4JMt247W/hHsVw7cMZDLY/dFyGl0MWnQwME3dj
W5h4jXS17TwfkqdpbLbDypEWbsgpBfgu1smHcwIZ5zwyrhYYqem3g14iVOdlPtQuudMcUXJk3Mnj
2K+A3twuiZ4jTQXzedrFiw7pdueF+EKf/h2HR+hmVYK/D7RCs7ztUrqXS1F/5EAY0eFijsERq33i
qns5zy6JdIMIyrwl3j0VzUqEfXnVPClsPzXtBGXeCk66WrJxaEsiwq42HpXTSCRgEk0lom6BGCUv
WGHvzNSk5zAlPn9K81I6d62fMZa858BewGQrLRy3JJTUSlFyROrBtLfnhzGY6VvHatc7NdQcGmuS
UWIltcVBMHIWkEeakUNMcqN03PDUngHD/q9QMdjVNpUQqu2WLn7hhwj3K0xx+CzTLShP3E7jIsjb
MOk0Jt5zjTMVbXFL8mxgprqZB4+hOR3WDboSgGJXVawOA7LmtTOjOT/HqkuUZD0gkUuzY0q0v3io
paCkN4PfpgJO4E4JcSe6P53s6u7hzzH6ZThiY+BKL8Dc0n14RvzJNEPiPy6iZQ7TGngeDpeMviGV
1ZVO3c4dcSfZhl8oT5y1iMfDteFFr8v1v0C8FEQ5WDcqJNpqtzWq6WOeQEwn5NK4995ruA5cTbU4
d/EK3Ui1lYEMUgxyTKmcMdkFflydEojecZ1kL1Z3VMHpfLhMmM6av35mTD0W49lXZ4gdjtDk+cTE
AW+j+ezUA8SqjT3BQCWPeQYBPA9ZGLPes6+qeIme5NyRGTv8b2q5dRtBh9V1lSRD+2vX/Qd8aJTY
kakWlyeYSOerTyGP9l57x7S7v5xROLFBUo7B6WXYiQoGP/K9LDXiVO0C6dyicNVWEzX1Fa9neykf
dJ+ByKq3zbBr26512/trSOakMyEVoNIwU5VcU3pYENYQawdARoAHXDWutkjgRDhZvG5/zRPRfs9W
Shqo4FlSoXmga3uq0Pu/0yWQKXikWPbBa+KBkXvG9sZ+DARpERnqP1tQ/ap1u1OBLPanrQ5EfJTi
/PSHrmwhlLrB6B7B89Ibc2Su+emK3uXng0qnvVm8DMCF+Ghw9zWJVx5FhPl330OhRfJPw4zJpbNU
+M98G5F2WIK3RY9PC4JRQkTI0zNnK30TxFW9YSkQ99hzCCzwGQhmt2qbl8q6N4UVpPTc14+VdVGx
vOTVQLIefaCRuXL7uDTrHBu2YFau6meJNPzCrie3zbXgk2y9tjtNS5ku7o2NOE80hblU2i+GAccD
C5IrCZH+yZ2NtFD9KAn0hyCyZ2SXXtZbvdJczSgwZGER8M9m+oZrnniqtP3edfE8l1ADA2czWfrs
4EqGkKFCwGnr/xSJxUOSivWfNm864t6eTjFQYA+fmDo3maiPWMkaF7wjpitRmvK6J+aypbNm8+e4
Ns5IxwVOohOSKv6b/Dd99VuMB7FI81TU9sFIbabreiHVCJ0HuSVQuGUFi/CsvsyjXBiRdMqtqFzn
s2OxOWAKKj1aYw3Wt62odJep4yHyhTSLNbkkPD9xSNmDnWX4CENGe7pvQ+KpoGDoltbUgVMFcX10
UzjkFGO6c2nxiwVNLVvib4zgj1KyKAZacobsfEcOTg0k8rqyD+00EE0SJ3dUxNKlqjjx1L8xZKSV
WIlSlyE6dn1Yor+162Eg+mv5T84+VxFfDbne+YLEUAVk4kK/vy9J4drcGiwpklZuuITlIDI8QIUe
TtPb0JtkdYL7E46Ce77MDB0t7n+l1+WVZ7G12XNx25CIFh4I0Xwlqh55HqbwdCPV6vF8e2iLGYdo
jNvFgR+XGWbPVQBzWSkhpoMbHF4R5+qNjbnojwjhzPh4sLGX5b4bCjJNQgYFGrts9RbaWwt2TgnU
/x3fwWF4EWMpM2mN2gmmoD5wY4qhPo0CeQglWOX5LDapcPKqwoALloqjfE7B5K5suNRv62NU43rs
xSQ2iyayfRLPYmB738L3Dtk5WzaVwXQbzOlyMWyB26AzXHkj/C9IrmtbnXSljEfVbMLvNVCZSFmV
VXmSa7wm8xQUSLSQtdKKxWE8EsyN4YtfRPat9DaJ3lch/rawimef/8jOiCu+T3uATQN7/beXkatb
KGHLKyXggAuM7klC39DLcS3DKczHHn0mI5I0CN++x9+T7CJ2d8GHlTRv1MZpDX9UNXnvVhZe3BHY
dRcGDuoojljnlhHf2IpYL2zC71VCZusbGtULd4rS8dFed6OHZ77Cj76fGuEpipw8pULCH2rFbGc1
3CUz3rMSpeLBKbL/8TrIdRNWFpZuzCUsVh2fvzBCf/YCpGoXBL5tiT8Hz1OVaEYIkCHKkC7XsVfZ
xiebeRPOC6xM9PfODHO+Q4sYPXr3LRZ/HtAeo2FF7+lVGRp6YSIcq8pzXkJNp9c/9teltgqjmt9W
4jgQlEBPpaUqABX/ywkKWZOQBS5rYk8ulnQFxpb31Pgll6bfOKyhic8fMMUnBC7rcSQm6XSOO9Xs
mdWUW5ssNO6M9SF3thHoL8QHzZYB0+tlsDuDcTqCQlVt+2WHMDAMZKLSq2Ht37J9yGm5yr8aim/6
WYH3aoyK21d/OmEEAhCrBkh8MdaLBB5D8WULW2iNiqWbjXnyuIY/dLSQr0nUUIBTtD+FxPeaI5lu
ovFJBB0b8WAE08R9GaPUZkfUjJyt0U+Ws2WyKlCewPV87l0YWr72Dxz56bXdw3I6rWr7ZICiCkcp
NRio5RZf5K4rBmVIhPR5Cv5fCtJh0tV5Tc+Q+J2Le5pv1MNK2cjKo1BzGXkjDht0yn5R+iL4v+6n
LvpjhDYtkTxMR0TdnRVxmopd0T94OIGimOyGltsAQcnSUFOCfzUtUxTuZ2l5MJoJ8+plxvzLnbd4
vwtNlWidcBk/XwXs7rauZhT3YT3p1JV8AAQMP7CJZpXG/xACQE+50bx1IICAd7l5mQfKha6DhPqO
a0+5SSOeRT9aWU/Y0P8bmSWiWdXE6w5GdIVRKJPrhOrWF0c2zi4FsfMSLUhSKhMSjgZfLp1Ex/50
kFq2825P7eN0C9SU5Yx8uNehPOdUaAwiCMj5VCOvVpWocw3/0OHFBfQGRAQG674JxJvTh6dUus/l
Wwu4VjdYTftf4NQocIqGVwKPW2QANiY+X5OLmmAn4OjPxlx4by8DPv+WdNF31dlG45k6L/DH3Riw
zMy6KebL0dtlaFb7w6oPqO9QM1TR81cot2bfUlPUbTBH7Dza/MHsg/pcrIdRyHs+cbLEy4BOoMUi
vOA4JGUNvXv/HQZqfEKADYElXmdRqbpwfdggU07DD7YtL/miLUMpLHGdOQJ7AgPGaWGrb268s56H
9SwjQnMFJTSKhdhOO34OtqdrnNOg3SYiGD3V6V6w1XrmYvE7antXC1vFkUhKr0CDpO/OC/QA1/PS
/iDAkqkf5v79X0xhlrHj7aDohzP+413d5Vkj+2oyy2aXoGFSWhj1pIAfZKa73YGlYhOaJmYahBaS
j52ON5QwJdeArSuOt4TkH7GukeoCPOKHPjujY9I3p6IEPETTapdnfLgtZoVaFU6PFLcJJjYkJytK
Inbq5lGlMb12MixI56L3Oowe/ObmipG2JOUgjCe4Wcg61p6m1OdG4NQsdUA2mTyMogp9BzXPOZAo
2j43AjITgZEpgXZkgUGaEXOgk1lwlAwDPlvhDB90wCGOmRJnGTrOZwHOlUgz0fkejhHZYnrzDZIP
EOg9uqj0SpU1M1paGgHldNbmAbFI6MYgNxk4hr1DH4C8++QYlEyQne9z8R3pz7SQSakxm+1IZ/7P
AkrrGf3oEJIWzIFNDGMS6Brn6hgcXN4gIV6CGMwRaorM3R7NU3HlTvHMVw2D95LXnxplOI5pneA6
c36vgo8IYNzEu0KJhdhz3gcVJh9fhkzkjrApXNjYqLjFeGvyV4Msgy3zPpUoQGtshAn7tnXYc9gK
K9k8eb7M2CvOeXH3COKy4yoCqF/oh7JG8tsNgohouB/clvFGn4NhOy5f+gSVbNrMMkiREoKFiRN8
Xq+sBk4ItSeeLGWoY5Cagj9DwtmpwKYnFeo/+dBixm0q3Qqie9xZGV680bLvWp+8P2MEzedUafZD
maweMvLSM54K+jiDCr1Mr+/TpLBS9cEYgmgxwJJ/CKp8JwxHkksDae6BMYFKqiCRmXhEp3KWBK+7
XySJHPsKdpl1bItsBJxn4/xrYWFTTYdcZYe83qfcEZAdV68J9iRzga4S+kW32hG9pJ4/GaHJYIU+
Hiim9W/aBw8jzhQjtmGS2Vq9xsoQNAOBcdqaxcO8xzfhz3FSAVeSZIsOGivsOMhQ3kLgC3WL56oJ
YPaiXJ3MVrsJtB3NNTyHRTkp2NuOifj6Ebw+TTSzMM5GuYwQs2Rqenc8T1yfnaoJiOPy93VvfbcG
xPDiIUmdR4fGQ/pSv/bKXlOLjY85mON4T8QevxYOYxuTuEc6AR+4epw6mBxUQvkEcCsv78xLptgt
HrBkE5mPVdtkBmuYEeuzFe6GKPYC6uOYeE2MzyFF/Lq14KA+myOsFUDO5jPOnKR6QiRZCpJqq7uI
fPCOZtqwzYJPGW6j3/o7eOBGEa350AM1fn0rD/DtWQvqlBNhCvoJh68mnEGCmcN7snSDGMLf+Wvj
PSFe7nGOrqxb67GgzIslaOnlhJm7hzTdqlp9kl2JMcXfez/cVLMH1nHV3VBgbo/W7mphTbm/mQO3
NPG6vDYrZH7lu/zkx/aTYaq2HsZTTH7Lao+z3Gb2UIVzh4PLJni+mjCG03kA1OPeZuz5r2B81is1
3LhuxbEpFLVomB1EY3BMW9Vl8cPyyB4zXRFS6j0ja62prWbWEqitzrunEe1sP7GYNJo6+MJHTFR7
g/5K5JppcZjLDyLu8X4tim8+rQfKd8n5iJX+yFLeF0MLAz5Jf0U0rbbYjxfEQEbluZSeT1D19xWm
IuyvnMkDkPs62PNcSotsb4Z6C19b38lFOhC5F5jVZn/0/aPAQMk24WmzbVZTr7W/55n6IL3PA01s
PObRq4rNMUbL1xpFIwU+k5TYP7jDEm2pDzLcnoTcplhidVlDCAHw0FPBVyd+8R97x7AthgkQDDg8
FmXhTaobNotoj8kvOKlbkR4VBRY/vCe+M2/pYoFuFpfq5MEXoCK9v3n+psQVjRlxrhTXXNQt6RQS
eE54G9zXDUcRM+K41XdHwUV6aqBFFUZgLmiLfYTVBmoZg3R4LZI8DFsTlUAS03iRI/mA8vSrzRNI
vazwe7DdjHBqvD4VPmXsX+Jwrgj4gSEE/Ch3pme8ObpwPIfpdnawkh086kM+v95CAMtRdwAM7fka
AZ3abonNOmdrbk12DErPZOi0VJ0gFnNQ5mZ6i5asZJA15xCSrE2SUPLOjgv3zbNLFw3udxVB6Hc3
17lFZKphPVGrbWjgp3C/qvWksjoRcjxNMCusp0bGdE/Ug4+J/YwpeqMSaR+M60CejaSk/Vs6JC39
wgjDw2puGoqYUVhwwqWzUV23JMeZvXqA8tXVu4RcUZ0JekK9ERkpftK3gnbu7K1WQ3WzUeQ9VyTk
c0pveAI2tOotiSO5nSY6AlPCyXqjfdzE66qD8Qk5u5sMRJjZREnHbie3rn7C76tCOPm3vkbh22lA
gro11h8Joldk87ziTWCyxp/oon+v64bOg1YVHX5s7mAPCEDolaRqKL5TxikPObAhTt7OM8BFCRqO
MMJ9VN6Xxhgn9wZuAGXpFyjkseQNDpt36vytkxAPEnHDlUOpFm5KgfL33Z82jAA00fc0TwhWovMN
7wkFElGlvKwCJHquwCcvzJYixYlHp99zFXoIFIeQ2ei6xteN4PD+znJdNsISp3yEVTlU0zjqM+GA
BzKc3d5qvngEvI29hcW9/L5V+poWtwHa/n5VZnK53OY+u/m4T80CAKdxllkVcX0Ks9HNF/VKn1fH
vIyrO/5QiIc8J0FSHWg/i2q76RbJCMoQieqUVwVLc12H83RCS8IxytzZQrCva3MrVgkKZDgYiRhq
wva5zNxiA/kaXhFfv+w6mHFvDrm2fc58JSk1+1R8ndIT97b7XiOdYdgGfQSDa6WZBH6ECUKLHLTK
0Lf/6v2OKQ2Io/XyDaw3MLFHqPRGq0Kw7PDtKtkO+9W5RM4L6ND3Cwuto6CFZ6S43VodMybYSND5
G3wzTzLknHKqwBdmhrVxQX96JutvvvSvNPlBqKDmpN/6g36G0L/UXA0aa6BdUnp7Nv03rWfFGZNs
0sMOUlBAsx1TYGFT4oqg3ncXcBYM+SKoU5dNXyBzT/uauYNQIdE/KChGIFjeB7421tpAp1wWcUPe
R7Nem0QCOlqjTdp+HMaMNg1yMNKy9Qvh7p5eHo1bchPWm2SzpXu/3dBohQQov9eO9+B2pAs24pTF
CjQT3AuvqbBZd1ioig78sbi9Ufp5l6c64lrvilyUnBjZL+pSBNannKzGPd2Qx7Yn2AWFQTPh4UmZ
u+xQ34ZeWUDIdP/4XSEteVjqyuhrrjcaBPc6MYvV+Y8nf1IUQfoFb1LAyaxQ2uYQYDRyqiggJRjj
XBDuf632RWvOMV8sAemxNfL3MZKCJ2xRZGW23Fiu1xatyAgvCEPOvId84+E+m9lbUOSH27FRMmzh
NbKLGL/GPj+jh5IMOF2Az21GA2GHdWTUbGOrA5QsOt/byBEf1BbrY7IXt9vCtESI3wFRrhDNKWx4
35i7ama3yaB5i+wi3awys7rzcpT1gzj+bWWnW4uJ+hQsU1YvCyEMLOJhRTiQI7/Y30U3fF2ZPWnU
puVGMDcU9E6t01TBt4bbNvqIBDMAc9BK0udsnnTtvedEOKwUuc1zUtJpk2LyLbG/uOL1qLGjiwNN
mCrX+PHuPtm4nC8nyenlH5zcef5D03mlSJkH3VpMMuS1TmNded4TAPmd/naRb6dFp2QjuImyPZJM
ok8HS3q2irfLV9+x4asySl7DNnyr3UU1SLGoD3D8PxouFcqYkWZwE1QR2nfpDzk2a8LH0T71YO0S
b4kJ9XbxTXpTs+S2Zigpd9ptnKaG/TYiYHfHG/S67S+UOc0qghV7eIDdOggcEgaagWfw2uSmn6Nr
Zx7megoH49V72CJ/YWo/L9HNeuaZd+q+O71uMXlT3V67g2st6rlt2owhdgm3cyUulZbKlDHA2HfU
hkBNiWDx1WjwCWQEQWnU/qifpGsb4d/mg4gsD3LQ6Ue5gCiG4Xgjl1kpZfRd1MyKugwi+D2eD7Mj
BHlnOPrR5308WW/VvvJmSg3yIp1wK3JByBoWfLiQAjOmKjsrjZC926kwULBLtutWexKIbXuxu64Z
odVpA7/SP1KzA7XXpfAkzkKjxNdB2txSClQofD6Dq5YWDbANuKsscF4i8bWhKinAGmpd02plrOJv
+pzDDF6hdqDdGH8Bf/hjic4QQxnESp66x2IcicC8+LB0ho/1XQ5dh4E7Iivak+Iiug1lQ8MnGnaM
yHuQroQCxyPz1rSYkYNYQoK4Nc5NZjYmqTZqMFduedwzdC6jHPYR2bLJuXl3PbZ7rV4uBrZetm1Z
w6zmdM5iYchI80d4CLw7i5GkImFnI3Wo+uVmFMymPWenKwJwwI59PLO95R1Iypvcw870vPPl0Qze
g95B+FOEkHHFSBs5l1LFoDoU5U9kr8w9mcXkBH9g/lmpbGFz9zPj2Ap6/yJP+9uF5yjyvL0cVkc2
HUKpxl9fkLMkeX0KHgp/Q/wh5Ga70a6w4aHiYXNnfXb0i/brd5+Lj1LmxRlD9Y/my+TesvzIFM6t
bAHI4rOF+2anU8CTLNPQcbOWsdVoTUqI0E98RO2o7PPmENEQjk1pwKaem7WFniZrVGnRuAxWDnbD
uPP+TW7x00Jls56roSK0RbII+SWbgrL8ufde23c82fpPdFXTZzPvO9gt8ZJ65b4p75bmvjdXUlW7
wBFmWgrD9r7NL1/9hW9J57X2jiMxPkaCC36aP+698KFUz2CTXG16tCzbwce14Uh13wKqb2tHAeFD
UGyTHVzwZdF8sdJPtdSR4SowVrhvO/FrPFKVjTNldC66Ms5WJnEo3rglZ6i6PKVYOXm7Ps1AM9Jo
BFx9z3LMnj5KhcCyjMRimO/c2NJLn1DmdU9143iXYru0Ll/vohEPBrdJ0DryiDzi3NWWfWZ5YhER
DZMb8cs6D6Agap3E60vE0dlBoNWERMBnoI1dD+1zosUp34JfSpxGdtd7z3ukcthVU33DRCCk4Z/j
JdLy7WQEyWJQsS6TW1NL4YbmRXpiE75AqGuudEz8NKNXtBU8WY0hdB18I8+rcNh3WBii9uGw78hC
h7hqZ2pupbpm0TFXmexPjUiNE4HoPGv4If5beD2oy2T8xGlqYASMrcoPYQ4IfyI5lN4RVhE2IZve
oq5sONnAfPpO++N/V69oJmKNc+F+ZiUpl0QNa/151ObzHLjCKl5Ctn08HkLhtKxKkA0sFmmC9cNe
XUvLfk+CJmfm6k+WNIC921Jhh8K6Sh00uGWnvPu9tLhc15lnWsWGw9oj/dLTjiCqraY0e6U7U0Gn
jBGzMvT5i3WFAng5kKOrgb3vOoYeZTb+Z76z4NwI1dWMA84QLb6BfFKIIuzBXwJWEVHSIVWW4kpx
/tsvOwB+xNKSNvc5fdo31lvL1pNpUF9VN7XwsOYvW8DH584sdCl74JBFuxgcjFxwhBzAPH72anIe
Wcuh8H4SUXpPeDdXT35+/3Ov9juhK2b4h7RL30YmWfqAR0FYplB5ivtgdAMAHnNdKzwpxkbIMV9v
JLDkyPgUbztCy4NkRO9oNuTExeYk8rF/TDbDFbKD+jy7q3TlnK33qI/6hXFn6n8Q65CjrvwgfuUJ
GcWsj99wJi1pFjtjeU9TzTcOksPxIpsS1eSgiPsY5BtCpU1iKHct8YKeu0ZkAnkGszcJa2SbWtYU
qIrQD5KoQ+UMzBEbXIDfTVbzhet4M65LDqp02RbDOM+TZqD602FOOKVL17KC7EaYRxMN0regcsLq
uq0aFsWv7NRIGCvAuk5wgaVnMFlS6BwbrM6qvQ4P5d6pEM92xaa5v5ZdfF5Q0Q0LP+mtfUVpD+Qn
E8s1wPu/fho9udW8r8nlJj18Sc6Uu6iqU2k3jdbCgKnKUULG6mupRZpLsgMa5VrnkmyzQBVMqqKR
6pPTRlC1AVG86KF+irlY8emk9HAMDQ4hjYalUz79GM5C3EgUd6DkaVLXrDZLISV6oWsaCR5bICu4
wjOoCIBW6QCUjGu9ncoRfKJokmTjItAYtzlAwGsJ8dxvZSRrf9cHfvHqibe/2xh+H/mF2QQfKtpb
MbS6RtPcQXlpFGbmZxplgQwBgdAYfH3QpNa+tnwo4D27qXE6YVpYixc1q4oiZmFMgvsQe2zP/7ka
r3hWv/ozBQtDGThR6ySqSQpbOlt8o0E8akIC7vkWTN/k5SL8VSeJT8oiaFBT+bvM9lNh+IFb0GRq
bw+frMuu6FM9GKpFd7H/e4I/zEm8rFiLYx12F+5wXcuIL5A6tRAUSOkNjVWAZiHOCBd+VyGsbuXw
gr2tHS576umuinWN7S5WyMnhsXDWFPYC1Jq99QkThhn1WCeHdDlVswdGPKI8AbTIovXZM7R8myf5
QQMsl/YRJ8L3gIWAd1LVYp9YrxNd9tkhS6sLqWPtT5Kb/we/C/onGZY512+SI7dResZ+uSIsLEm1
czumWJmcTczqY1IagEyIwJ4EOtgkD0FowZEKHKRrW51IQU9VHxeWGLgnGbQkwYvpF0f+Nnyn84KI
krvA2PAZ3aFQloKw9H9r7lqZ0r7ES5NPWr+iuINpuDYtodUQGl11tLuYA4ePgddBf4WjaMKTJ+uL
9Or4ixoa+zsMs2Vu9AXljZ9R3uCRlioH2I8GmaCZ8/+3AnAMh6vxUF4TZNkb5xT0jO1mOss78SJE
TtIkRPPOBt2fCFN4611MYFaFxopj/W+3OZ8tCW7Mveq5FsuS1pDZ4FQkPVofzqDkFLc6Ct7fQ3iY
vaP1cpsIrPuZoIjlGx+EqOT+7cZ55EGIDrh+v4q4389IDn8F7oRJ5V9sKLi0Ym1OzNqkkfPLpOlz
lKFKCU4/NK+jd/L06muMH264fxLv6PJd5SVFY1HLKgBeSevbmSsghv11eHftqjabh5aQ9Q/soUBh
kmaE9WwqvQovLdqXn+14oNcL/ep++PiGv+NXePlupFBpbGuRs2N9emWx7F6iO3EQPwXML7++s5l5
e3Ta+6BEEx0OLIHKdrEKELj3S1CEeR+cCa+ZXOp0ewgQmos/vc8LAYE5ZRycshlncS/3Bd+YHIvr
c5X7Jj6Lzf9Ens9qeYBxhYTpzMyNUlvccCoW3aZwjGZuD9rRDBJrgk2A6q3/V+Z0T9RjE1TTV3tb
EVPoRZvPsblO+UnIzGo9Gfxfo01DC6hp0qzCvFtKouM6bVqbPLW4AO6TBxpGzPFTUaOqci86LPFh
az4Or8aasYJpBwn18OWv3RQl4ufkq81o4vh+hLGsAwVOPXUOWDqu0aTfv/vI3I9BtQ0zMA9fY9pY
A0wmwwEyj/4yncbQwToDz0ahucJ4VojNZtGVzxBZKpXHdmbtn9gqLBToEDQguI2xyVt8xj2uKzCG
vQJzPXFt6Jr1h2RtMhGsRH74RQlL29Y0ntyujnuj2LBjdkZoBM2Kaz9byXU5FJT6DbVFGRjKPYQe
5EGogv5KA1uPWTwFoflxHdSpObjXdGkCrQNGDkndgliytTCtLcZhKheBlMIcf6FfH9Wzj3rvEJlF
cZMk9Td6zO3/gFEw1lHHpMu8tZPuH9icS0Ma5+Ps3Udf7Q6yLzo1y2FE29xhGcRGYx7NHlC7rE8u
k81F0NKrgYuLjBBISpccEoLllVe1RWEcmVNrDJEitEiMwzAYPAtm08Kv9J4N760ykp0juJArdsLI
6VHmG8xMVjHb4A4BPzyk3fVr5CqApRTk/tkqTMuRFaMhJGFBUbwMLKFVU3O3VQP3k2sg53Wn1htL
RJqth7gJXEzRB7XrgNo1AjpkeXPlheXyL0jfid5MJwOqSS/dLr7hopzgnjq0hjcfuniGL099y97z
vfDkCTW9tld2I6+r1zpT3Xr1hfvw2jjAGJrt4qwXRBYEQAOEukio+0g6jSl5xe1fqmsGGAm3npHi
xx/QOiP/jfldnlY2DgIxFI+iqkbZuy38NFyTwPV9GcMVorXGgYhv1XQn8yYm/VgSaYvfe47fRh8f
9hPZrBX2/baUW9jrleLRQIWWS1QZU0v/YX0Pxn3+mpt0yAblcJ6xuY7tV/WoCn/SwAZGaZA6YUKI
x4O3sJuaKhHwT1WoBK2GHld21wkGwqxTMQeVenw0clL/W/jYD6mxTSWbWQ73FREMwAzW0WOObiND
CJ99XnnS6/UOQXY1ctHwlib06qQDVdL4/ovpEQOIdKK8b3za+6ZOeCy9sMB/p+fl06580pxn9P1K
DFe83DMJSMWGW+heWWA/WHMnJSYfGRAbuLAwYwDMBlR50yxm3tBEBxiiRfh3W28st1PLvKv640+j
EIqK3vGXdEFhmdQFaEp4mGTzm4bIHWdVLtgorBOG4N7IH06wpZcBSk3VWM/ng7gLpRC8MvJQm2lx
aJQe35JqR4NDql39FnreOzVPnc/FeQEJbxTZ5qIicdbnXxJIS7BmXIs4HGPF4EfLTeOU+ViSyOM0
2ss2JzM0SVSDJvfETnlh9q5EM8EWi+6X0WCx8+WULMPsnnQh3oGfWpqluMh0hGUI4CxfETVPVIoG
XYVB/gWTq6td/1D+bPR8MdXtwuQsjui/D0VIV2M9QyyEbFVrchPPpxNv3g367vv/FqaD/U0n8N6h
OiektyKlv/GMCVJMD6lEutxAvUAT2X/lTD2rBlQo4MPbgbAHbdxKQyiZLJRiN+8ARVICP+gFCOqM
iKG+q0CoNH17nvmYoStAXahWjJnUc1V9L0pHBYwYvgFw+hB8Z2psCGVLz0RUISLOrY3z1K0dcI82
0R/UaWXl5GI6jriZAppZwnaAIkkADbGhHWYIdHkyOXZnsdfgLSgsm2fQ/iJeGMydR0WvzVRPEOoe
JA63xqouUkjCJ/MUL3VF354imR3uV9/FLwD+IKSaatFYCih4WhLUjrfgscPL5J9KZ3VcHugB8OWI
wufohGrIIdcEvoZmCPJusUin//k6ye8u4Z+Q89ack3w8aJzEoXGgLFIYfvMcwQUCFcPdjFLyH7ap
Zh3l5Q9xqeMio7w5zgXr1TMmTHtgyuuPmujtv1L6cIqFHopEmkJk8+JdvNAFhgqL3G43tHdwpsmm
j8e+ZPKS4HxlesF5dn9+tHE4rToGIHytQjM64RX52ZmFHjA5P4ivl3wObEd+mUNjT2vaWOFgq48w
jkSKe8rTgRbd9R8RMTJGvKAIlBci2cEjv+RgjjoECqmvsNvSo2B30tUi+9ZsDhiktOQJJwLkVRa9
zFhTE1rDfnUiRVYkaLRt4ik+RXknTPTM65GghwMrbDCCibhnGF0u2zlr2HpWsjdWx4CRYXoyarGN
k/VfWZVUb+rlHupzdNihApt78faCKD7HOaG4ykxZbpDRzAbO3t0MRumPytBWyR3RvaNHxgwXmbpI
xDqXcfv09m2cRHL08Gd3XHJi/9ewo8CDVdtF6AnpFUkBXaQSrILajubQ6+lncrCENjGpCrQyfY0t
Mfjg4c+SiQJ/7TGXW7n5/RvbpMbhgZiqoAfknntEhivYM+l5WNHKCWBpd/PydC7e4MaiF8pRgE4C
o7w2Mjdz088+pDT+eQt619YtqXa3BNuUj1n2M0rd6xa3eXfWJ7qvXuiduAdhVdmYDikSidXPAOtg
1RjyJctzsU5cmrSsSGcyCzyMR8/8QKntqC7etGWfd9za7khWQHLqQRQImGdsxLUHp/gs4pPAQzT8
xcu8OpF5dQAHYMnKQyh45pkHTZRAjr+PgaG1mRHY1Caejo7A61T6TxVpH+C+lPtUj4na18367Ny+
BF8lztOOdobECPdG5S3q5U+JGLwVlHESgi7m+kAAl/RIWu5uc0+Ok/itaZFQ/pkE3MRYYLBQ0Shm
ZgPjxXbQtXcER4Vy+2vjcNlYRLOkusmLyASUR+IuZh4xYSpfeBHg3mllqEudtgx55cu94wjVvcba
GmZif3OfMSHDueWIiOBrstwfa91UROeVDQWXR9h5mbpeTm4OcmwtIe7xNObN0FsUKc9cQrn1a1+w
uQ6LVTUR/zKqAr35GVvctllejmNVUDX/zWzd9E4dPS1sGScPUHG9ATljdatmv7gjRfJACNNXbi6A
LFazog5B1fZ9uGJYRjPxbCWD066Pv4vpJNMcKKIZelN1bKqj7jbJbMqJix3sfzwcAucn+nxjp8kt
d2dwJfnhsKfqUEkPvCNSIWKJP7t3zr08RElJQEJAIHpEZGO5i1s6I5+50SLwItuDv5JimbW0nJNL
5PgJrWrjo808Dz64Smene6ncgEuSWuP6Rl/8mY2kuQdj1+xIp1IafjJVN06VR/qmPs7sF7Rlx2oz
E+7y42wChRl2NhYQetRfX38egqPKoTEH/iNKgK+DfQ1iTF4vI5jUUflJrDMRM7souTmCueRyg4eP
DdA9ky1AWCim0lmq9LudDAvdWs4Oq7DBgok07szFC19V4xa2HGiFnoUccpXGw0IbQWP2LkDKyWXt
tXK3RLc2Re6BxqlnXa9K8+QeBzQyibWJwkjC1HcyRax70g3/mA7aT0jM7KMsYAVRtRIIcylpxTHw
qhGcRdYXoWPSKFJfl35Ue0PzMmBZKEUJ2ulxx1FbF5ASmygqaeQZjHaYjzcuAIidUP2W4TDC/i98
roX7EcybD4/l0Sin/j/u5SqAb1edw0nAIoHZSWEen9FCZvJtKMDEuxlFI0UuxBY2fXngce9NKlwk
hfyuUoaMHHxcTQ/rihr4VkrlMHob/C3qSmTE3A98+lYY7v2NcpHiN44muzH8PPfmjpwnjP4Jh+Kj
TTcKj9r63RP93z8h+dXtTgnxL8EMf/6w9EptYTOuxE0Nx+LMUlMWSNL3ni11BOz2rFl7es1mwbN5
Qk3cyNMSALZBa1hDS6NHP4oH2S+GdYz492W62l7O9qtZXnKoBUus2Q9vlRYl/nSTgFJnp29ZZ8sF
MeoJZ3shIzYe5N/W9+/ZOSFssnJDfndFlKCGPAVG7R0597+zrkJ7gYSY2+3wZs02qF5qXL8HK/UW
z8GaJdMZUhLBRvVVRnNqMW6Id7cMz4mMJ/4LcOAQxE1Ci/DueYcoMOBEbZErD7lmIQl31USUstTI
hPVOzBNSU04dlJ5sCohb5ekOOATh7SS0z9UrH4WslU7pO3P6eC99ji5siscp41mrqHSjNgWl5ljC
lwU6Z8LYLlouo/b7mdmiqNVqe3L4qG4YcLKzMuUlnrcP+skcp5ovyms6C2BxSK3G+b62feDv86g2
R2IoAwYuS1EVcH3PDzb3EQBCju2KaZcFgxN0srdSaH6ADThPM/QuTFQ5lbLD3KUTolFQryQYF9RO
0X7JIle3qKkjSiSoCpE7gZmLPvzeQ6JenT1gZmlrzGDwi/C7ZVUBhM0NUHptL9RonHRsdWUgbP06
vcqZDhEa40iek8kF8ntyU8uIrzhdd315v72aMgP6T0TLtWPfm40N60SSYVzpae7pMiZVYE4wUglL
o70r8X89pAOE7qAUKo7VhX/lcD4OxwyUodVCf3CAsh21GuLM9MIT/MvIwrLvfOSJ+cQyH5OSBTs2
oyCxWEis/D4P0Wla/ul8nCltDoSvsWs3GF7X6pmJifujNC/JWo75u+DOLLqCzI0C+asbFEGJivbB
rfpZ0iEpvntbeQUKTc3EEYTGxZHFeTViD08yFIYZKqXq1vHzrpoBWNE+HbkbJMLiI0EV/i95qSng
iQHADrsrgBbWNe8n9lrnz1liER6SKPQ+dWjhRV1L4Q3Q7fWm1XNjSkZCpC54nd7xgLygqV6Fa84K
ARYXeQhqDLrvz/M7dByFdvCHQMSCMaFdE0npUU5FVraKMkbPJsBQEXCRnJIcUuQE2Vn9QdWHc4/X
bt+sSU/mCLP+HpFE80Qak2SM7kqRzTHX5Pgib+k+PpMY0p2QZi8741T/YmLd7LEaGoyQcLVLkxwG
YUWgSQtA420u1R6JJhO09ihpMvvnWOzEWvfMDGe7W8Dt7+60LaJPY4hUz5lzpzbkbudcZY5zu9bE
AL4CIEBs2FzV9OEdkFkZJGIhz7hDjTdfXn0i8i6lD/UqB+xvx1z0wbei5B9UZQf5HXR72dLhKjXk
gVwJ9yI47s9BU5xZTiROPM1LNpRXItVFiUCJs0dsFxQYWgkzq4TeuyCiC8SuSv8dps7Zs6iiinA4
0+1ib20D52u78TY+vnvSVo9awK7Sg+X7hCdYgkKt9wUXFc6OJLiF96aB5B2CG5Nh0SLU147ycO/e
6MKQYkvx9DxO7BKKz1VNOiHRztNWm/My/QtPrPXpYfUDpOl0E+FGSnKqdhOq8rTRnkVGQdrz9+98
cGyvLzEemN/44JBzKRay3lm5MiMRSAsCJkvf1KYIaiee27ZxNAwSIG2HXmt3QPqdJKTNpBy4vaJ7
yKTdEoYH8JQfi6hCLpmKU1c62TRy05onGZEjEzEoZws/M94loSdeVjoEjCHqobGE6cxF1gAGI4Xb
QK3MuR1zyX+m+v3EA0kFuqG3cZ71EL2WIj29nD1AY99iJlFjZGv5lidMZTD+3r/bCb1Pd6CgSrhH
9faQg1/UyRKODVDWeLowtsu2qd3Wl+v6xGfiIzd/dLmu1wmfV6LKiXZL6ZXWwtvummBb/jNiv9Wn
d5j6cm0OYbMuO9ysBVqU+dIkmqNqb+IdD+1TvXexjhAZXEQoKQk5wbdidpC7pKqo8oblUa/HsMlM
0oNPJjmWk1UfbiMvIwzTWkTq2kloOe92FRGtaAw4POEKuCb6jzBf8JwxKFw2hs6U9l3OxaI5f8NB
UHUCMoUzTkWZ+7zZUX+nl/5xNKEwT344oBsu/ZcE5nsNzXAgEvOns8GB9dZjFld03RoEDIhTVWFm
OhBRjwvk+TmGtObhgjaUS2FQAqe9dMokJ6Yv6NSg0DOEY9nJEFzujHkhUEPTMeaGxVt9b9AVhnoQ
NF4iHrj+3IN58fIjBGGp29ph9/D0fz0GVamPfdQzHLDsDJ0lrHLzvGDdqccx03yOY822insIci0B
Q3k1nY+/MbUa7XV7R1iwLcwzFl6vXj1ba8QnIgucBQAIV6mKz8GeslxjOGOWmJrB4EJ6WjQcgK4v
uSoCFrKOD+5EpiRDRbJDyx+8r6w/YvNNp+UysOZS/HDLAoC98qp8+siFsOVqlYZ0fRI9i3OX1xNV
e9oaa5Kubt7mAVrX3U39bXDK5oA6k6yNbHi39/l0Ls1H7zVJkWXnCmoz+wYNZs5sxV3JXR0UIY6G
kQ37sHrnR1lyrUKa13ZBH0FFYGrDmcXOmXHs9XWM7n8r77fZiXt4Vyo/ujNtPHKLwVa+faPTzY3Z
Hn/RejPNc8myI3PT8QTu+zaNbtrE7srSK374krokTMUeVBrB9zGlBINFr/PQuECWv8/efdYwZY7L
sDJTlth4GQ3zJRU27V56u5ZcVKaTpeAA/zgYC+ArQZ/l7sQm2LSqbWju6+/d/i0eewqG5YHINgGj
KyVeLMILXf2qbcP+AiKmrOk8odJwQk9AkqGWRvuxF9sZ7tIdJqh3dn5dUZUJS9iBdpJI4dm8WiUb
9XZlK7gAajxokSzj0ga3uUxiker3cOn3RRZhob5xxWzT4OLMj6R5HiiZuv8jQCY/GYh+Id5md4HC
NNjdWIW/spbB2N1WasAEuEWB7GVnqZEVVRPIXH9XKEVa0cK+44DYkqy0CD4oOR4ZZZbQaRLln0jL
zU7ZFuoIFXhxRZUYeu+Owl5iaI/GzqPfyKKx8CfZq+qnNnnkxrb82h+mOkY1kKgM5S0TZiHG12Gr
0OT6+Gk9B7t27qZUwsQJj9xWXPuedTEKiT46qBXralucwb16n3NRG5pK0CKmmVS9V7WVMmlDAujb
jaggEkI9M0d+FkH7SEkWWaxBASUNt1B1Mo7OmoG1FW9y3Yc0tIDdLDAALJQNpdfr50oMiAkr2T/E
oe1JdIOaKO6lzaz4VXpQaqpdD5tAHCOF/uQGPHiQvcYeoxrXGRVz9hk6r3uu/gYnRvCwyempaSfE
iAUtPZY+KxXiE6jUYnmvsID4dkUcSFax5P3E10Am1MVxXsafkS5xIIEnpEqFd9bzQh1ht6RirVvR
+LzViEUtmCwDfvdeuWDqsOHYyb7k8+5KucqPbY0Zxq4sGU1nBXOXZD1e88O7sH80lHF7D9BX7cFr
ClyL+8+SjFUrYqqSfHNHN1kxUaCn4eazE7IrfLhddBIkYFOr3tMPTk8FnmJvDjURcfuj9CxOu8sS
usgcAuS/xv60uFtHJ5Y6Lok0L8plXai7j2HEZdcqeOrf2Fgw+3/T15peCB7KU/quN2tMyHZsdKJv
gO4OzBW4u0DYe04x2R/CiAb6EeD5mx7Brbl4RxkFIlw7Z/YWeodIeJkgJOTjxL49qnSpqNCLrYwm
YeIBCcU38Iv4BxRnqHBd13H9v1zAP6h0DntoKcurHlXZFlgFw7mghRAwTMeDPIRvADqyj/ey9P1l
TOlLWu7kEP09sFquU8+OZOqVM9iIlRztNMEFIL76jBsu9fMH9hC5TySfda/y7LqzzodKMgRC7Nab
CDY+zs3WsWkvxN4PqICDrrQFayHD/umK7WjeLPQQr6QL5pkjG+ZI01LRQxfKamXRBN5amlzV9yIr
HPS4u62PYszBXvTryg5OqiXPL0UlOpli6aXb1eawui0hvPEO/UhqA3IJM1nh0Fs47AMVcfhwoBsC
W2iXUGqPeIbDgKoyrcSFjGwk/OLa3omgMDNe8LnVl/0bss38yKqzDEXKsm43AMfOZ5EB8Mddk/1R
GGEuoQpq5u5xVkp9fcr61w95yqSQd67jY4KeCR0ALAHXt/8mzhtIX3MrUu9PM30XwZs3J8dJlBBX
diU2Wbl9ZqUeoLN2pCgI0n8ugVwOjdC3w4cnDEL040MkBZGqHLURpc4ZXqfYBQZdLs3RYqWKFEzM
Az2OUvMia1ETm2byMFqvKnpTENOPZ+hbuT5txVcH21l2xVUPkIBNKKG1ashDfjKOXihOd6XpCfEL
MwHyVkDNAGBRwtsgqrkM0qYp2gXTQsU5chXGXl6WOz5zCsxGuUasSvFql8kxeFZ7c1vA6MMN+qQm
hHuM3mXQWYDWrgBptDIXYtFpgK0XAkS/UsYhvpI4+ZIpVAe/GZHEi/1NVuOWd6jMWTeWz8a1epnE
N0Ks2m3qfdag9nVw80oNzelqCP/vu4J21gTEXpdICFgR5fmQ1swx1X//MZOftLIE9nznVLyt0BxQ
dMvoflyAC+KiV8LiCYrvN/M5+gRY/imvg+U6XyYUPJhSmoWb77JIBcxmD1G+MHmg4ZoXNPV98nf3
PhIIgWoBcB6jC0lRgEkf8Bx1Rifd3u1R+s4QidT1koA3kiCJ94x2hxOh+q+q63CwHafTAeJrbXkO
pZT64JMJ4ZDQhfcYDeACrjFI9Ddmcu92Z2BNd2s1qYkASNraI7Uqsuo8BdWfisyK3AdFkwFbuQIK
3pOLgWFSXi1vEtFNw4EEVmdGmZVMZKkS7uRbdP1XGLG3A9sFHgXJOvyEduC3FcZldGHQ0ruHMHiM
L3GxjOKvgxstzpy8QgGSErunuvQGxGK6okk77141/Eit2PU2bp2LQN8eYbpk7bjnYq9skY2R3V/B
OSyNA/iaLbLUjLS5AaIBDq0b/zJLx4JIlsLG/woA7FhS5VUvqnp5BAPN+Uko7dQpX7gEbrcKg56n
HuVby4qLaXpZRHtSSKnTbSyf1zgnFEf9pi5NFWRhK6ze/XTop3TMkgHJ/jg2x0pia2JePEid5Coc
Lga4JxSHup6/GlvJuQaMqN7+tABqoxVA1XQ8pN6plmQkGOdcTUUC9/fAauHB+g/3GL4Km8lE11mx
KPani2L9htjAyqqPeu4gy0JI1VgGK+berzXWLifhFE/WSdJSkxP7yb9qeUokSlyC24drBp46ZG9J
MMdSs5jtqdVy67tReh32ytgYK+XyOC4EpVAve1lXQGz1Andlz0DVnzE3e78TexMOdI0iV+ztpsPG
prkpqQeV2vCXZrdZkPEBf8ghmjlGU1WYmyuaAdrkEPG+4/+7UMmFA0cMdpP9rwYOKEwsoWihZQME
3SNE8N29f0PLzNuzX3WOO5GnUz2cEvfa6zRlBR75TtQkD7eaKUgmqTBfjSUl7t+25P0C4tUJVWVi
DURXSgF+82AuSdFvjuiHhXSzAjRFHdGuAG/pupIG9aX4aVdwqLYVW48syjkQ+uftpCfvMp6JvwUg
z8IPCBeDtseo6TOMSgoxiZuEr+zyeSeuOtccGc0ysR0XwBZ/RLFcvXrtT1UNxPCGkJIGqZPtSFFM
sinajWQ8I3JZIjUznaSh+Hz5Sv6ZUAmihmyv7NxqP+a+WxjvrnNl4uaObQtH1b1qs3SjugioLr0X
kwCrlFl3k2foIQJUeBwr410vbYu+RdWIO6K1udZr7jiFS+EslXefe0QE7FO9op9KyiVMtpXBQ9q3
KrG+oSSk166Uk6+PdlymkSSPQm+7KlBQh8znr8/p+pF38iW7wDvIBa57IUxe2P5+//TJNEMdBEt2
ybs6uiRJ++UX3mawaJa+JCubRPbznlGjaRMD6pawBe/4Yz+9CoAmi6aOfaCujK7+Qwgw4KhE47bs
5gbMKEaY2cXF9OiKmUcHPPqsULDPefx7Jzm+P5+R2zZtM4DQKvP1GQwETeOdRIKowy41CFCb33uV
3MNdrWegpbL5z8qofbuI88MtQHF+UksnSQE555pi+IquNsRaEvL2r44fSXYNLSAmJz4VKUWo83EU
B63WgOzhC8di+Fn4zhiuD97p/MCYHNaDbsoSCtuhROa+SCbKABqPpKXFkwQrc6qfVZNQE5lDF3Hf
khfpMke3xDDRmIombauLb+s963GYint3RwGLBS+g7od9dBC12qawYgmb/oE5p8u5Vn61q3mqYV28
9FCwp9yjK09j6Yc0On84FPR97XCNrzKC+3iegGRs2UmX8BQu8/D2FSNpBYNCrknQgWT2nMpLlAxa
QJnirEpfotFKsvq1b7+OoXAmW2uApaHd3VSyLFClv4rrzhnpCpIAU/JuU8HejOpTAkhZoUEZ3jDe
2usmgeHvwcEXSJ4jzAr5f4VDJh61vPq9VXavnVvLh6drZdNQw1VyE8nTcQrTTV0CRcnHdrunIJuM
a97YnO+Rz3qn2I7GCPzrZDr2hBUlwRWiTrFP2QQx+DBsihbkxOpr+X8E/U3WAGstwOFAI0ALxrRa
jVuT28GeJjpZNcuEn9Ody6MWlY9ySY22qZCq0tviSCtKd9SxDRFZ9qeUovsGu7AIN5LHGUi9eIfA
4qoWgQLb4XPfMhaiTuMRVAJSSJFAAmNrSusHXLrp56OvNc3Ut0Pbj4qQVaE4Hn9w5GmlprqB9yk7
unkMpjLBI9LVLqHMFCTQttzSipJfInnS9hqkooWKHyPwmQYU4pFNhzTZNZAfVDV5IfwGPBkKmVcb
1ayRMKxD4C9DFFQQGnWJQ3RmEQlys14HbbxxH1n2YlUNnlbTImLO8kXA+VeVN0wYvtwBoqOtlfym
yXi2ZXTEVZWlHxA5TujXGfegzMT/S/HpDD+AT1fvgMtcVKUrSZhx1/vmqAKSTU6W4unm5m5B1twR
PKmFuHAaia4PF587rwvWY3UkvyxYfCGA+O0mURoniSAG5ZRAfgVZAQjMIoSQxEBLUAKmF+0NmDUW
mlY3KJbwci8+XKCM9hqHq6/0QzExxnsKH3e/CZbXFzCwFVYdc+71/ibnkcOHkOOImhq/BSpy8IVr
UNqJE6gb/8ooEh4rXlXUAaprHjDfIHLGqZ8P6sbuBSLO3zdi5ppDpCNOntnunqUztM7+++HwiXXj
pEuFMhlP71piKYFNMEVdwDbrp4llsNwCLB9Jm0NCRnuUqET1JiyrRARlBHwWOqY2j5Xpzou4Obny
fH+a0izkUd0wWcfcYPFp4YpKk/2tM3j77sbDjx1reABjNwg+SK+zFELKzD6nCdjoL7UdtFeth9+D
ADAUGaU/mzinMPcqDgVtBFQoz1AVXvVvq4Lnt5M3Pnu9INCxZe5zuUWe9gTkU3giuZntEKqV8Jd8
wKqP8PB4tJaj2KvxUNSuluOQBy4y9jasw5mz6xQFk/FW4d3LX6Z/N7Nz66hozFz0To719r8q5Y2Z
1V4cRZlIIizePGulfrDFkT2FbhpKxLQMnQZMwGAlU/V0OCcrY+goKlX1gDAWIQ2hYW+7ybD05G57
yK87ctNKKi8EFxlPN7RTM0lIc8Zp49vesyAAxRJSVxUMonN5FtNAeqYCY9omJDmQb+Llgp4cqGDG
MjkVDDcWu7b4rx5wox/X8iT42XXxeZZKmJJoMIDCYfesb3Hs91y4xHQbmvTVdwOb895ilehyqRQ6
ycQkm02bQ/kIe8Zjid6fdSej3O3eQPWpYQS02MU0BfanJtKvxuW2DxM3w148UkbwpBRN6+JrzDy4
kSExyNrTHx5lrKOWf/zLBKxsFOXcvIZ2L97/82EwrAAke7TJiLh+9wbmfVv0tVPohoCtPIolrzZR
Zsu4zS8Q/Au5EnWdA42ppb4fwwMias6G0Rbo3Dhr1rvwaCmdhxrSHnSSmVi4IEA/jzOtwjVcnyu8
tkdYEyiyqyGYE4pUQn9oEi2BZ2f1St8ArUcYDbq+0Mfsu9p6Hc9CoK0cWB9Ag3CSZ6ATS4DbtSGN
RsPSvqsicRyoti9iEjSZzfJU1oqGZi60GMaweBZS3+xl9uzoyihS/Vt+DGLWI65TUxcSdyLmD72k
f9fWZTopzcpZeH6nwhiiIbP3dUJF3Qxhb1Zf1VyVdgbtbD6UVu4eKALThK2GnxLrcZaEBccrP9a2
Q2vslBpfgny+cxzIEd4AVpINR3hwbAILnnbCc3fCkUPNJYiMUF4ZLMZo0uD7nGKY5U2nuoyxXr5V
v67Ubj8I1Y4M9NwaBPPYnMbhivYduQNySicBnbzIfYrQladrDyPsUwiC5RpZ6xrgUd2JuZjSS6/u
TLwZqZ+Dqo39mokLgNWuNQdoQem3aDpPK4Ub+9TUoG8jY5E6ggVBaY1HxhhiODLPsMUTfJexoLPy
AJ0V542MxGlqq9N+IcJDBvy29LGgdevQYKJkExkF5jHJ2AtTQ7rT8RR08FgE+PGRAZELb0HVq61e
NCj15nBlGd1jNTn427bhGooO2R9pjFJKPOSAvcx5J650INw6SBU5/lETkvxj8RKWv7DlmXQcV06o
bEAASpPKKbbanheebs3z7v+580W0lx0deVL2W03L83xXxK2Ar60VPYtOz6mpIpJbnWKbvrnsEt0J
ttgHzy44BfM2ljjCf3Rn8MaATf8jBYV24u6O9kcgkUZjOsst6V5oCTAkEfk4Iozo4Mt7Xe7o7JUQ
xSoGrfQOW1JjyclRvu90BlI/WgN/BjSN0VPK1HIMjvnCrX/H+t3fXsX9vb41d7Iz9/7EiTjIdO3A
6e1nVhZKQmyQaOp7LdOK/vqMPYVhUDq+TVt+LtFyzs6eTBOpBUwNdJwd0fElcadMr097rOsPlDRl
yIwPMTwL82fJOI+Poi3er3gjySGtAlFgy4AoKJu3b0juYLeMDc1M1adATHR8C938I1HDbZ2hwLvT
AFF7w6Hptz9xJuy+uX/55LiBvRXbfZ2DAGSC8PmuuFOWPrQxXlevexPJ/Exz41eg4xfspcFWspbg
Jh+OjIbcsxOJ92nFYN3L8xBMUYijQVn18Oriw6+ghWgJxO3MAEv41VSnnA02WQAyfVyn9evIQYZT
pBkXzru6n89I52WnWLYkAOboNuuDCd6xOzgK4mdyFXrMAkvp/DXwsCtp1VcYGLjWw9tIgtzLE9bS
Gbmt5QIYXyb3BYMJMTegjpi5wRGHcbkRhVb5BHfZvtmY1rZ+1knv6YxBWpt78wap/ERFy4XShpAZ
5KwK00uYdrKsYv0k+DRdENlJJ4DckHr4DdFaNDykQV4NMHqo9aBtH375vYZl4yhIvnTRlLjsnylO
HR8yq6Dl2L1q7v6LfGGv5PCa5TVEkUDBx4SDk+CbMDfI0ZsdG/B+u6z9c3I5n+E6MfWsf0eakDdF
2OZn+jDVTbq4nYyOSWHBiicdiYdEgTRMU/FpUgcJt+ldX0nS0NHFRnlk5jebnb2mTl/3GdIprtF8
BYXmPO6uxoKOaUBt+4jroyBV6qv+FbhTgMbCPOPFXUI70bDiyCl4ZkVrAuVO3k9Q3PiE/IJwIyib
7OlLa+LjmC/pIIRVV0u7FwypF5Zpo61iFa+SeSBKRL04tP3UKUGtzT1m9ZX9ovjt+sqKHMyHr7hO
LS0qnwoQuAYaMakkXmaoCApTq4HvwMRypRWq6j2f0P2oSXQNz9dgiQej2ospzUjId+R/ZuU8S7cs
sZ9R9RWU8/71JIIVvMNuvyBZQlQBOvZcgn0tLL5nPWlTUvIfA1WW0mKw6zKvAiJ6Bgbsz8pCUkn8
UfkAufYz/kK767hcyQaT64XSnxTVjoOONxbzDyQ6Bi9J7q6LD7Fc3/0AX2O+Gteb42i5hOm68BYG
YLVNauP41ZSzjLp/PmvaNcKMJ+gHO4iXO3kDzZteId7LeK6IkZGeC2N8DjbFZsHHJxwzrBPbnTDr
dF1xhuE/r8hEaIWZYOKdR2KAqGEQ16zbUHbywbY3e4LmOCldIGgMZwvnbLWe4korf6I8QpSN5gep
Ksqa5FDWE9ZiivbTTi0EXLadvQCLWUP5ENzCAlA/v1PmasekwOGyXPaJ72SjXzu1wA/swvcl8oy7
ooO3SdDLqUK3TuUY3dY5jkyRD5U7xw64089Fw8yg8uSb3gQ90ThDKnYCGkIbIyEvEghoNjtZwJkM
zf45xM3zk0exK/Zc6DpHl3RxMW2Tr8L/ysqaA5zJfYJSW6Lj/1ij4+IJU2Irc4BuanirkHQYW1wG
qisDQSg+aZ8KVlgz6yRGIy9A42MTpcd5+LNmsMr/g59XSuakDBwR2+jruGNeWnlB7yavgN5IflhI
ACiWnqKRCdWZ/afmT6CPBWWg0c/68PfMvjvXnUKgJr/9b7+ueSmIvJB4eDcYgCC+KN/Yddja3KSE
xhA3te5iB1vuI2WcFkDt8VGoChq2IYI+HPPLww60iZUsID250yZjJWf9Irbr9wIFCjDcz8ML9WYa
dUZJigvQrqO44Ym0hsZGLBTAG/1UmXhN5oPxTUN9ezXxpUe5Di+aFop9R5XlcUia+tQw55MiQ1h1
M0ZgyEbALe4UHYi9r/eymInCFTVao836gkVtwaIIcD1EGTjqBvCAqJzxlRaCcInM7c1w4ZwMpzgu
9m2Czy7NlmBWy6I0nTPowPyloTnxVqciy6Yo9gd3lBn2STIL3Sh5U7Bmk8zjqGlfWfxwB0p6Ha+1
JSdCypCZDNZw9vpBGnx4LK4NiNCh/VTGY36va3rRCwM8N4HMCkR31ySJBV5SPUmyEFic3PP7gw1w
9OLVBCA5mVhFZ0zcO2YK2cN49E7KtFVkj2cwYI8kSKw5pGfiMrNlUGXUl+fgBFco4pXJlBssZwfh
yjG0H8MZI6434GvMu1WmUS0dUrL5uxvMhO2he4Ib3LnW+FzaiTIyidgX3W8i5DNfFlgTkUVNVcLt
5h+s3kr1Nt8ZRLloKBgSoAXZ1yIXLym3a/gBC1odU9kyXFC/VTNiGlCQ16x+IinVjMulNGLCJmmD
LX4CFny5ZkZ7u0ov9XKNR0AoOh6tR1fFWHPDB8+3Lq9WzgUzHv9eRrc7zxEXeFCzo5o+nEFe1HMR
JL7jAr3WToy/G4R0QT7EjugJo38wULjXOHpthq9byJ+UzPtr9F+8qivzNKAfXfYhTs/kySu7f5+n
ZbXkKUTQl/kiHX1L3r72X58+A7uGN8MFEZEoZadXCJoJ31wlmu5n9GL7RnhM3J+KYl7ohDeyueOq
SouGnNU3HfaErgoCYvMqJTbWVvRFT9cMSzTTxZz7BEgA584eujf62nWqqrWzCBE43QtFdRXpzHvb
v1P+InUl5Cr5jM7uHY6w+RqGEMFo2eLl2Lyntd98DBrR6J3ywENn7FWl5SgH48/JID48xgpXF9Y/
mgGdkK756xfMIxyph9in1UW8d8QE7+Kd5yHXCSoBxzEGlw1iDB9X5y5aEUdqL3uB5GVgtFVumD2D
ulu5J2uxnWgrCfQi+JJOPfWaDG0pHk5Dy3zcDvXrrCNgNeGpP2AdgHnSyZo6pZIdvVzLhY1p9kIt
7cMUzWicrOMMwjTYHEU2Dv/B8TDyedPMdy+Y6t5qFj7nuqU1yQ03Ht+koQjFUjzpt0QWwldTgMZo
aXi8MBKmByQaS66ejOsKpDJMUHKMOQNrkANXfyml62h2HNCDEA5ldDmsOdtZ8FYgwsXWxVLN18Fm
+W75ZqLpOsb7+y7Dw5gBkQhXOBPnwQbLrTnk+cCM9SSPM8YtGWZ7jpWHKygYkb5b3eOxmW0PpaP7
iW+zF2PnfSnWWIt1zF7As22enJD75XcTCeWBEe5mYW6fIU0cEn7hdX7hkJ4YwHxXd353WiiZ5P/+
mwqV3OfoMv9x/rKlOyGpGyDs+4VbN5DcoNCp178dgaZd/1sAB86716Y/GM51Vxvohvu4MS8XdbiB
fxWIf8ENvNDibRd3UzoIdlsLFngVj2cpLFI8z09aXPTnxovcdR6U/7hYE/HNJS78dmBXUsC9PhBG
V64NewJKlQBP/kYMRHDIeeNogPmSCvFVLV6kH1JngcENTfW1BGxHFdtp6T2m4FGLkgibnpAC7hMK
v/OUnEkRDK64Nu84UwBiZL0QFqu37+fAFe5AsG2s2nnTBo8eKeNq0rKuFCAl/Ro+EGq5vOakPtVW
MN2Lu8HjYKNXANEv621MxRNTCTysJbq66S6+AOltnKxa/d0969Rrdqmu5zNQGBTFKHMaPoIqd1q6
BSJj0wpB6jkSH8ah/JkqHuYRTZHVHxSS6CZ8iRMXFsbNv9/u2xjuBmhZ1XXe3Vtu4vP/Oevyy176
7IEjVni3ZVefT9oqinS9PoPA078NOZSyHXgq+ZkGsJFnIlh4ighFg69ru0epC/mE/iD3CsfKRJTe
ft72wohTt42bgKZnFVYpbMxMuvdF6bECbYDd6z7h3mAyDCs0QPer7IwUBsoM3PH49x4w+z5uIzE0
4x35whjABBRwE3e/V+ZizYgoYHbzPCCFUA/EoEfCeA/79R7dtOAtFwQrs12tsVUT4XAKFvXxB8W7
eCvHFJJJxqhtx+TYn/whlI5esRK3HDj0jWa5NvPdPI9B5xq5KQQTFGCFDb1Kyal7cbS8PF4FHFeV
vRZkjbdmBPr1Ecpb/L/dY8tlZOUCEjH9bvD2jmpBxEyCQlCsvF5wt3tOCFk9L+uWqVE3XFGx3Gd3
KBvJfKj+DW6go9ibDfuDEGMP6ZxV1VLqFrWJ5UavqyRdy8MWvLkBMsCnXH3xOfYVufVoC1f3aWG3
nnHlWew/KyTWbK3pDDfekqeT6ovNBo8/Gdtx+8wqsmtxZVYDxbQtOF2w+uXZ9+h1vx4NtEwUdqC3
BwBC9fajHIv43GXQndHt2arIe4JojKbldDMyT4VtaFtf0Le/pI++fbsVxt3/Slesjm2itGasLYNQ
OhXpZcb+WjtzIMeAUfzapDAbQZtkXggJJOpyelJaQ5ljO0HIKJn/4A8s1SpERGbYdN52bwbRxWUE
7zfGteflmf+oW/TG0/PFtjQqE3/nKB4CA+NgResQ1nEskfFXYV9g6VI0PM+nxMLIsqeTU5elpgHS
KQu2vMYN6dsNbXwsIyxUjmh7DpNNPnGbEFzPx0Qov7CmjDNBwoTyPgs/KWDgS1FhxWQFK/bKVmr4
2qWnqq0Wlwt0cOW0QmQyblRl5W7g7bXbfbOsCCsw3r8fW2L9lPjDVLFpduR3gMtpCjjCqu84l7xJ
m+Bm5T3s+vw2CEk5squ2IWgAXuzdLXtKowOhltUWAPnN8izkHId1UZHpYliAsWJVMFYE7uHoyAyZ
0RS/flrE/9w7xO/uqFJ1oHDxKJHSRRsbnotTRRPOLYFLXthn4PWcuBHnnar+kklUscX6+PM42abt
NjgjpdEYKgwSaw0nLHIz5pHf9oOAUTE2frYfLLOFQTCw5x32PrYRoGRDSuZw7uKJ+wgohxGRrQ2b
vrmaqhRyCxZ1ZmUu1d9rfbgJnpk/TjMMyglVfLaLoHOpiwggmrIprckZoRsFNbHgLJZ+B69eDHVF
wEZtIenFLXBOTEZYFNKmMvi4gDHNyOD/QyEOTm6PyF1j23l4P3xAxN4/iSVMboG5X2utYVhGC+jX
VwWcAHVFWzZH38A0wqfM+Ipzrw888S00XNn7/pBg3eSXVNORnC8t0CSifpREzmbAsF8OJLC9bCEG
PAFDR3KDkh3zquZg1UsXoZ/Dt1Erul/zPMJPnQRqnXnZDRszv44sYKwSFcxOm7XbGhvMkemmK1Xc
fdGfC9dk6YA8yvbxw1q47ZHVed8mRntCAxfcrnQMb/Zy7bDhun7u9/rLrZvh3AJNrnjEMsX8sYeV
Dm7W1A5GhQMWuJ68k8EUJEIKhuSmRAuKT7lrQXrw2v15LsHH4i1N7uTY4ebKDwzrwPv61PxsNWLd
wTmal3rVAmjCMbCmo+1keDqEVNPWny9YIqehYp82QfXHIAsFCuA1H4FRpQkhJygbm2ltJhEmeujV
X9R0GrKkA5wN38f61q2+DSC9aNRdF65piM7ktmvv2tHFNU/5gLOQrE2Eejr+MBN9I+x7+VV8mp22
c2cqdl9a5j8zCw85jI+YrLFmtCWPbPh1fJC3sFXLGm2Qos5mdhu7W1Z7r0hrv/xKT0/6nEQlgw7w
ia2RjesgJBTYnRAhi1S24rk1ZjegHlrvMh1VMPqO/YHMKvxAOOkNGUEWy65qBAsxHFhQszDW9Zo0
35jlCaHI0YJ3hkiUpwHyXhY2FNQMSY+KGKMoJAlWwJtkjGjOs5c6J2ySIC6mHqMVkfIWb/vRXEgR
6D8kz9ApO+U/eoEFeiqL+uvlfNEmm/BoPFwseUvHBTogQCQOufCAuEyz2QeHX3Vul9L8tzix2JtT
BLJmptkOtuTJ0EjM8yNhMvuLGMjUJhRf7uTB0yuIsCskafeaWkBJdq21SAa47QbrZ6Azy7pzEeQb
EnEM5eMEQo0NYeawaWC7I2elmZ8z2P4xK4dAb+1VvMbn+MFKDSFCbNX6wgj5muEqOJ/H4IB6YE0K
Fkq/AJsZvmmK+PrcQNG/gv0teaQE2iNzjJ/8tEWF5PaN6JlxVuD5BuaWVDKmdjDbjRgD6N10Y74l
oHk36MKCjtH39Qx1lZfl228a8oQwbvEd4b0pnGv9Kf2aD8olHIAHZR0MfSC7Di9wIuohVWzLo1lP
c4ndxCmlhw7geKejyyY/Tmxo3HrQmPwCDggpCjEwPSFb3GrOz91ySuos0YSxpjg/60yqCG5Xg8Uo
eCk3XO599H37ZLFTj1qT8B9H6uKMAkG2eayIFzZVpDXuQ9qs7v7CNofDZfQoCVodCmc4sTLbEpFi
u+awztM/xniposMe+xPyflSLjzESqWNx2/YvBNCJyA4K4hQAJ9HoQA4gx6S4RGLFZsmg/q17UKeJ
++C5KHo/ugscFLrZcSJ/sP6oXVYtjTlU7fxnF5N2QLwGB3jMm9D2NRHBBljz1Ai334hrh+mF5t/X
JIJ2V2beSQtfSBBANLKEz8Egpn0zWLbiD3gTruWlv87CCmxw8m9CHG8y0wPK+EfkMSqvqH3VRxO4
Rco8yv1oC+9QzMwSA8zXych3IQ2Er12oW3aKwwiNhT8tm+v8UFUIUYwKSJ7D9oA+IwT7vO6F6qmq
QXk2fws00e/d+eGCQYv2Nb8kD72UCbLWil2Bk3bhF2NnYhLMbtvupt8CpHA/mmosFtiDiLBK5Vno
I7SgfgxKUk09y8+REDUyi7FToim/WjG9QyMxi/lz8zXgskK/obYqd56NMb/Ax345/evk3QZZL7GK
gh8I236DGcc9LRpWOQPyh2nrLn6wPxUNMt/EeOh6XrOWY7cRiGIYjbZw6SogjP3KHMc57MsoTRVR
Hdzan6sQjEatvIldBK7UVb3nboxasv57cV3g0yOlEboYx6n34/GIi5EX132NLOEdyMvYHqO/VfNx
NAyK4whgE2KBqSM7tjKkj8IDbf/9IF2vMAVepldJFMnvOotgX6Ao8pVUTfsZ5M+98xJJmnK0/VIi
+RWD26vo9wJKd2hWTEQ7FCFq/fQ9rEdHPr7VC69oOWQSNDDS2OY8IGktaaP8drMZhaNMigfxZmvu
4TD9u3u9IDpxAXVd3XF/heLgyOtANajnj0+TMNbsw2Cg5re5ngUZKF8LWNK64hGZ3cIGr7QWN00c
s+rhun6ammAqaLWyzHI=
`pragma protect end_protected
