// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1PiUiEPI7AdxrXWqGfX0nS2KQUw6OlvxADK773WxQZTqJ6OCmJK/bYrN/EdZBqkBmzJjCRI4OmDl
DJCHYOngHW9yS+GI55o4MofbJbZlIuMC42IfieTibz2414JxJq/C3XP/75rz+M4xyzJxCxP0Gg30
9QRr67BKv8HzJAAJiQKif0Z6uhC8YhwquqSkU1FZEuBlf1aswp2FYzNc5mxD67p+LvlkmMIPSoiA
OEKmFB0RdiL/djfGl0bXkCTYzC+HYV8kvnRMzz8nxILI63AzfxHj/Lef6WhMO3FketdEXJIxVeO2
wZvigVFibM637DvHJF/fOEqJnB4olPSTCqJFQw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 34640)
UuDOmtuX6Eqkgm6pr68vKYUQOXrO2fU2JF0vbABF++10IMLUZJ0oLdYI/++iMDvZF0jEZRRjn55W
yAYKh2GyvviOoH49RIjDWU4p9/T+ChEbVjXOV8DAA7Y2KpNjKVcrfaUzJuPuSIiUx3xbe6q2hoAW
ekwKpJBHhW65g10PQWrMerWa/lqWmo7iOZJLsAezsvmcnAVH8FPJrlVnc3FGIu9Xm9ITQEwo+GhT
3pkWuHX17D3E58nd+r2ZXDIr4xQOR3U0g85Ryz97/VGXWug22S61tuOn0lVO8E+RDRRXcldVIeB7
c/lkLSBDSCramBRPadgZM0JLAF8dpQyww7FTmGSy23r1fjqOl0XOGWk3nE44H1JCxgQ5UXjS+B44
YuRAigCaK0ljzxdn9ouUdgvWDdYOpLFEFd1N+Qjv0LWW/xLI+rIoK3vmsqv1eJU4Tfdg1/uVybuV
FOqIDTIHaEedMTbjcYwZUsNbo+9DYD8zx1vSD539ENCqckvNpUfH5SltLLCFr0+oeJdaRsY67zLc
eNNkFZr5isbuGmiRcSeHJS1ulDkCww+5X2+iGM+7I0D/dNzaQlXOPH+uDnIGdaquxaEQwY+G9Umh
MtVoUwLkLc4rvH0KltUbc4BhBMqrOPF+A/INqtOzyJI3xfTUCo2zWs1NQZrH7u9jwJtd46UEaShg
5q/CZkSB27TR9+3hQD61S7eaGjb78SvMIY0vnWY12MyHGhM8gyQzqLLrFH6PbBjiaBDT2IMhcMfv
bm985B0NBLm0HKCYAyekjCvNNfmNl7yEdz/WYnsGHEqNizZXOBlnT8sBQ0zF8y1c02pNrUUoGa+D
mDFZIZGZSQo+sxrNu6M4yJP7kOvppNF/uGHti7kYksCe3RYUQsW8ZupDJUap7xQibGK61lHbqkEk
uxK3Gx08NZrpJrXjTnVMThSsHqgTQ4zupWvXsFywwau8NuD542a5t/3bjVe9Y8+upzSfUZ54CuXt
X8oRrGZu7sWxLlabHw2OcSrp7OtDgN4IFtGTRyKPKIf8bZieDbgOReGP8Bf4a61yCyYgS/tYDDe1
FKvmEVCDVvYeAiDTT8ekXmKYIqlFVdyTijmKQXjWTN65KYWv1Ui+ROAMhqF7E/vA0tZ7CBwfhISZ
U1nm2Lo8QRvePXYD8yLSNKhxxHD0f9Bx2KL11DylmOUTfdzdarOvKI2d4QGzE9GSZWjyDg8BiL3B
OZbHNSqhGGnbb0oVSBt8Lus1vt1yuxW/EvSJkxWDr8OG4axgvops6MCCGyRU/yNtuBxrcyjvts2Y
ZICfa5mYggNvjhan4lt/93mfp3xj8f41FUbI11kcWD5crf27UWAwZtdDJXDsjbncKrZMnwoghNFD
YCISrtGXO6c6RtayfIiRMiyvcLFbR2smOXDV4kpAFDzoc+AGG9VZ/0tCo8oL4xCUwQBEZoMXXjk5
cvEn5Jn4Y46DWoZOCx2abNAJcVm/YHxebmV19IGW8Mg4NlzI9xWMmxYW2fFEsgXyWEMh/A0nuA1p
PeAxDmzoNXfq4oZqqP8anUjaLUs3rxDN7xxmVD7eXiFQC4FHtlDBfAfEEQc6smVXUm3H+9U05CTc
3r8unxtKfzWh4pYh30sjiFhjKFKs10yNe/BXMHSjjtJiVqSVzr5Z5E0DPElQrtUx5aMmtiGaHqnE
KJxNehY+wwEKexx10gfBnfo3MTRMn9MN0xEpX5iV6YvJLvLCIXlUqjn4P2mlmv/YTsSm6F4X6Y3/
tkYWqvirMuLLPasMQmLaWjjxZtuVrpt+dReFpI3OkJNbRgXBe7b6ceWhgtW6kb+bFS18OZLOcnAS
0g5KXXXf3Fbj2JYmf+rG1C55Aq/JB53CuDLPRXGYAIU7SiEY33TF3ZoHYHPY495XCToRN7xQtRFv
vddEdV2h3PvPEQ5ThDGa2YC2gbRYpa1tCqvySS+2Q1ZkRGlYFhWhOkwnccrgidzMNhlRQpLuJ16+
zYQkfh7PAflLnXbxmYXrOSGNAbiAZ4Uin+W9Q+qvAx5nq0dt0OEiAQ3FTCISx52Z5484va4VcaVa
8mexirjEa81QyTsK/72btol9IodzI+VW/58/qQN4hSU0B1B8KTkvKR/6d0gAzHDREKp7sSiTdMQF
Fiy2eExGH5/9NY4HFoFS7jcVsNM4zw0tpaSZ9khP5QIu311j0SUa94SW7p5Hzf4uznyqga4BsNUB
FcwD0qQU+K2z2L6++czoIfIudZdZYYgIvv3P7Rf5RGYeoFiZb3TuhNq9Lq7RcQlf4I+lz1WvbnZJ
Engcd3ZLD855AAEsovs/jzYeoXzcDNvqUdvz9u2NgaGTMp+LWGOdpGj7Sg1obrFRjq4Cr/RGNUS6
F16syfZq1zXd94ZbpMB1JdsmnroShjKUQ2E8tibUQyWICRXKulr9kupRBBl3DrReZC9mo8aUr2o5
+wjtQqAibyy9I4ZPHnu4oLLhVi08Lh+vYPd/AOT5muWZBfq8GvF+WGui8bcl56mYvSUuEI6eoZvG
Or/6NlcCadVez2GLDjSi5NivuSFXjAIjZ+zub7kiAhujxhen8hvPICeGLxFDbWMUWI6JUw8Dha6x
XDaBcPcbzW32Bg1dx//HsJuXdSGm5KSq4u4f/J63ro6Bn2knaoDjH/qTCQKF3afVZTxSNU3W3aDH
Ou4+Xw93V4KPuD4owgy5d13yVfqMTpomZnx84C1UiQ88DDmaq/qzjkC27P5YjA/jdPSqhZJOUYyl
3jDUM0eJ96p64osBIr4W9QI5tv0m4LIz4LRYXAUUtyjUOYh7wugq0qMjMsGMq091D39e1JVOtOmW
ifJ+8ykipG5+dgiRk+Cl8whEkTWr88W+kVMUJuO5BvyFKl/jmQLjoTpMlSnZ+XaTTdmyC13KORlz
49W7gwQRTrbeIxWD5UI6pDgVinKtyKVH9YdxOpsQMzSRKit/dfntJzc/ssn7FIpS5ejRUwt0UDvj
YIW8IhXkeDjh0pvGlAraLAWJ1aScIsf06NUlJ8pejbvgSiXV6bW4OiRNmWlD0wXctgQ5DDYAoRe1
aU5KtkwsrX1hGXPhdeSCNzqrOuqa+I6bEBclZznpWJ+rD8LNvnY9u3b6CQbTYUfLWBTSKNr/uVA1
jSYIzWYx3CPFxbsRisGj0EyybthjAG1OzITgGLtCU3esUlGpTOIEUOz28teNp/6jaFvC2LOfB86Z
SYJyjHv+QbuFI7RVh7BCXuteiAOOy3X29DP+QCKBNODVbE0OCAd72h6AR/Y+zEAAyAuEUkt6apNu
Gexxzsidaq3VvMv31iW7aiAMNk3WFs9J6EBHmHyDEQOyFIuvQCc65P//P+1J4QhspZ9MBcxtK0EC
drPpbO7/7Vw9rJdbNszA8P6RX0wk3L6tnej7onZtc/VdcQVO3Z36FJKTuoIHGy5l8eI8eiBKTZRz
Jk5VQ05mwNESRqyZqCSPa5wMvi4CICNTc/oscRxLaSa9zpnCG20NOYJ6GO/s250Ol8VCqcXGZQ6x
AkpWbsJx2GW3tZ0hDSw6NQq4Yl/n9x7wmj+zdIFonrJXETxhEgYubMVYD+lcRqeIq4w5LfKsPiwU
dlO4X+fB+3gDajZApNFwoihoNf/HY1nqtVw+/HDcwhlTVE0bhD8vyUAjlmTCmadSI6zuL0cfxikJ
Hu9w1uTi0RBJ9DGahmcFZPsLtulPECTK5OXnFkBk1lF3bQPWzR4jZQ5X2KEFIXtWSQc3qw+1ZGb4
TvTNhM/PcQQQ5YhVL9nPZzHwCBquX3NmmnOgk0Qe6JuqRj6eVArmnHORg1iEY86nx4af7/5ZEz83
o1ripZBvFZp3AUkFJqyklVaoycxBkHK/Np0rLXBzNxgrAZa0ynfZXpO+VBjKu3XYZ/vJm1twa4Eu
qaP+vc+uGA4xqDruik2GsWfBipCdKphqPeF+PLT5AMAluYeQe+5WFolO2Rl56P8289/qDoxMeLe8
jovIDTRZ0xldnWE/N67iTc/7UxamuKCaD52YMYEs6vAjSrocSFnB/ISOJbeAtlHbAFWVQ1i6fL/Z
q4LIbPsVfrxwuKGqZwdBAZDCPfOemd+N+cgbqOesmz+6d8Xq1mTOt/blL0vaH4G9l/KOq5gaasEy
/ZyiebmegVvJ6l8w6/LZuJ5UQdiTC8QiEbTBeNgw95jjpWY53e/hM5cim5FJVvymlVPR1MPRP3hW
YpVnWvzcu2eyE7Lv0yrskKjvLoZ0uGaEet1+7QtqAkdPZZksQzrTEJMiIH10a1ZK3X2MRdthgoKy
VIw1wel65rLggdMPJXChlXq09Fd+mXButd/pSZdQ1EcxCD/QUZaa83r3l5XNHiijZeL8H+krwiEn
Ay4KwJ84yNl8GCXd+/hK+IBQ6EasckyaSCoGveZGgLZWlDUym9+Bpt70JAI1B4eeDyZU8eurE/92
3Im8gToFzRXuFfodmntGeS+1dKz2fSzq7qhrjMYb5XSjbLTAKJTcr4EA51ZXGLBTdevMby2zEzS/
kRIrZXCgJkjR3K9ZwPS6PGwEV5E0PlrspvyFA8WODfs5m3llVA/DA6iDjtLarChWGpGKe9dik4w0
Pl//WgeH+mV0x5Gnugb9Nm3z2xroefDZ14UBSGHFpnSzL5IAG56Rjvh5k2UHKqpl89qj+tewhPO/
tpsndFMB5LVUW2GAWJ2rQLVC+opxM6ehh2r8c4mfk5oznqVHXWyQco3XHRN+47syX2iZ5KiwY1Se
Ga+q3JrDI+BdeVF2NRL/j/Z1Z2I/m86Razii5gkst8vloJnKjS8Q+zonQ6YN3icROrTMXd9UfzgV
Mh+B+aAJpsQUOgGJC6afvlx43PJe9SjO+AuYVLQPnd3BQCxOavsfQe9mW/zhPCRgXivLaVUYlrPl
1bRXAoCGIUfz9+oXvW17be9U/i3jZkmqBM2dQa3dNz/VvAlhn5WShca5ilX8ySJuU0GV9iaaDl98
v4An36qKYjA1p1hMHiLjJqrLUqloZBi7R2mtlM8GvDyeX+vs9nwboDeeZAUYld0craoFZISBfmWe
bU/yuPDf3axmrSdjHvwGUtRSlOSrNQhcMWrEfyV4jmcQR1udkiqkmRFqtWcoSkFBCUYqwbGafEq/
GB1hzydHy7csnEGfFv4Ahv/sVLVDa1FV7mCQjAdrc2bofPAH/L8b+XgQldagzOYmAr6omZxu5WBL
2M5bVKo+paP9mp5Wy53cyLukXkh+ygF8yQ3hJujUpdsybFoCdQSbENUtVOsCm1F84I/3hUbtHX4w
1TT91Zq3xAm5/bwi9oLz9uffDdgh+kLiwL9Lgrg+mZHVbuTt1TQ/y3c8SDSEvVWqqTYlIb6rgOd0
BzT73a7yS/dR3YsStOaoT+mQqIns5DyGBRasQpSOUL3gTVzsLiZSzjRtxC3BM8MzTtpnSH+VyahC
tIi6zLQNPp/wf1g1be/7HJfgUz4aRX9DPJKiQc79w1In/lE1kPVhUjoik5vP2t2heymes68U+AOK
S5gZT5Ua204bxAPzVK79X5RGO+CdDUyZvjPmQOMNXTTp2n3w9OAfCkR/Zkj0jCz49leTQFT1C4u3
S4AM2/yMaRobFzHOJO1bjuXSqDb9U7VhgLJubtDGN2vD+UlyyQWqGofm+NL5BN3ZDcVBCkFDvHX7
2/MVRC2Ks48fP3JWn6NkNu6fyHe467K2CxJCIs3XfvzG1AtjWGDxms/EfPGL6LP4mMc0sInOeMip
FChg15dgzbU85uFZEaffgPppwJE7+04W0m70XO7/spDyn8oMU/kfFTCLnKVjmeqvr0qwvAMKZtI0
xOqLYGgqxvaE0m+i8S6eC9T4OyZ/6IITRg2cMHE7qYVpw/2lmiiT+9B4wd2HqScFx4PWstLbB9Bb
y2xD8N+TjpsWHKmaMQ2/TOoqrn40+wy7G9w4ogNL55kVj9535e2WblNiTXIFcyAMKh02jEo67sFb
947zLWKu23cBrsRPnnCoQzejleaOCic5Nco8Jxu4kX0qcVxRSF77wJK4k8zZPZMfNirHcUyYJT1W
shDPzw63knrVBu1aKRaXd3RUsngVJWN7TJkbzgYMqBkm1LiTmw08JeyrOZaJlBtLx/pHOalU+26R
tqH1YAyhI+9G/bHIIgcv6lzGaYSNR7b7UR09LvCaN5nqQEJqIOjPASybIuNuC6oQ9H/hUoX5miSE
qL0o48+8Yij0Y0aO9284ovAqImdOibh7YPTar0uj2jIaMTCkK3nd0n/qOUM8GeWLXB9wCLbhjjkr
qfUaHoQUGpPaaVDVFD5vsf9ph/luC/7KLmRz9wPEIjU9KcjJcq26Vj1fQaP25LOUDFAgsLsmADA9
qLLLgKm/JvhJji8zbBGky5OUg+8EgBGbjn+vF3+jejFmn7UDceFx5WkdDsZ9VbV9hm4mSHvoC7Nr
P3XgoxXcVvc85Es1A4i7SSICLo5uz1ukyjfjbE32PuwBEABzcJ3W/sHq+pnuyqUOgyGCWmwmGsdV
8sZYxv01tZuhmvtrLjAg/xBDGQrSr3yFMnE8s2GczMW2ucMjl7wno8821KaxCvMh91SrNwvKGcuc
C+YYhrxrqa4gPjhNZV1saaYRddmWfxr15lQux41KXGzGgqlQysyNHNSDwNhuU9gKk4GjxF9+LJxY
i8oh9mVIQPetRdXSCvXmoYF9l9iM4RAz3HOsD15V0CalCA0HottZzUk9QvUSrcBMtM06YB6pX93J
BZ/hcnlShiNv8J3uQ8immpF2Sqm54Kg1xrftYeJ0SRraTCxDHokQRvZ2q0GJf1KW0Vlib0zaF3To
V2SW5WadI3WPpPfc1hYncXCFj/vr2Rw6AbdxydeGqE50a3G8QI2i4uYz203H6+H7gR/q8ZvFdsMr
zLWMq8K8KapoRtgyQpbOxQ65E2qTMvGQzab8SskgN8WhypnWg9a9l9dGZT94VlhWlfoYuH76g42v
OSF4AoLZp89zRh54PT3FuNj2hbjaXLSylKdwaBz+wKWbetBtd8U23Pmgao1ZyVCe904keOPxdrN2
EmNrrxb7n2fj1kOkewjYVQP+cDICEtyhMfYvuH3yH0pkwFgMgjRqZvv+ZPs5frqRWXe8hn7PbyK1
2fs1Eo6iTtbV8esYcthpPmUluQtUg7HZpCSxz95qXwv4dk386TFph63DdmNbqMjvxBFSyhzmjLx7
qtPQyMDfRyVm9VqLuESnjWLhiZdowvTimAyg58eIA8vdIApojmk4nky4SNdcXs8N8FSacDtRWbhm
7aRODgbG2O5oVolpDef5OFYUkxAhfPtX7tmpOrex6Q2BvZz+C4FcCEMWvRddcK780qS5EPGZSgxR
16onoDb24Ljef163ADAjsUtT0mEPxTmS5PNWstmwzdBJg/92DwUQQY5enPGYc1Vj2AbRJK7HI44W
d0/sozDoPQ10Y7JyHYUhbdpo24nuaCchZo0SNOAhGKFcQIFoDHzA4XggvESCDe5S+k2Zags07CFZ
u3zGzhVlH6dGld/MXEbxRcI7wm6i+soU11rZ6gHq5WjgVPiLpofl5r3fZXqtg5ysoQVhhfRKpdWP
vyn5P7w3K35npZDYk2CBps6ekSAyazpHe+gAndMSE0wz3W3o1JoWkxqG2ZgJu0oR0eiJqANaAEpC
RXssoVtkVqy6o/qHf71XDzDpbrxuWUz/BSaEg3ej4DxxNZQTXjT0/bWWestIrnoYXsbQ33aEebrM
6x9tmXTv/Jn+pah9JNmqVwF/2GLpWCfP1CWctmbIs8JQ29gDQLpliemR1QduYFMdalDK9nTNYSrN
/qsLET+o5Qj0zUITnOMvzxoJz9PFbzS3a1S1V5RjWnBYfwCmpdwWctCzoyQ2trQcvF60JQRG7j2l
5b9jtMg8CKwL3+jLdTXd2NbbCYgwRQ+Z7EF34A9FBQWPgXXKU56JVXHOjMGq0mjnnfc/JoLmnLhA
Y5usU3EuIti9ULeRviN03yAaFQ4hFM6MZ+L2p94YceL0ExGK53+eRCtj9owMBM4FM1Uoqdal+9hS
B9T0DfdIZr8Rs9gvUAm3LCe17uygvdensYbc5hCbjHbrm3aatFWxlIDmY/vHG5rzGOoQYrKnj/wK
y7AKkIzb3w9Bcf0LSL+ukVrKgBTZ3UgUC2OuU8LGu22sEtrbtCJ3JCWMcOk3YieyBllRmHk/N3i2
zRCoh65GbWphFHAdeC20dWeLI+HExIwwl+9vrdtbi+XrUoBRTdXaTAlIbvoOF4BAPb9OjUiuNTGP
S0pZlSBkodhYYd5ZS/4euZ+03/uJsfGcsRhJcJrvyNJPeKQxCQSptXleZxKrMIdkX6XvU0k/Yrc+
oCDkSt7FiNi24v1c462Hv0kbZFQC0ISb0taZ79tNfisFp8/+LaSjKz6NvaPW8ce8eltMH6DaBHXp
b4MfebrDtAKX8j00q7c1Tg7/zAK2ToBxSnEqGttSWFnT2eNZft9n3ENftpK/0qhQhGWgd70zu2xM
2RPmaj3r+6JqW1JK0U38ddTZ+PwmxZdwgFPOQuPz9pisW5YSMzMfZj1ZDMgFYL/tvhQVd6ADqweE
WtFb6f1Nsy0JDfZGtwKrc5VXqf/jaF5HC8Ftj+XokTT8Lxmym5M0K854ik/mit6KSsIN3DRDdYEv
tkdfJb351rjoJAHpkHR97sJRxqkNrSrlK4x+dQj1woFk5YkxHDyoieBGWEF+kdaLsJOV509LzXPY
qcqRCimHHHKi0nv++cgOQ3L2C4/E9vldk6qe+INhTj+zTOgF4dJX5u3RH3eFoUYcAq0zItJwAPO4
GGFJCFBRO9s7Ln8QZaLXTxs72cEWsbmZDXgYjoLwi64iYitSm+zvFcHGGfvCd5OsWcSA9w2bSSFN
PhEcbaSHOgwXb8sr8TgwcZhGIa1QkRJA2fXVdggCq4f8E/esYvYRVpat8P9RAPnmy0lHK/wwM/pd
XBj9s0m3vcnm0e5sN70tnMViAqyW/QdrO/JV32XkmtoJgG0VpAodBZD0rDEQOXrPtnGZkAl9GW5+
oKp2k4Ew7s7np6f1Y4carLps8UBZYLqGEZk9eFFkwRQNdfo1+kM3JgZWQ9DvBwhbi1WJLdmBocCG
JYClfnrQYcl98R8aj96PfDeBdRy1xbkoLqmGXMQPtNyV/EEUbc3cw8zq1anhDp2pyhHrXL3ZxjBn
Nji4w94i/leITDXezQWmIuVaHxEkb+tghbJjkJLosFIaO5p3RBlxlPxb8uRgV1ueZvLLngIKoKSG
VERNmluraixqMDG+7Z79Kg1O38IFUnpzbofasMcOzZMUMPzP/Lce26pKY/dram+Uv2z96v00ElvF
LA+ovYA3U8/4VVVl+A97H7Yv2nNDTHM8wKs1nZF3iBv4bIQrCfVSrMqt7e5w7sd0zXYevxOW7wY/
BWZBoYtNpA5C4iLGiscfal+5cFEmFx+SHmRXLyssBjYVdrhtLSWar72MyIREtu910mxntDD07ZPw
tzv17rw/FVVkQ0R2Tw8vZIzKicikH00yZqZScID9/F4/KOsuNwIF69OVOVphWLIL9mS4RBNtndJA
wU5tNtoYG8K4qP1ukQhTR267/9kmVRnQOV0F44KbYeqVuDeN3KMdyzWbJAq4I1xxlSfcH1ZcnbmS
CkzNEvUH2qYxfDJkXc+5oMr9WKnKw8RdSTT5JvC/nv5N63bodxH+m/IxHnKIceCM2psmQFM/o1lK
D1nzhe2oZ1RRc/TMF5x+GTdSN8dP04ATRpoJmBSRSGAF5chznI9FoyPwc2s6vJSp37hbd1wxotrI
trFWwa7eMfUB6Vzjh05KJTKtdh+3cYDKW742Qmec15X+kjU/1TLLiw1/YNsERjrDVS1b6IsKJp8e
DgJdLj+Uh10q4mGbkKi5FaNC6A6LgmV1mceAWkmI0ETKRTtS0U1PZdOOm3E/R8XoXEjY+bqAfdFH
N8uRLqG9eul4+Fsy5S3X4lJubf3jDnVgPKZojBrUFDUwFjuZBtmMnSlENqp9ZKejhOUFx6Y/aQnH
b1rf6KjeEW9PP513wan4RPrjPJvCfTJE+PhQlQ7EXNngFkM4+YbJ4XgitqqpZpjOaAVdLzKSf05+
nh+/lFlpD/h3NrTt5PXscdR+CanJDn93rFZLfgwBunYyJ8x348Onhrjzwzc0Ch0ijjimVKsVC3eu
tLwKBglj7lJrMiQWZksb4RwDaNXdWwpZTmdua3nEPoF42ZymWOCNP3sFaAxyWiaLJoSdfnPGFDZG
OYZQRueNkzID7P194UpkX4rRz4WUJJnqKSk9533vclOjzrqixoA8uzqIDeG1uvn91N6to+PdmpR0
GAxqZkaiozycDUHdyb0PdfKQ8O1Ot9m1k1V+P63YtCNnNDaT0TbyeZ3vjBbh8xpLb61RvwOqjCW2
niFQ7u11vf3mertEhFALYBFFjIt2U8HdTxwdvw4AZuD6rvdsjs8Be9BvflFIIdxuj0Rhlg63VSQ+
t6cZbIHrlGiTX61viKq/6T/RCgfoZCnJ5GTCsAuFck9/xOUbyCySmyo/xcdqZ8F2yyNyYxit/dAd
gZEplSAA7wOCdkcG/vEwf6iMc3VD5uXU30hveqfkez2TxvktTKOvzpnGQL2omK0eqy0lhxjqZ5eJ
e5HSsduQd4p1Y9VNprK5xYSxp0rBpfAC+bzyMWNe0GCoc5EFT1U7CYzZTH1hZbW70tpUcxv0rqcs
hgPnhHTDnC6se5CZWH28WUxL/q5oYh2/xuEEax5VZ16N2k2uac+3XrynKL3V4kgN4kLXj+yRXB1H
13jgmO3SxyoyvkW95H2B6qtGe8J7cqQ85yLk0EHTy2ngF28Gt4B/iwAmpDoGrF4ojAnAsYr7YmV1
I/l8BTiqXcgfnNrKkWLsRmVmBSTQmF73/T9Up7nRLzYi42Gf5yCBJFAFiTE4lKABdBpbaHGlqmRw
3OgFa77iYr9RqJN9ouwPHtssmqzTGwVSrBpI2AF+MeVIrM5pUOBRajqe7i+bh+7vCUPLBXes5eyH
6a9hqW/OApVTnSZrR8CYyZm8YxNhKH7OUanWvL6E1HNMOi7LXszftdd+lRgZf/x8R4rJlQl+4r8I
YaEy+YU1HVxZX6BVrRKctTRB8qtcXUGz/qQ7VHtUCJbhO8X5KqVW8bxiNFFWQeq8hyqCFlJQPLEa
dhcfpJs/gIolkW7Q6DDTcMb0itax+tyaiKzkvR32tkQ21DkzWlIv1MhkjcS160LD7P/21xNzhooa
c5VWFtrVkH6KcVc9zjnEueN3CDHQcqMYrOkLznJb/cG9rlNuRcrApMSM1fCYMxR0jThMIy7ld3EH
73w1zKHj01Xz9S4nIXaZ1zlVuDXqAxMXeQHxSPr2uPry9LS64Ekl6Np/fTm8LF0o821W+SnRU8ph
FQ5L+xmElDyo0CxOoQQ8MebPt1auoO/k1Z5c9QY7uJgT6lqFhF3c9KpTElCe0yoONMXjG/l3nib4
cfy+/YGuzCUWBW0sgqxqEe6WDH2QrQvz1F0EXPZgZ52q+pzbhSZ9diy6BD5m0o45OTxko6H6O5zZ
xgN3A/vYFgQsl1bxrbA/p8IYmP4I2MPuqkZfSio7N2ROJzFXrx7w/gzeGXejKzDR2OFltwJYZJ5K
6F4V+QSbHaQFWEjHfyw9uLmdMY/zjl6kz4+yfI2CBzV8Fmic5ps8BRBFcQLC4UfuD0I3ozqaKOuV
cnzMNkzRfMBr45d06Y2bqkNxBFbNY21rPtTu/Hi94prqWtX8pZREKO1x2Uyyz6IXA7IxXhj/ieRC
aaIS6JhI7otQ04xOP0dsaytDMpqvsKhO4UOW16dYjVt0m1YNDuIgysHVom3+suoito9DfBY6UgSF
ov1u8MLRKkZXCIzFIT45bmBGWVcMuaLY6sHSjpxm/meyTxA5nsjTwt4782E6cIdRXPT7XFgvBhDY
yMFQ6ODPHqVCyPOJKJzbqST6ny60MYvszwvIPtYJVyrFDHZ5RSFGD2+d9SWX801WC7WYdcRE5v5w
bgVGsKDurLEZ2mk3aWpNT4m2tPgUA2mf+OM2d38ceRxTgfXOsTGOPFSiJqFOHQoFMOw98pE5VwYU
wdHlvsBOMrjOAAjtB8D8+tKaE2/24KJKeoeT9IzmSU4yLOY3PxHC5E4u6JpUIeIMEfuf+dt03MBc
xFJ1WZH08NS6bPexm5wFyzCMs9LrElgHRkWbVeow9WVB7NIIs/ykGP0kYu2RLy1CFZ7ZpdIgCXbK
kvUrOH0s17BoyUrX1s6eNnGu/8YPSB9/DcSrHH7+4ufbx5BsZ7Hv+mlSd5197vbMVoVD7Gyqsgq6
4md9H/QsI/Tg5iJD30K73UL9uAayvv8gYJQ+sgZXpdYb5lAw/3UP+pXyJcvha2uA9mgMMOrqfNtT
UIxtY0hhJd/olGNtsa57lxIaY4W2ok1aF/gYAyRwhD9vTlNhjZ+D82J1QGcbIHikicyRC0Syy03a
LA9hSr9aWUSBoyc3ungdYlDDtlqYdNiEfqjWN81Grm6TZFIkf61fz2GQeoxTwR4KBTKxFoAlcAHQ
04ayDgbBTorOEaL0DRElqGz1MK63myN1i62kNzcat7cy9lYQofb+ktsQPD0c9VTLmzQ4xqLt1S+v
NVYgdmyaGW+MZdGgTEy4m8lvUZG3azuyY1Y04CilBXj5wavQlR5ovu7LvT8XHr/Ysczku7X9LK17
AeTUMQYz6eyK8/xPAtdUkX8yhcJvAQtGrKDNkPo1mJpn9+RzTiPfr0DBKaXhb+7qIkA14NmdwPm9
/78dvfmUmynA36RUVbugkM/KSnBEhPUT/IBKt1G5wy29MTkcdNmgcaw2Z1zbmMz41X6f22Uo4LPV
pYJaExqaDUiXcvIs/OsOwLKDektXN6GYdcF9kwvdUfrFHAiRwfLAnjn2TFlo5m2S9e0Fo58hlTuS
2v5MihvUA5iwRBspBRP8Ks404UOVUeKNywsh0JP2E9DQRIEZ1jO6XSG5tfMWYl85ioQIRWJLr0QU
Ifo2GhUyr+gJ7q5Z+hxN+ygdTKu/oxMpBXoJk5TcPNqueWStbTNticL1eKSu/l/Yc9UfxZPMder4
wJvCGTwMo8OM9uULkcxXcImdopifFSbNaUuGeov3udn3l2hT042ESCv4Ay01URDGDSk1vwfxd+W1
b+DvJLstk6ZyOl8wRo0YnjPu7dx8sIHJVwTAE/MVT3woiH+3vzYz+JS3yOysznosD6qHfvmt+Rc3
Pfwd/VAkGo/3hsQQpWEMXyg1MKmJrmXNRduBLCm88ylFvnDkH3ZBGefQmu5qTavZSzjAZ3bBSvqn
iJbD9PKN4WuXiO9jY0dyaiUNa72DxM673/rh9onxEvRp8/T+V9aumDY5FZqI4U4LGWO8/l+jegr3
iJDdgvR2ofw+F+Hr9z5T56VLUDWoDes325ASiD4CEjL2x3ebUxoL4guL8uxoq7xgwO56hspgj3FD
BQJ4HHdTjELEeMM1yF4nnwWqTES97T3f8Kdzl1HkvmOTHtElekiKMZAE8/D/bk/zzQut5eO3JeAf
1+a0US2M8t9KY36gxk9dXGVSSrbB9qJ3+8Dpj4y358ASqs8BQvQOZ6qMUCRisij6blt+cTpuNNTB
DQFuGN+r22id7HFVVgNJQyOm3OTfhg5uayd8x4R07VatrbI5skI87/cBQsZKNGPVRrYYCBLL2v5U
LDRfFg+/0AzJ8wyeL8vHEoRz/pHwIM1/Fk+9XOOImG1CPRSqdc6gkuEVy1KWyY3KvJtf7daL6nbS
SMz3GzW7TNeOXwR5wDNLB4DTJdPoI1zRVmTAVzvN3jDYVXAvJTdyVTkzGuzOrXW6GuCzCKwFQzQa
O3nr5YJ6gQoK4HJxBU1tEpPHi3clVKSJBHGqtFzg2e/YJY7hJJM3d5/ef58hrDVGsqSlm5tzFlAu
q8L4hxJ7LpHMcqZQ4ZOzmw46KkSV/eXLLERtouKgiG+XZY7E2nbsj6aP23xJCF6XlXfrA/2eUdeI
qMz7ZEyyUSnGF86tLnFE3XcepSk0n7sMe2OyVDHrFOlsMSUOMhkhrORF2t2rIxfONR0v26l9NM89
I7IShFx4BZHQpgZdykn2lCGSVD+494S9gNihZ5it9jzJj4hBv3YdKNhl9/vKP91E0jDx0dHZHDii
YmafeYBeKG1heVlhlVUq/58OlRoEo4v9b2rd4PbcTcXGEi1UvllESnIonEUMVfX4XX8wYXx/Ywwe
wOS5+zijV1rxxmleh2UA8jayH1UC1UwHKLhFCesfMhQ9qcwVfPgql6q0/5bf/1gtO8zn7fRxQjUU
mksxB+L/bxxx/WD0yGMg+YkRDw9Do04PWUs/ulB2rqB4TvP/R+JWad+QdxqnXMvOmKQ+kVSZFEnR
bZECzptnvwZ56sPUiD2lR49WCQ4Ai9ZSBMNQiC0Zn4eiKFh8lMgXhFdl/smLTsmfjWTZXfoErdBv
Jst13kyK6Olq2brH/IWYhhn55Pg8mwzoTnaNZBI/vYYKtW3nm0pVcte0JbjoXjJ/AXxJaCrOKsz8
xNTBWvr7cS5TKZaHp+bBuU433ru6VzYovmLXhWW4KrOy8kIoremkYA6+A7tY7WcWpDAQN3+Kxa5D
tYQ2irTlEn2aH2QprS2JK6KI1ckhZbfobiagzGAlFQ9QX1HsQa7H01+3GnDyNEy3/H7usbshaQ9l
MPT6bADtOB5rxjTh8EUy5vXrbVXnIWCnLaglF4XsIFMKWghVIoH9lygWN/vlJ3cf2DHoZUdFukoT
edDIp7f0x6xkzUNteqVBSSS9jmQxidxXkL8L3xu9X1nBXVplwNvZ6XnRm0S1NNOi82CpmuUr4hHr
GDP+O23Rz2OUakX2sDB8clMlpXWRe5iZST8CSPi28Vq8roEmYTvVl0HOMtoDfwILiFmd2IKIGtpR
jkD1hHAZ/P/544VVUI8OAdohKGU8cs6odPw1qaVCMYkI0zqlBhoqxLCKOagQ0lFEPFT9f/zBx2o2
6MEc2rh9iIJvAjCtikzZJ1gWCNmESNVRmqIvyEN+Rye/K1VuPXmV+VxXNSXBrz7fy3fzN3tcet67
kQLPIkSfWR0EvesaVpr79Lt9TyidnqFHBABdT2cXHYiEX48Gj/i6wDS2L8ZxEHYB+1sz0cK1sKQ2
ttGK/7uY6x6ENzYYcMHynEGgVNvZxFOL06kLdY25/OWLg1MUCZ5drvz0bgM2lcnGQfeohAOguNRJ
RDFfRA8g09QdQfUFy9iz6QwtRtR2EUd3EQmUB5pYoCyiXAX518z+hL2d/2qAyoQvf1GG/Bo3XEnw
fHO0g35zkhp/wVma7WbHXqUGsXf+h9sivoH8BZPKKfsCKhfE0SXwZHW6XLmVHx2QgjIvLhyVMV4b
AcIbbNu7JzPXRoas1ZGMWOahGInTids8Qm2rsUcjJN41Y3Kabbsp9PDWR9zTJg+A3av9U6qJg789
N6y53KOwpQkx/zo2yES4ZFlLepikD6cvuDt0c0r34f9/CgBbtBtphn/lZyrOqYn+CJkmAePEiKeX
Efas+Aeh+X3GFBTlvZgBGshBIPUrDDvHGuRv5lLSxxX8Xz3rjfPzr4zZgYHP7kYqrMTBSxUXYIVB
W5+a3ueV5WP2N7hQTZ1t3b0SosR5jANxuyHSC0ubDSHxy40DqESL0jm/JCL3FNHax0H2xJfci/SL
/w1M+oj/f74VSAq2zE1byx1STjw243uV6km6cXU48QJmBU25UAh6na4sF1AgP9K+RsEWJKsl5yZ7
Mz6ikvPjMwzo7OD+nmZmlR+wfZj9I2IEYxTfi1PC1qvuhq/nogAxoCqxEPBmoAC3lz2+xtCFjajQ
deI/t7sirWIxedI+fkm+tMG+aEkGHdiCG+Lum3Vf5699x8Gx+rXfVeGIDRXyxnF6kz8M+9R9fEaJ
ug0Pgl1EblJ1KhDAgmyllpbY9xvAwtO5Xgs2P9/ljk01jm7z0xe4uK4h3XDMrK258Qpa5Ez3B2dC
ajVNFGpdZKBh/A9tlyp6yk1Q42Qry29DG0n0yHg46Toalm8BMkgGAiEj+jpPE2TlyHK4xHJx84vf
v6qwfiWcolDJHm7LUf6M4/CXZstyGZ5hYso1s76Z7iTDlNBhoyr1QjNIpfFu+bjDqmFHPdjF6d+C
k19zy6TSyFVj5BWOx2AQzFoL/fmuKT585SNsX4fVuBfdyrMG/ePAIdIfKDzuzuugWbdUgXPSX0HS
QT+Wb6Wi9I8DCJr74oq1fN/mb3UHNlY6DvtC7ZjbjOrcDwNVKOvufIeS0TUHZAY1I07oEtF+ZG7b
8ZtS5mztRijkIXhlrjb3WVIIXc8sdUH7V2jqBDtXhIjHDrG4ZcZq+vZ0Kg71j489GbitNH5dBpH7
S6BHM+BzAeriSQnT7ED7r4AUyM237TS51e42Y6cYFnnoGz+oIDdnG+SpO/2eEAU7SBUadIKiseQM
7bvaFXbYXqkLZghM5mL/JIY2jRUcvpjle7ppK37od1+gNwrFPFXaDI94lmNPmS0Tc9KOIVh4hBxc
cqYsS94xfk9njHMbcueY07iJylW1XT92P5OzKxd/SI6WfHJlUc42IHrIUWJDDHzsd+dnLnpTBg8x
G3Vl2dfm6L4bmrcmRMIqk0dsTipbyNPNf1LkK3MVKtrw4w60rNdUnlsM4mFzzBMoYhD0jBCKvV2x
bdUN/BhsNSToEG59OQa9tb7bOE0mIjtAhSXdNr3PfJUOQMdDBG/ZpjyA+4yRDFfJfWgUi+AJhNQQ
uwPKNjMK0T72VC/m0vTAYBbc19Gn/t3z9UAtBNRyOWBGIUUKVd9pub1Rw5VRZRt7wZll5oXgJHe8
DBg0mau1+ZeksBbb8kv530tvP/1qIJAaZsdL8/RBlKumYruYdXtqBg6je6/CYsjlpYAELp20Jpfg
KigjNIRlo3ICc+UszJ8oOef7JJyo//gW+NlXFms+GsYrzXRx7/003eONDF0rmi638A2TzC1jlsDV
f8jotYff0RVFsyQ/9d2a8FfvzQyc2hqxrQOHbp6MDFtQ4Iu8cMu4EwQ3tPy+tY1j8lwmGlcJL+Zx
bQ1Umb2AraZeEO0EBz5aE50+RT2InrK/NlmBfad1akvwkd0YNARymkkT2I6U/tsvy2J29iAVik0C
54FBZxlCrBVNIzmBMHLFohYMTovnK82Wjt6MHkV6TZ0s9I8mYg2raE6gJUXrta6WmWdHTomtdCWA
r07xAdmoA7vGpt4cbhB1XV4KxMNEyzDHKaELFD3YNbjR1SsiXX+BlbDysxX6VYvu3JqjWOgW/4Ew
yQT11HQdaEBVHHdiKQS2FOU3Dazp5r5HAOcBXK2Zdfyrln1JNKhg8cT7L9/dbL15SaNaCcJUnzFR
mhji24q8jeUzx9SjCNSjCXvq0TvstiNY8v9cFice59xAXbrl/RNoww2lpnQNdA7S3OvU3UwszJqn
ZpqKjykQBk/nZl85cZHa+vu2ITMORpWvdWf2Hwkfs1J0h6XiSaePDaWsOWYeAmbhfWhzvGP6RYC4
5GjmN6d/H6hcyJwmtqvStAe3dEFsnq+xGEx7ksmckzmQTRJUS0a7psCH05j1iEWjdh438NV5MDrn
3xE9BfKxcoCBzMpTXSGP9Q2V7HGz0EpcBnPAf8pjy4jQ02I2YuJSSJZT4odrt7kwQUFQaVxzwC8w
7uUa9p9K/TdlT+tyJ4WGLWaU4Tl4CCCIpaXr+zpI1wyhwJ/JFNkZ0w5YncAak+a5YfPtZ/0TeCYC
/z6UFdYNxakP+VLfY44qvcaAZl98e6TICWVQtCCWV9IGWTwDCjGNrwKRbNL0K4plaj6d88hxr5GD
jP4y3154RMQvXv3/LksFaP5xh4NN+uP4/tpoRCIrFOUFOvXgLgoYy9sGbbCCaxDPJ4OG0zDvxH/T
6riXEa+PUbAz6hZpE2ALFldUURwu9XQ4Dp0Dp5Tu1Mc+yeOgyuIjDIGyyR3zMBH2ni2TptcPuEKx
76hfBFIYZtTZ2WnBTtYZ9Zenu1fp0QeV/j3HhnDOybX6leaKPj8y+/qRouZuX8+/TPuJCad8hfpU
AOxaNNVRVDhwwBItGtC5MVvrD8CngocgbPc2JZQzpSk6x+ifaQISaOW9PpNV0oOgnngKSu7x1IrY
s0Z14GjiQ1jHGyuqRj2fyGtqofRb56K+3cNfUJ3AgV3AgBHWpKTM13mFkfTajVonU9G4Z18cQ69s
Rvx4XEVHurWJ5nAaS0tmfItI81DLN34Bi7T2+JaGnXQnn4KCnu9dZcm42TZ5ca9hfWNGK2ImraqR
Ggyup3mzDcI8kDdCXWohDdAGt8K9RPRBgz+X7sHX+HoHTXFbZtQV+FB78NnP2TEyXAQi2xxbpCyo
pR6MV57fJ1sVzD7iPZHDVpZQZRXD8HLzp0SADIm+GJqnWBTEzbnBXiurm0saatl9YjpOKjymMHkz
v9BLaMyCWKi6j1ifhZFP0r/WkY8t168WF0tDA5k/l4mbc22A9ejKSpqly2nLYMfXz8Tq1NQg+8QC
rD17+TJEb+APIWfqdopE+4VHokDRshhFCTnlQh0VuwIdx5vAoyXy4T+BQlZhwT9vOveA6t/Ut1et
iWs+zyYPiom4tq12yncm+6r9khULFOcpA3cPxn9Jl+V7Qwjs3w28Xz+/UAC7gH3VOZUb3zX3j/y4
8SVvgdtvSYylbfGeX19IvXj9zBDbMSHvZj7D/G+vqwnDdD/eNHAeuZqud7t2ll8u00nq8PRFtdK8
rpioXkd3uq8wGA1hTetRsPlITR3QKXnwlQunNB83ofQJT9iEuSOJmoXNuH0Ti1mBdocvEErqQRFH
FDtGiDaOvNueG56oZ4yrbqcsIpChiUYE3uQyzs4ECd/rTnupDIPzC12RdAfiIq79NAVncZosrpzY
KZ2uknzv8ZjCFwzgPQwi7M1wr0wn06l4e0dp2mVYnN/oBBX9SJUfbYbI78yhSJ6/pSPwTspPqmJa
Fmctn+OP0x5UDyTVMw+ISUTC32lSDhITRP38nTk7tXKSg+LDdMF90RKsCOyfNG85VNtuglh3peWn
bKztMk+atMuC/AS0//9CNdH8xgm7/lTqXDIK1BqGPd/4fvqz8EYvCaef3L4UQsVR0Vk9aaloTt3Y
NXLmAw+vXo2bDHxpeBNCBNPvrKdhCH0XFuu4flbv+WXmUYZB6cabtu5hwIg6oWjUBlRCeXejR41t
aG8h8VeSCNrtZb3KK9Bvv1YXzdoWKxGH1xfmTzeOZ4aVYt5jWcdFSCQVnwMRk1gk2oJhrhyq0Xe4
OwTDpGQTHvJSK02VtFswDKzN1Zw/lw00d0ODhrl4FPmscCMEQhGguJKjFjYjnnCwdgIlkR1uQ2/F
tzRvW1/gXmQDtIvCDx4GZgGOvfAfK933GKT4X9d2QwU+wuS+69j85A+IhCYpRxoKnObw3l3se330
ascYDxHWZAZhHdl//8hwv77c8CA5F9FGU7GAQHO/PM51/SjQAUTmLF8ByNEkoYJtE6HUgjNOrsXn
WDRkYDU2+vZEz7PHALGDqnFHzifHWmuc5f8ONsiL252ecYRwgn50QoYz1bhbfbHh0hapLw/nnLGc
PTAKx91K1gXmgTzAZYe4Oz+rmDRmwPIDTRLPsDQhIaRp0ppa8piNCpyOYyAPOhceBsyfRs+btHah
VPBfG/FnIm9SPee5pbdxLNPILxYnxVlpty6AzkSiW25CdW4HoPwcRX63wiNfC4Rs+afWwI04p6Mn
5t4l3BZJJxnWPMoyo1eDsz/RwoeCprxiFvhkP+/YI0ZAZBWoaE6plNYIh26PVOf6xTdX+aNEERgM
r9t+7Js/eX9/XILU1zBxliUaxMQnqjzbw3ifW7cJ1KvEPN06NOetLnuWmF/2qAN959nLimIUCfx3
3r0racqRV4R8K1hvWeaOIGnIMM6Ll1q5eKd5xSI9mSfDoWrti+t9JjIVEmLZ8g292b44d8rUZ+TS
2SK/03YhxvsRNcXg1Jh7jWeJGYLc++b3eNezBMXkN7x4WyminP4fWKsLaY1tYZKO7RCW8kAKXB6Q
rIIRXUtoGbOjiY/96loawLPFIZ2jBhu1B4AUphGYb6RWNWZAUNpvh8Pg4l/CCghSpoeiTIJPEl9t
Et6Dm1wCuTNZ6vB8CeDF9kl6n2xpoZ1k/4aLINRsur6E+yT0+Afi5NbqtEI7Y0NcSH9APlvMf4Bv
2Raaj5AQN5hzgXE+mo9g9Lq+V+Oop2pUfCW9mX6BI+LhuELqCR0appEPKHMky51HwzEXm0rZ2gBq
C1xdrANDced7Fq4w5uanLeIT0LWR571GqyzEgChesprrpeWIfnaQzCSX+fePEkS2cY1um05/YL7z
9Z4M05twhh8POm/otOxdn5ujqzUU7/Q6jqC/IJrcHrc0GVS99/C/anZq/FJpgaMGGWTp+/AflRC+
HGAxTGuF58e95bl6O+70hZRl29uFfCH4Qf0KrA3Zs8ZbvoaZRLACCCM72cdkQtnvYuGD42ejw1U5
i3jxmn7GwtC3v/sSVZtwRQuCCozcp2TPucJkAMKRwbV09MweLy6BKdorR9Ju0UFJ2gW69hsiqFke
Qx4Y1Ji7SeKhIRHpjEVjo2SYGQo5EAZ1E+I0fOXhGYIflx8MyntVb16RMnXQLlGam+AbfE4wzHfn
9NzC9GkuMwIy9XlVs4nHWlqaz2rmyheXdxV67q5hnGLMbvkjie3FUnaXYIUy05++kLGDuHFSwiqz
TEkhCbvv9rIwuF1HIlJ+sdaGRj53r2SqCh52vsI8oSirnJkz8GnUu+qSKsFKV12N7PrUW+asXfAN
bacQEggLuwoVXc/Ikd3ZfQdCWxxnW8QAoHBsiyLbHcAj//E4uMo4L8FuTF8CbsDHiRXS+gAlYGQ5
RuIg0c1BrKj9AdSfbBESoAecSMfrpp9OMCTSfMuIjdzyoOXvaaUm4xNTbuHZGHW00ZWxIiH84N7Z
2j43u/y/bqtOlV0N7yka5pDkq2Y4ENW+9rKD4XD5uiViKApo1Cfr6VeaRNtJGyY3BCq5JcZy6sqU
/TNwcVqebdlKU/jhFELxrFb/SGLLl1xAKdVCNPqH6/+nLUwaKY+DQ3VXfRJdC6SL+9L3GYlSS8sg
hUWiaA7DnkHQAbWDkuBxwpkr5Zt43cmKoN9AX7dyDqTYgrD//rfdI6FC+Yg8SFUJG0kego0jJbi+
5L2TxPzUj8jXuaRgHdNgPIJEUdjAPEw3eLOEdmNKuM6u9JsvKybX8m06wb32LzSeJw5Oio8BeQ1+
A80gtUhpG0jchhy2jYtPxbGEBn3PfNTCBkJSy6xAt85m7ZqCpVI5Ti9Rgq88I7eLXYDjosmfV4O1
WsonSyxYsZXx/WNdRizpYhd8hVG5AahIZ//TiLFnxSPxgCZVSvK1+5AVxrkWp+nVy/NyZVDm4Jf6
jolkdDPclWsSrNeTiFGtQNfYE4NHuiqJm8V8L39bNKmSBPe70u+NDTz5bbPTbcBBW1y+H7pZlTVY
DmJeZxQ2us3Ym8tf5IXooqKUmYb/ao/JvbPKl9+GR4azhmxfZub+ZYGlMGebVgxeW3XFWzFC9QY3
5ToCY5d6d1VIotQqN0HQ8HRiWz4irLOmF1/+r9ZE9zLmzLScsRPaFMiNIlLBSsK4wBt/BDaeqnK+
HA6CIqKUi0vA1mhTjpCgBBQ2UtkrdcZdAdV3vczi7o2A1SFcvSK8nrOhoqZDh40O3ZnyLfEMKwz4
F2iFLqnZMV8a9gdGUcPyzeRuQoV74AFppaBWIwSbLjGCE4G0rJKsbEr9MPzUpnrCv+qEPo5E8edn
x/ie0VpqqSySIxW3UeTsAxNhkSyYmS6bq0y8Dro15C7lop1wXy+zgZbA70OVD7ry5AnI7xqUqsjx
RxXirAhExLCxApYwMUjrDYmYk2oP0ZV0RZAZYJfbN4Xtk6zHbEQiVw+NYqCjbJegU+L1KV7tDlqq
XreW3i0nzCj9SdL+TqTTqTQpyBBQ29dBMj9ADOpNzJ30O2XWHoCNain/in5tAd112gAjF7667uMN
gJ12ufebjoDUw59HgJGu8oA9x1E+6KTMjPMX3/R5QPPMhqinf2/RtX/3dGOBuIRyNJ7nxUd2Fiko
VmutieglKGLtzI67mY2EYCNnZm/G0fEg3tCuc3zvhyUkFMVZLD8ysg4ZSPJj6g8cEaWsR3lhrIo7
Z2AYcqCuEGBRMeWVTIWSDrq6ZNyCMiAHJEGN6v2D8HDTxGt9kQH034yhzC+f9dRF+kJxMmR0vpTt
T/bYzG++fy1KHAzt8Et2f0zZuzMaTnU/Hwt23SMqktHEIMpN9ETp0viW7LuwxVEocehVT32ZxyO/
6YJpmTgMC/2Bhfdc1gtafMPcF5gRSXnKtyFHfrJIUfoLXo4+KoNcaGkjIFqtIzfzD0idh4YUvxJr
Bqm7h6F1dIgwiqVcG0ppaudpqpp8xfQZyVIAJQZFEKfIQJhZ3EZxf79PY8wzhiJNPZwkZQrgWNKy
c/gVUC965zz5f9C30hwB5KMKfQEU8nWHa5Y+rP36Ecu25yE+Pw3ttFvfbVDz9sCu1OUoMXKUogmH
xyA5JnHmENzw3VGeHWTZOJA4Bmqp0Zo/jwVaqRRUYYgMD0ws1bLPxXZF6zG0Pnv0mt7qJtN0tgI2
1yX8xWUNyPkwyCw4BDhIEyyxgscbicVERrb7EnuhQaqgV5vZ97PIfcpCobdPJGZBucp5L0wr+PMI
D7Dg9d+46K/uEgd7oHp+ziUCBWcsv6wkU3lVnUm9pTWR2TuupnLZm9XU4r5wdmPCi5RLsmx1k0m2
xQobFH4p/XT28o35p5aScnqovVzVrPYXD4bI2WkzZ2BiRQyWsFVLxlMgzHBiD1NaQAMZR0xY39Bl
nrtfHqseTIYEqMu4/H/A1eZOSnpE1Tixr4cSvh0RnxMVCsyWq+ovJPbzYGn34Vb+5MoLePAsJOQ9
vBBcSEuWBtEJ7tbDXL7ZLDk51db0FoJRxYicqnM+SZd7dgBiXt79tlRtZt3VH4EB9t4E8tz+uNol
qWgPDGP8+fRxzBBa8Cou53o5uY+jxYGO9BMgLUbN+BFwvW+Ojv6T563KoxkURli3UCahg3Ws2aL+
Es7OsakCJ9jp6mxXzm60MVHRYyskGB6RALA9frLO63RhCvkUE6Dpyw814Bt/FiyTjven2pc2uqyj
6zUDgHhG8KJ4y6N1u/OeKoPNjCdtSVJfGtIC2u3WKcSk05VBxofMVsJo+zqYRgMib7ow0JzYEOvf
uO0o2zwijyOqUzaEtrIJESVl0Ej84DfQhJviw2h2qKdv05XJhiLc5DQlhl6oPeLUDghezFIVwg2l
9UoYV5cEChRfrqy07F+HDheABBz8XmTKjhBKUkdn9aWRASgmMjkb7+OyasZrlKF/vNoDrQ1xUwPu
s0ykbmxmKves3td1PZ6a7Z6+XaX4KXL4JZ5iU1rpL5PDCZMgbj5Fl650XfR9Aug85wp4fP6MHUNu
yX3A9A53skjxy+wL+tB0kCuGycYGO5SxPJeHmFu5qv2RtyFGATUR+lLgE7tzF+IlcrIVga2GRkPz
j5BN72/biTm2MvFEE3if66hGhadYB4JSNGllQh1OHIDqab0x6JGoBYibnBwFhIrEzGvk2QDAr3er
+rGZy08kqn4zUs7KXVvG9Z5HdpgN6JFuni94AvCwnvsXSj1SMEp0BE3fLLbpVDsgE0nuLx+YOH2v
InVshhg/cEWD8AZ5fA0vFME1jZynLPtt0x8E27tRq/hYXlDfz9amBsKx33jLQxA3ScyYNZT+36xy
04CG084+9d2luEMOUj1STFkr/U+pcA/TJuxgsBQArFeOH5sM0ULLdkbUVZmmAhuLFrzGkPX9E8VR
Mu2eNZQJfUP7YFwvSc1CASbO38zoW/vIM/5pJYet0DI692zroOep0497Ad5Bm416CO2Tf0gDgYBZ
gKL4pHmsJSpwIKrbVV9RG/55AdIxktNxPbhvTPEcD+96nnLgpPIAxGL6QP46FopmmLeiMBOr2gbN
ofAS/fUVT6WLkP9bdbuId6lroO3LKCCtR+qZPCz5uy2aqAOUx8B8BOmbM3BxeawdMwEOHmpOQqFl
W2HPA2kUFmD5LSmouodY9L2spL6bqfBX1MzhRshUURKUxldHEz6qf0lYzHQ6QU/m7uE5ll+WSDa8
IB0zyTKBWOe4vKQ9TKJ2ttonk4XWLKfTTftVIlUCa7gTvj3exfL+0U4jo2abvzW+1DvGxsBdumxW
zalgoqZTqlYEC6napFFimmmJEcLSdurTITR7u023j02Kgm9yvgKBpjKQ2b9nCpHsxRfARkS2Mgtc
yrnVALHww8GKaMrCCKyXcjWduu+whUTkPgVtJOnQj4F0Z8wGRNX91o/eeYsDlnMRTPOwGJZ/uhF1
C+bOnk1rOCFNcbqKcr89J40FzvzU63wBLODR/kpTWHBrn7Mpo5ekSEc2uqKI6NfVLwsWXlaYZ3zt
qEP8O7v8PMV4Nq3/0rZWaveV1neXAy010eM+Rylr00kx/d/aCp2U+cHxJxwsompVXXbAy6YA4TN+
cnrLObM297+HOsLJS5zI7uQGPMJH2QWMvL5t4BpAbDTd16aL3QtRpDzOpIUeuzxO26oCEXDYwLyY
wKbdB40XuZFGsjQ9d5wbsyMZnP/r4GM3dPfXxsE1yxdteQ6whO9lmP9ZZQwvsVnEg9F4GuDMncgB
/OLKjksN0SbutR7W1Mlij4VLIJt89W+nmUQytjkzTI/LWRFcTIO+eqqd9uzk0kyOoRrQUZfIZxND
U4Nck7A4orjfmUG264cAvMPkhIinZU574qs7+Xt6uOplbmbXz9NML0GKTJQEw+dmYjemQB00e6nM
hQT84o32adzzynaBbIIdtYoNILwDRe1lc7JOtfwvfrdvDmQhBE+G8NObs4aEUEgv8vZx02qWWfw3
7hoYgJ6nUWo1VKIN4YWrByZDiwQHBDWM/xqoIUz0VhggHb23yWECVgRSHf+4zgUQ+hz8PvsOMpGN
n4FGSPWAesc6JjC/trwgds3SdO3Cqb2YAm+hrEJMV1vfg77YRbSy345KJO8txefaDDB/D4mmFMIv
oBUldmGDSU4Avm+UlXYohlYOyeEXXn1VDhLuLKYZ5eFlaCvJvtM/oWTqeR8DcULFdSoSDaLTGh18
Py4a7gICcGoJHBOmkI/374xCjGxdYR5vY4mLubaJht9GtaOIBZ87VssFnQdk6EfCtE/BviQBVL0g
PsuOPnfCufOBOAcTm2mkPCr1IT4GJo7zYvPIC8aO9TrflCLopg4WmFe0q+EeurYk/M4SBHSkfILu
Tz09yNrOFeoKrDdGO24n7mqm4ielhpgCZRlZPrVx0ew1s8cb9zCLgPho94/g84mdt6gSj19FKpVa
dJ716ZXhPou55YlIhIEmkGMjSUI/9vAT3YFXvshHWZCpxAtztxphk+13eHREyT/odBCdfdVjD6uV
7yI8f5kQtHcjJpFE2B9j4XzUijgEFbcC63vEejbr/bqafrrOCFTk9HbyGYSdcUPNjCa8stcKgr4K
8gaCiGn/1KB0r+n2plzHq2ibbJFVVB2PEWKUE14M2/SN7lobn1/4Ww7TWOnrZpMtqtHVa20GJwES
K88429NQRfNV4KENt4H/MjOi9o8p7h4ttIT/YDgCZ3GfJXO1t5wjEkXSINQNOeJc3amVoHViE5Ja
wI/txBs5W1MMTb3p3arpmmmtUtxwC8Mg7VxYcSqRQ8S4cWjM9Dq31aC72HLz0pcoP0hAqm0f5ssc
obSsauV6KxsAcWIEwzxsFRTuYartffbcyaFmmwA0b4+LSlY7vZITAueu0KsPYQMhOkvabvM+7E3y
phjmSNMBd9LDrmWYV6QP+PykbGuOAj0jEIAwX6uQMpI0HOAvxo/9crWEj8Cn77f6PghCbeI4zNJx
qDHKV9iKBY7ziNxdflyf4nIQIu93Gc7oO7LXdBrjD+e8kSQKsd3nwuYNwb4DzrF/bI1p2jLLhRly
vCZ9ibnK/KaMfFc4XyqC2BTgNyuum0USWe1pqAQ/t4fPBVBTszZGOoCTpF01xxXYRjGUhwr9hXwp
NJSEW75lqBT4DpgBaH2/y45AWTQrO1ncwE8IVuhQq1HrgIUKpJxPiGUWe2Cx6esk539Q936PJLYn
Zw2ZX+AkDrCPOfs0C6Dy0TIPPzvDCZEfaNO+OyClPMMzAX6yMlFvXxZV7mjKi+2OWj0Zbw9ZNPmp
9wBemPsItVr4q1LEh82AZtDXAooZfI733mvlhBdrFgX2REN/tI4MZCaew+Kr6gp0a1NJk8Pi0ftV
dVTkwQhJdhkyZCmvAwqGn2fXuwJg3YPksRUEvc/ln10fxuqoUUsT4vG0n2gV7tppO6v01VUya5fA
hGSkFRl1ukJZJmgDqYef2z82/xMeMjk8DggAwfJTowpurJA37MJZ3zMg6oRGkE98H/vm80Db9koK
gOwSr/sp45iq0drvzlalHQiXLCn1pt07xda5+tG5gvuDOJUKD0lQUzYMLEr3LYZvluakHymDKjWi
sTP5C6651lZgyz9kCeGFyUuMw/h1FbKvcIBcABwtDJM2Ivfyc2wsfvZs9ud0kC7ImRR5/anDl3oB
8562jB63kLk7rYRz5TUJF+APpWiErlhyOF3AwrD9m88oBt83GJkm3yQgZy6JvqTG8ZrmV8JVKMg9
iHeUYnKswq51KGmCDMEYjDeaxBF7bC3mYVO11doIwxAX7OWCmxqSFnOOPx2YmeSwVHSNiuWFC+DL
8o63isEvkX8L9y5Hy3rno1jafmsmKB9mfBzpf2kkEiOy5aOvc2jrFMvkOGv21FFXX43HnnUeAZ4W
KsuiweYP94A3x1SAtLpcjZvNJG1DVPPP9yku5Za2JMIyKUs2NLGsFuVlr1MlRf64eHy83wm2gOMZ
XzYUPTyOE7+cfcYdeyXW8MLpBM/yZOLR/xs/zMXBNyI7R+2vhAh46jVbo5+jZizWiOlyQZhJHHfR
RjWdC5xHqfdVf5yXVlg/JtCMS0Var25prKNxGf58dH6lknKHIBuCilwSdi86moLoO8s8rdR79MiW
WDeQcGxWnQlaTJJ6c/KFN/9XwcKTFMmyHzvdBvMsjGbtDcfTYqQ2KjY/C3XGC4iBKkRMemnx7Njl
iMTVPcBqf51xYRMMtmyr9YjDuXSL+xwVhNzNrQM0ggsMXO3k4DcwRb5p7Bg3CPBcvjrwCBH8lCO9
ZR2GANKdlsxm73jvOavughPFqnSWidZqjsHy1pmQt7vritI824PBQOISdy/9WcS8M96dhRT/hRVV
Qm/J9dViFiEP8zWXO8aAPT+MOhEzEzpMo3CKE8+9oiEfvanqbbtKbNa/jiWwpmy0zD5kBSJzARXt
DVT2Rt4F8Y7eo8KsSEGlfgGbpqFdFsokUSttvRExjRG5roaYQEUJMMyXAfN9Ush9l2pK1KhtAt5Y
XrzzExM7OjtSNrNY5WqpdW3qSuZRR2KgfWuXpTLUeSdqZ2xtWospJ7eIxFdmxuqTT9QFs/d89pD0
oT5ET7pnyA+fAoIsKnbNP4Vel9ZQk7jxMDlBA/KEf0Nt70kKgj7/23ZL+5hYbjTPKLeLzbG3Iuet
HrYcCNLn6nYLKap2BsBzRAb8CMVnxXIp8hIs4R1E13MyANiN8RhDn/aKSDCdwqQCgNgH1/ZZVWg7
mLa8YborzNDSrSm+XRqOmbD3+8gyDSlGwBncLoQ3Qmt6G3wvfSXHvHukvSW6jF+O49CleK+Cxark
S068SHRys6pKKsIWvRF2DP9n/VS3lSTN7cSYYM6v0nKgcRU6y9QE3xXNmc4MxtmxHCW7AHYWsUOU
gvJInr+zlrUcBf5gSM6BbV5PSIBT1YgSzqRHERAOd7mqpaE7NSuZEQPK9Ca+I7lIK9uJXfdajzdX
jKrmB5CzZ5tRxGPXcdu8xhhxuHgH/3j0/bmu6Mhv+j8bTd5DYhLJwqz2mdFfJFMe17UJfXEnXe9p
lECY2zTQI7thFCy5wRBkhCmZOtTlKX3o/APJjlA+GP1D2PMJct0fmW/UvSp6RQPUY2PazYgBL3ho
0cj6i1CzfxwfxhmTqakBN/T2iy4zcdD3r0FIxoM6jue8t4L9VfJ3tUswNJCmGytXo5Wf0jIUudhd
te0Mk5Lzb23VhUTwkYyli/6amkD4Vx/alOhbifPH9tQuP6xWfYEXdt9EyKMM7l2k+OFb9FScehX4
xZvRJuNqxyv1m9EDFeioaj2tfn6Xx+wX2D+kvTIdh3tyTk5bMS8qz/e9wS+1tzH73UFvAb3bkgNS
tkWpODuoaaPEWXHqcfM2C446QeASWUqy/5Rd5CH1vFnuRy11UD+d/0Xc/qBTRov7Db8o8j5ZkxwZ
4d5dckD+Hp7uiP9vox+D67dSf0hLGk7hq7nqz9sMIhnLykuvjNTEsnvFyMffuH3KaJFM4BhIBCSR
rX7+Y9wjQ9JPByJ21ErLa0hyAq+DW/hy/aJKxfrEbBi+X7wRaCTTCFEZJOhAGoY76XJvF6eqY1Lu
DYOhNNjKQnp2dQFrEA1zL8+l2xwfZe99XUCxd/VdNqmGaXGBujWmVj6vQAgJWuT2HIveg1PvJIhI
MT388lSnjW57GczCgd2j90QZbJcTcLrwDLgV3Tp22l+VXJ9QnkamGq3OHVYveKXnRd8VjbqHDWno
vAcy+YZwwBpThTeILJnYGZ9ZruPtlcXQhtFsELqQrZpz7CRpUnOkpap3UDJx10Hm//wl6hVwmSpS
Yo8RFN9BV79NfzE4cUmcjOwPuqs4E30LhK/3rQzL47P+TXGHAkY47OQHKfI7/uCvPhwQCGkMeEdw
FDRpDBgjSVUFAXFRlaRQFazMFp2VpfXcDqdjciVymTDscbDhv92ry22fHfbe+LFN8MqcUKbyIbX2
0g3LUS+j21awY+Y6RhxXSkuWwMZiKau0D7wr0DGE1kW5zmoj008foaTxsSOTOnrczu/iJftatrUd
Pi9FkCfoAuPC6jtIuFFsGVssJLxVQAk3xc1MhFgVILq2XjIGiKj8cXykwR0l0eVm1EbizpWO7XfS
DBZYqIrdnU6yjkuJTQ/AGiasTfGcU0K3lumLfA3rlASgzsC/gqAIVw9RUE6IIsyhM9F9UWUtKDYr
dDDDg1UwMgOrMs7v6YwwKcGk+tEdL6owfeDTJRRZxS/4BycG4aqWhO3nCQmI1OZxPpCPyrsjQlQ4
Ms6ZVniKuGFj204TYr4/eUM9WFV24B6QthogUr8S8fK1GZ0oJxDs8jVvmeIYQ+zd/dqqBUwdxfWK
SiK8OZUdh+RTl7jWLwyIOAavZiBRhUl0aB+lq/KXDrAKqLEf1JCvmuyxExrtDIgopDP4ebA3ECzq
ePDxjIXvhu9Y/q8zx+pWcgDxKQBZH2RlMybHEwrw7Eu3xRppuFbOFeFNg/74z39QhX3iwkTs5Eb0
5GqA/OprW9qwkNLYeg0rTNwZVK2KedY7+mu69HXFGcgpjt01D8WhJyDXR8kshkHQwPU/FMyq8x20
GOIb0P79u2UW77KZgAuVRAguWo4FDbQQiBP9Cws5yF6g68jvG1aRWAQa5VADM9yHOxIwUwBAt/Yf
Va+Eh37HfZuIhSrxJmnlVD0oqx0V04pVvbxgKfiiTbGY/YDavKJtoTXIHkkbt8WOV7NIUW+16Wp6
UGxxBa4w0fETSrxdXtmEce7yGfsKBKZhmSmuOWRt9dqH4HCiCQGSbsQTJfrODQZkrP4BjJsBGEWU
uhE9zayD8rGKnzrakF0x0dNAgkG1OKV4BLpZ48gmRLnCR3LMLtvBLcdrl/wsPl2QV8ucNWVpcR7E
bBk5Y6B3uzIjFzE3B4TZ1gr6oeWbqhledbeLX3SQisUFeImTNC+ojBVIRPduiz3d/+o5fsEBZTO5
J0Jh70vL0Gn3TAA1IZuuqrhaJXjhBxanmjvcUDRztPjsR/GDtEzNMfnHHFPnfa8i6DrVcFOjut5f
SUAz0sO9XA2+QbM3nqUKUQwpjvA5xev61AwZF2tO0Wt0FfA66YmHbsXnVLNbKhttTZUegCjeTheC
ergKwYJML486mo2Sc30IElYdrf0qLCxWrIE36BZ/6jFmLQQPwnlh+7qSYEfa96h32Amq6GqWIvjB
lpVNsUlp8dmkXNAiK3YlrED9sYu10n43XeVkTWG5VmPPJqgP8prFIfIwhtK8UYdA+a7heS1/2AWB
pYKBRS71RA25LW91EFdRlQA6Udj8p/l2zgQhCe9A3KVg/Ov+FJxnqDSQt6H1iq89nGUvZhACOMKP
creTe123N7e6irUpzzV2J/rjwr6c8iNDQi9VCQfVQSHw9jPI6fSAGN6TIaqBk2GgKzlh6rFJHE3Q
dnNCjFYcmxASTkzUVbV9BOt39EmhD7kLPv9IAVwxD5d+/TZqikSV7qLBTRWLRXNCQ0V+1CJsGV03
ZfNrhXUQNreTCh4BmHagbbPPyOd70eAPrG2oYKRzvOhvv97qBoOrPT8u6yMHVhPh1KlE87m67HtA
M+EBuWkYxU06LQvcBqL0UQZLwh+EuZ44cPODdWfQqilUF86klTNcD4pXgU2+P/gFYSJHms8Pyfm1
lAubTzHcCNXNmecNdUC34Po8KsvrFAcGxmckrNiehBWeXSfjp4ICyilEF0QygpbiivaIvHJBUu6c
5z+5qJ4uW+Is6/GuvfWTVBNG/1uIVQcybFvfuHhfTk+T8U6vM8m5n2tGVhAn7NeP65bDwEai20G2
1dwwSLMuVgJaH9pvRwRFyH10fUVGm080rXG9NJUWrT8tEa4pGC8QS1q2fZLszR4ey4a3xcS7Ba3K
Vk6P6P+f2Eua7ujilXCOezeWZrwpqMRqWOezxx0ydH5zbro2CcWTFQd4eHJiv5PEM4twIgY83oKG
z/CYONuO51CUMk1ybk24sJ0SyTAeltOX3l5E//NtQwIQWiDDYQobvtz943CeAAF2HsEh6u9Bwm+k
8N99w6f3s2TetgxVb6908QF1KTtgw1GicukvOw45G6iqMw3L+PFY1ZmBlfBwwAdJDrBjBRaXLqmH
Rl7ntluP8nZKJsKp6fZ7DwfACJkH+rVCh4QdGu0JrJF1BjF6aFHobNWLJeQMdcyy54nHCMvcsUdE
pD1uVaeIQd9uF7ZGSvsZJA0JTIyWLmuHkfIt3l7oygixbECwQQQp0TteBLVlKyv8nJWcdHcKTuWt
Yk3uf4s8MGeRpxJL8xtMJoFfymcZMEC0MXqE5XcQXRyUC9ZQ8/lEZbwR+Erb4GMtDROSXLUkfYPm
UmSShliIt1B/2AM3Z3k+CmVxeSx8LpleZW1MOM7j1knjBdFOOTuIDK0JTWPKP7MAMA/xx7Axh1VI
pM5NMPiWGHgQvsqAoFvsouty5khavUOxIanQEGVRsZqy9QzVmwA0GvPpfjy97KYaT/trjckIlfQe
QgssrpSVa8irP+ZDkrTupOXRtN4eK+Jn1jtT4Qi6KCTqM2eWKFNKsQXJEPCt45JA+8FLRXom1sTC
xmxECKxAVYfUlNzbW2FX2dI78ho76//DAk6rgcYNqdAS1QJ0Od0ofa74J6TBuqDMG0tuedch6zX9
dnO9zQ0AzDC8LWGv+csLaaeyXgMAG1KsJAeaYXkJ2w6Qu9SG0AGfbb3BtilstPQNZrZkTcqjggpr
i4J9f6+ED4QWbCzRTDWhb/mBQwdO3oC+TD2mywAAqPFnAXjW7GF2qpjJh0K7ETNen+EMGLw85WVs
YDw4WQK5T7KyRc93G0OyBhjcZOcHhdqXy4QmM01JQFSGrKb6bbWyj4atorSz0IV9XLMb5KQzOVAs
bH02L2RonH90P7l7cvkybRZp/9FXrthzATKmmUuOIFjiKk9IDCMJXb6Riq6sYprXIaqAkT91SHEf
Vj307q21d1vr3kRDTJCHibNWptrRPf7CowUm0/G3GzxMeGq+5Ezp8Tyb6jXsxgOPXZNN+SdoKQ5o
zczMZSeE5ycfV8KjefYZNJfTvaMlQvclxhCxRNMgrxpvTgaO9wSlLwHdUeeWvatQXs/WOnITpRR0
reYmyvrL2Lcq0gJiD/XQenkArhesVjvBZvpJ5hIHnSrkLn8njA9k/nNXMCC+fgv7rezobLX3Q+fg
5a8ysGnbJ24Bd+ytseMuFpSvDLBiPNTcV3umaNX79wopqOEuPppt60cjkKvzHWGIZYtCo2AbOaPL
31uNfitFezbllk2WuKKNAmICwKgE7lZI/yFHTQhGXKA96m61pLy4Ij+WiDYk9r5+QjLSqsIVv5oP
j6J4HqSLsr3N5bktfjlJYkGSYN5KslHDRlCEyk1inhSOgBK5BP7xtTbIGJLheF75mJ5YMvHvsDlr
9mZU3jWPAHam/7BDSXG2MLHH6LGwAJHtg4pBkSkwcExHJUeLx7+JWUoNKbJ2D61swCV3nqUs2wfO
OIjBoT0CK7ap5GoiT9/32lG0bZ9LBvZxLg9XMb6MHCjG0IeOxPpP82tCal55F/JJuEiONh4JioHv
Iu5t5RzvCo8+4fbI7WCzZwPKKFJ+QfF2UrUlPQJwQqjouMJ4XaEBLuihmejVrKS8WbBUiLNNwudZ
hSp9YD7lN900s9TJulx8rWy8cjlDAiIUQXDQyaPEgl/J0QU8wigeZq3TrlGRdg/kRpBQcJQfFT+6
ur8JnXzNYSnmHe505qP2z/oxwq2E80Kq9x4AEqTP9GG8YJgT5qRAnjOrR293XHCedltBJFr+XHJD
Bu6kb+J0Vl+QQmvb7u9Ycvv6lNiBzIPDX51tr8/Dh1MOTCY3c/kM7C6REDst6/TBhJncEYRqBMqs
CeZGEOqFSWrvIOkSgKlEaxEhAJSIDkNWvSctDKkjNeNOtjMClfgc9tASddIqPkEZxar5ix0a7aGs
KmBmcuCaXVt9H4j1YHJivUH2RQAOXpde0P1ilH0SdH1MugZllto66J2Mzn9d84PsdMfs+bJos1dv
c6NYHtJ0hjGiXJ5zApwsVzX6GJCBDSijU6p+PL+NmsWVdt0z13Crr/ieQMnz2cG37jRRXzA0MsxQ
jQfQoh1h/i3uK0puoicjSKE/+fnuk9wIJYBBa4Gs9It+5+QXO4Qh4+axE717ebfmwEUGYCUlxeiF
EZtsQlrmnor6240xpfG/xvJzmm5WsEuKm1wXPXWeuIKQWKjWlC1DrjdloLI/8hDPxNjW/+UHRc+D
yBy280FWr4U6oZTk+Dqm+Kqkroo2k8z6AY+VLfpVxxivgsPhFuGHDLTPaRF2eboCY1Fd4sGC6MZT
Yd8C/VK1KahEtL4ov03JSRfi111BtKhA7BKUcUbT+FfbQ/g3Oh7ODhDfnnUmiK8I15ysAu8Y7tda
ocllf57FSKXPXTTt4K+AAFIiDuDRTQhygC3p0E1Mk6XiVD4/5CvPqwMzT2XR0N/U5wLOMH8cu1+f
XuUDWTB355B2UBxLWJ0gJMoQGikRmv3msbPxZIPl4Cq6KzOFUqzfz92/scoT0AOzBHOCHxsZQd3f
sss9LtRfnCAQ7I8OmVXaQwp0NurUrNyseWp16hNLaBIcwZcVz0iZDtbK4eNhO0X0g7q6bSNkprJN
t7m03Ez8xxAwLqVEi6QQ2Ux+0asD7PFebNWeqbZYlCCNYHI+o/1Qgp+mlhCCxwiJXLVNWOdVjNQx
2NIMC0cH9cDApxwFOf8nbcZuUujysPSa6SxGByhya+PE0XIFo1EG4wmejwEqoUZlwQyA4RWo6Uqr
zw531Fq1TK9ob+Sxe9fKsObRQ9n01dXvObCE+XhI7XblhzcV5VWMCgll6HnWRgpboCC/Dq1XbgqO
PsEu697Tf9J/Z2CrOkaoPOPbUUtk3FOE5oC/forMjix1IXhDZ1Mj5Sh8ir4a1PENkYhmzcIr/aV4
ycv1gGf6P7hrRK0KVTqIqwl5ZFDCG/7aiBRo7I+I3hEGPzUK4xksMDX0h48Ufy4gLE05HtnyUCuX
ygA26ljmrtFZHWb7zDUrm7td0CvFCeIKsJkJtfTFoO7oM15v03vpfhBJrXJSGQi9b8uhJqNeCZtl
fstF1v3tNhSAGfhRMzY7akGie1pmH6JX311r4/KDit0CpIn/lp0rwwhsoK20zfTXexC1hblTQA1t
Jmc1XgOLzmv802M0zurjVOYLYTB/QyfrP4X2uSp/r0iG2UHiiq1/NYXJxO7SKrIe1BU5GHnWoYKK
Y+R4OJS3eBhMvrHbQG8n0hfgyUT47Nn/IraGx2pVeg+JWbxUVjeeQj1ug8m6Y5Jdwc1Sv08DuI0B
1WYrBiqSklbnt+5eu+XX6OhpxnEbPrjPw8mSN/6PT6oExYd6ZOYvsep4rUdY2dIymoYaM6Qwutf0
1LMSCLvjew7iMO+KeyxvodIrpS2cLEdBKH9DIs0Y/oqulvL1ly0g0EzfLCfntGn1C94xEBdXbUTE
iR7pcFsZsZnmGttQt4zRGSS3tr8hmP7mZu/bRNu+M1U8vn2YiNihnB0olu8rNH+r0gINbF6VJ2Ln
EpClxD7nEwPo7sBz+Cwf9DvuSijKGrtBo0PTDdBGsFnt6AJPCHO/TNu6Oge8IlHqrgxMT/my+Wh3
rqY7RsKo17BmySLlzUjsPT2IUm52dCpkJ1kH9gvP+0mKbb4sF0NECG9R7Ja7Hkh2yCUTbIKyXv7v
m68c4R2lmoApx0SH1P0YEOTjaBMVOrOIBPrmSYc3U9K5mApefF4x577fwCRN+kH4dl+j5HhQiuXI
GUSvSAVpTAJ04YahmvrehEmqlvP4V49iGVaOnlGB3cDZLqSuoy5eOh8JGfBWsontOk3fBV+2GGmN
W7grwXq08Kh2JYjkaPxjLLZnaEcqBmqR+N05x2fIi1ipRzwAySLyG1Bs1nWrVcN7bVxBXIPKiT5P
UPfdh4TXXiYtpK1Ja4LEL1zGuPelfO4VK2jdhKz+hITqG4/VES4t25gISr7nvYNwch13fTWQSzhu
1RIm6huBm4z2FxZol5ipOjUEsTBwMbHCA60fo4UXLYqPBRjwDDO+qweDhAlni7crVHjwvP3gdsDd
bbbiwLWk4fT6bNSK4ANZJVJ/VZqK59WYS1neOHCZ1L3DslvmiGczmz0j73zCJJ3d/1Q7oAssXvi/
s/nty/w9xHvwWfY4SvQmGI2E7nTqa+gpRhp9mL2Hz2CxINqJ6JygzDCXq9kmcatzYfOC3amAdfp2
eFefMuPuonnlVW30srDqnyHsyE81iYGRTrcvwwzvtQTyeCrnkJ2xvADmwz924G+Rr5RAtY+PqTsc
h7BnCjVkojIpD2Sab3YyLSQzZFWfQ4kyCHQsrcvW54/ESZbjfCI6ijnE8TPNn69vY4gO2rtTh1Gh
6TKfPtZOyVzouDvZoqbGdIPbKK9P1KIKnc0JBlV6R9P6+719pw61BBdX5XyLtlDPW4cdYqjaWgb8
Qxx1VBZIygQ2Qmpjjtn7+GOWfz5+9dQLER8hFqZz27SrfD+gPZsdccKPOVCT4NaMNyUo67G8296Y
aEaZ5sSAW1s56dLMFxaRN9dtmWtkJydMvPMq47dG42CTPXaXitF3VAJFshRbUc05KTxwcQhsmMx6
Cjz928YNTL4H8NhBjVOaxMto1RyVcwg/M7e5H0Ri9GpIjgI95VrmvrnvlDf1kvtCDih7bYCF9Z1M
+/eiPFg4I9+TlYBwZSqnoMmouJJnGzpRIRSSNqDZFnVZ5i535XJK6+VxQ2MMa5f/UYN1TCpwn0LU
la9wp6bXCH9PBErYSiPSVsn4sQBEaPgGUDOhm1Uh2ogW59Fm6N1pC+IiTd7gXg215zH5bArfom2G
AmmOSpMg4xGMcjXoZ3UOlF7FBgIWrGJKBgLdS0IuGsN2BFueaOld2o1+LzwJ+2ZsvOJy1rezmMfh
hbFfFqgP27KWZ4un5l9+5y9zEyRPTlsCIVycutB5ceGGXU/CpfFuat66/QFXRL0b+wXvKHpTYS3n
hni9QRepGIMu55+AXEo5BRglVcIjg0JqBMhQ9qnp083GiEAHWH1Np3EqDCoStvgsdQkgxCTN42TQ
dkwcVT5BUBYPvXWfcqznmortYp9trrq5Kq2SqRdEXG/3eF2HWRAvGR0TSRLg4Lx5YVZfyZgtSyKn
7nRC6IY+Zj2j7ZtAcjV5D2aR7Mr/CsIuYADwY0K4aIz4gQsaZwxenESRUqARdf+VdmZW5GBDLe/p
Qwibi/CDlmBpM8ZxX5ICmOZYZAgYbuXDgO6Ozq9kliLKWXZ40WCGWZhCJm+uNaBgGxaROylXaJIo
WuDiOcEFlIt1OQGeYmxxkqwbBcXQCgm2LQjNDusM34yVISHrkR3Wen5oXftd4hJjlnp4W0ZrYzcV
VcZbYJnKyJ1wWnG+pJXg8IEbs7WeZ5w8KmhREXJ21FzYCwkAv2xxiFLJe1FgfWxvaOBsVr3SGolI
Ivb/265ur/Fflv6Sq1EgZM1wZbJuxg+J6YvmWpyu/+6c+l/J+Eiaz5SoiPWJByZA9NFvb1LV4iS8
OmyxpL2gPbU+dAE8w9oLSxarVsUj74/wDAIdpLWUT0EN+xqZ7xJbmEp3csJgLRnpap5/RwSL7UOW
98DpC2HXlgI81OaMDUaVKkSenzdbrz45flLQ0THHBNnQuPy65sQFNWVbxAYaIjpLKP5q/rVHcpkl
DRSiN1x3AiVoq7ra+jsVxMZWy7ypgxQ181ofQV9onnnKHuaSbujoBfRE59c1btRhZaFaYUaB/jor
lYKdL9P+wr35Wgz9JOmXUZNlJniZ8LRC75iHiOuVWObHB6uvm0L7HVV9VVxh1Qj1/kn8vUPyg1Ci
TPHIYsJZp74ie5WrvC+FSINpchqxieTZRp8d2p2sxqdorAtyZ/W/vmdp7KFiPONfbtSbjvfz9EWw
i1uo9KHePMjPYVrJ4JwTTsBnqg+Z3+WoCZ/DivBw4yHxsHhdPBu9mAS+1D6wVlKqcuNn/uZ1Gag0
7LxMTFRp1S5fXy+nY5DwYtGfXRXlGPw0VTJZivlbveM4JOzl7qUdK11i1QaNqcF1LY0MTtvflEvk
Rqhszm8CvGfdfpCs5lHgNCg4P7u5Tl6/U1DiHm+py1ol1Mbu7GAZWGgPR6d8JPqMD06cNcGrQFE7
l+zV1k5ifKgO+ZXjcoZeIie36DpQRE0vy/gTJc8X3x4Ds1/H3fx8v2mIYD3kJjbmDJKjrAQIWFB7
KYDg4POmkpzWuHMvr1qt1ziD9QOb8Hksrr/JxTO19c9tLceLX0MZn9hfQ8qPSeHNgRY6+meXz1yG
cTakdzyuJyspVquT/rsYeFC043aIhu6nF9Sb+tCwQr/pW2BB9Ua+gY6Zp0zTMqsptS9LoiagWFKM
SO6E/dCGyAWx2GM0/mPudUa0gqQBUNzNdxAxL7echiU4LY5QM/Fl7F+zdNkK799S3qhWxDjMCv8J
rXIkQMBs054n3KYz9pnzjeFyx61ByawTMFSjaq3VAd8GPnamfH+hb59iab+17mTamLfLjdIWwCb/
jP44ijtPOszJw+ZB21ocVYs/BuaiMeTQkmj13YmB/liba8/Zrpuf2iDJroST/3TLYpKdO4ITB2UU
90xclhgw7wEV4TR2nrr+2V0fqk1tkpVOBhVFhilzftgzgjCA447Muz06nN168x3AnALMWFDggYDP
DFSdYy+V/U5wJgOPGaOq2SE/qRFJrWIJkmNpCZBCt8+v3b9AiA6DdMr6k0Ry69jlw3j2KSIKZB6t
PNruA1Ubi7DGGdEEJURgnIOrOKvXLopqATDTvpaXuSOsfs0nwMApsNxi/fJrMkigTIIjiC0Y4jY0
wrbFr9zvDrcG3rtwBWGGtyl0NdGAVYBrblZmvGrHlon28ZZ1zI35nYG7yF/sC/jRoGaBJchOorDa
f1Kasb42/kh5Mgu6gteQimTK7MFH3NNfctJv9Rs84l/d1m22Xnq4pQKya1dPsbHFQdhoR0jiBtfV
a9bahzs2Pvfpts7OLSh1gU/xa+gSSn7F6m+Z3efuC0C3w4s9qIdyZdi/hmPlpT60HZTMm8dImi0c
JaKKwTM5EI5WNGteyMO76VlVgNs1enPlYztjhn5kCsgqjoqJT23a7U5qEu7BmPkmCfQ2WIpeSEsF
sAaiiP7z8uXRBviVzzHOYNvLst8Pka59K0T+VEbshYDnLrcGL2IpO1ElqG3ptZT20HKPllQxgRHy
L6+x9q2+Y6fYvsRTNu16ujyf1wOHlvDz4sfL+m4oIE9qkr61WDHVUY0XJZ8NSLj+wbs5YUGoW6nD
pZ+Jh++EU0/i+9GRyh3PfC48pNYCoJeQwdW2K3PL+l5BlEz52A6pPzVYCFkP/RzmjQ9fm7v4jd1F
NdJhOsPq8svhhWW0O0DAuZea2YkytEeRZGt1x6QjSEOdg1km+gQKHuSJTql34fVZq/K91ESQJ+eP
7RFJeAYr6C5sYEIc+F0pprvLswaP3+Lr0gpN59jmtdy1ORxV4lZ3DTvnxIVIVjOWgsgLK356MMiH
OOWSNtzbh/ZDZdfDeDTSJkQOKg6iP3Mloe3AtnIgaB0I9gTmAaKNYVsMPb+Ou6K7dQj+sGaikoXB
UAJE9E/yFS0PeVgsQMfGOFFiffvXvqf6uiDStEJ0tIfCnRFXSYJ4AN1wlcsGvHdgcMOcUsasG6pp
HArYq7SAe9/QRrsCBP88mPLzk+9PpzhDeMDp0d9xXFuWv1KMCcqvmancUjm84fNWt4hviSPWP8Gg
nIzGz0JsdrxR/8swH6n2q3e0f8sCdGroUplnjTBqISOjdCukXgudKh91E4pIDqL7ETqdiamjQ1wu
PxmUO0OWad8Kb92eE61JV681adLyPfHVlzjO+XDEkWue7hJEjUyyYRqUBE6klLlrqzOTuD8uyvt9
otFvEHh7hPYgWUSK5qhmawQJynWNsEj1sd4tMIQDQBTIbDMZAUT37aAfrUM+rNJLjJHtUxsNiJMM
i5DdHZvJFL+Q49ttXcbT5ido7TB9/hOU4GBEIpsGxHg8+ZFmbT0CbqRhfukfeh6UC9/2L7igrdK1
7gNueycLuDNlUHnMep7K/b6bC9U3mjknj9ykg7q8ZnWZGTErtlUiK98oPjanpwEdkYqVK/vSUBs/
Ega4JdvPwklf/o7zuZAiXt+vObojtMFH1k7VWP4+4fbrpHSonrrGpovdluqs4H0tHZRsWRwY0yMc
HpdgmF6uCgNaXATRDtyWZH5KdkGRBEFLt6vpU1oA0gc0BQiiq6RlrvZSae2KIUzlxRLWCE8o+jeu
pxjUsLXLFGNW7ifQFsQEwwbbRZ/yWyB4W3mPu+pglPgJGKvdlForTbllsUrp54nVMMhu6S/rdShD
ogqyyMbt7S/Xj1udXsfP0CrOSY1kqm3B7V0SNNs1wgkf72p7TgPiE4Jczm/WzTr4Nw901QHyciN1
bAM0PoPxe7vDbBiVyd6A+TgQ33OZ0/Aeaa/DS3ZAVU/35KK40hKjD/kqfkgdAmTcZUGcw5vRADzG
n7Iy43OAXFUmXvZlZASDoG5kB4IpriQoUKrDXmrtMuyDC7ZZqWmKRHTDhoyVCYwYYCoS9jIq7SdN
GJLJhCbznhWT62qTUEu1pFXzZeh0StD5ZbWHMbfI4aBUfO2H6NQuP7ZQF9NbJxX1veuTcH0gef4G
BMhdtR2MxWytzQsF0L5GuXTA1LqNxXHlNM6n7OmZckrZI/jYOhsrRWp7Ciw5fZ2NJVyT1BlOHuZh
chNnIaSGQuL2Ss9/HZOvFWb5kbb3jLn2arEzsjhOeyMIOTaw2j//HipyDekYDHa1LiNJlNh7ht1H
vsQYsqo+CTEVVSHdu1pj0iL+zrw2dciYlXk827N5htNGU0EQZp6xIWZz4BzqMTpjATdSdpc9Fl2V
jo1xrsvRsdFfAZHEMSpCb9erv4nnRTPgs1hPwLAYENw1JfrZ5vjTyrp/SoG+IlbUVXjmYnkKg1E3
tCW0GnBPciScFfX8w43XdqksPVqmIKaiVc2JP6XhEBfOOAWXXWsub2nutNvMOeVrQq6EOEnlrb8Q
4mvZW379jpw9SvMNEvOul/8Wi7cjxGtogT2h8J1JQDInWWLp99cERCbUsybJXGiCHPazzTOZ0eQz
AGiS2S04QkDDIdH2XF84Mtz9K3tC0jdfafrrm1xdjxQ63qyrpKVl0j4+O5Dtig3IMd4UGD6zy99X
alMt89AshYeBbQrZWBFMuKHr647v/iYxZe0sIU0t8mLws4jFg1IOS59O8ospHQhRP4feWMCDWII9
fQz0aw1xV6qSzgqbiM1kGmrI3apBU3iHk8LP4WeQMF6uFi2mFHkXsVls52L61DskT2K2QorYWePr
A8UL7ndjnsmpCrWldJMx1xvGpxgVWqYV+yuw8lCI7/GTDU0JCtrRQHoKsIYWhkq1ucao7Imb3aOw
Trs3VcyP+LBdBTdXTV6DAP/NjEUVYLpLhijdtmIi9CtqImfjNcm+098GLoCtjm/4SPuZ1iiN82CF
rGcIjt8YyTe1PQVvOrk+YJwp+4BuFm6FQDr4oyxYV7JNm2YfagZdAGifOVMa90yac8+bjtI+d4gQ
IHxb5L6eAFcPq2Srs/P/xeJk8HJJi5lGShJkxXdJWd8RKTF4aS452MCUHeaJLCBDAnQzLWi4QUNE
uSdBhiztPcoVin5B68tP8QmFNBwlcmGGvC345tSrhnJ8seEdSVQ7iGNISoa6hhTnEl9f3fbJvM+O
Gzeatir6jJ95M5BCdUntzXIBJ+fFZzzt1Xcd96t2fgS/GLYMuAocHwXqwlTdmq+xgtnrYhRm9vsY
Wq9I219YMBJsCf4X4bArHphN+KWoi1fdu4Zq0a5+Z6VLO4C1tBbsEtr/iBJjgF5mcCBHbhFsQ+vM
9G8MPS/X6CYQwU3HbYew45SL4kyhE+kaqAIIDLTzHhTzVvKOPgV39x1uSugJ9fyZLg1cuCwKSM/B
XsPwkTl2+LKkT9JhowjxLvJKgUvjfiSGO4+TJvx16JMjzBkAY7wF5Ou8Hxl5xFj/QvlRlINBqZeq
4c/oU+fqUGSocgfsDQeCsGjijbvHMY5FBPHYT95eTCSXmy2Qmm5fye6/mkyrpx9EwgCHOv5NOOag
xnDjh9dy0wBPTU6yCFixr99iE5anuq+HIaGvaFWslyJGaN6rMJGdnJ3GAkASu3kgOEBoqrHdczTZ
cNVQIjGRfw47dxemqenZ+qdvC/uSlBsutSST/xUA3Y7tABoePswpoH9rj6eH8/WMKI6A6I2H5yl8
6GNoBZ/avbKaiFlbHQj/t1sg+95rdeU6sK6Hwh8Ecc4ZZDRmVb/ct8NTGOCHMZOpVmxiQCWL53wg
uIUxTCZf35TlmgAGB2mb6MTZGevYn4aYZ6Wu856jUMJ7bsvI+kea+VjnJ2/PystvDPIodm0PW0lO
vyZLWHSNX4VE0ldI2VB+F7r3Kj8+rLdZxcLpMkjUOB5qZtSLpePyV9dX7+Bnk8uuljrloEYdR7BR
RITnTOH31rBRag/HyWjJYoJSH7t+/UOY1/X3KhH67jQKrwxkGQfVhpIBiNUdGDSIDwKdsIzk9Tv+
VsXBMCMpGdaeKKT04SEbRvIFF4C1lZdbt0v4I8ZqrIGzd1DoY0aG/iT8uhVqGU6+59IRgyjakcK7
YpKafo0Kv+XfAh9bJ29Hp8Ck5YOcIeU+qH8iW9XOajhd9bxHgXjprE46ATB0BpFGuMZdrH5zNzaj
e0hAQn3qDuGqMjiIObYm4Y2G2gGel/uML6vH9bhOLohUwyK/4SABNwCCnEVXh21WwRavTkL//Zuv
09iawZmwpYyvqJfmY6ZmIABhsGfCYcoQiYh4AnrFVTP0/+D/Oh364ixXGzBztC+WKcKv74LStyNE
WltJGJ+UdGwDiyqq5cP+IcES4GMeEpXJF3ODr34VFGhTeemwNkAGFbbVWibXDp1brrtLG2iWCo6Q
7YqyO5WX50UjcjUBVZiuxyj9PCT7OUj2TMTnKqtFPeOKLTSkkFJf/KAwSHexo0iIyBdksMzF0Nas
zRHZtPEN0UHu6b+tBajMGB4z/C/pfVoZGi4NgACwxzJ3tya2td037yVE+lBzavUj4ZC0MgON2hui
VMln379tbDuL71BElUjWI4++CQ1RkWc2/Zf86cVXKcWk2+J8HgoyvhdUXr8XcIhuGHNdqohhTUnQ
IaUr+ioLv2SiEOOd1Vux03wafSq0jZglRDu8CEvMO83VuSbqVPji7QRPzHCGc8f1A+YD3J2kqJy6
4FrZSBurtEMQ/k298wpA1lmvsJqN10k2QzHAYkjpg920c3SuEpxK89pXO4uD93rXBN4+7JpvGPze
iDv2Z6/b1GQf7bIwtdzUqNxYm45GWb5EaeyYPH0qmSXHI6saP3um+/WVAISW4yFlaUhBlQnLeUeg
4a9wKhnLsy49JMPP+Ne5NLx2DfTXLPTqwg63dJSUlcKCOOglsFMx78WXpJn+COdzQbZfqNsMnR+f
CvAh4KnC7xx1RhWrt2GkBePZR3/Vbi0a4Xw8+EWue4JsLnRGdT57gbJR96R3QWKh9I2BFMDzujs9
ZkTFdyKOdU5CixErdb7EG7SdXJILDPbdFil1az8jXqYJGL3rRCPrLxgrk2+qzhKqLEQ53VF34uFk
bkURxfZ+s5e8uk9QSxHZREZfjQ7qWhzouK4Q9mvlTUDF+r9AERq1TWpwvtbblq67ST73royRSYyT
dedBEl2FRfGljP5g8wSt1Mra2BUMzZzrGVajQg6XW1/RoVMpsR15qWVEreCvITjYN2Iovkzg42GA
X+U5aEiyTxUhP2Nfwe4Bi7IpLbJeLOkYmWyTLdQW54+1uBsej5XHu7+GY2a0On40X44sGpCYiEhP
tvQs/bG/KnnZC1OChpnal8YLPYimFz58pJ/KTwvVPsblvWFrlM4wWIRn8UelS6Ibmk9MvcIGtCuO
yKzmzpv6vp1uV/mmqeXvc3W3vTU8AYh5AEFx2JKrVHezSH4Dl3u3D1mdw5y5IK/n8phOlReScfuu
pjn+5tx81+5MtHWrUCxnrxDcjwOuiSSJqXsAXBEwRJEFErikqI5Dr93jT3cAQXUM+caQf0qrVPVW
CX9mIU1v4kNaJJ3cufVwZJkyNOAX97l8Rbzb4OOTR9Y0hRuiKbIOejeQZyKimD/WOSfvy5765ytP
mlrjYoLA2/M/t5A1PVQ7whp8cSPLRi/RWpueO3cDNHBz2c+GPuq3BsfWJ1AHRsgMM7bc+OYMxW/t
lBFaHoB/UnJuEr0/3Di/xC1Jt/gsNqzGe/6RN2IEw1wdJ/r8MkfEUJcSbMqGuZkPumZvvThPBzNn
lbWSkn81nnAWcW6Ro2oUjyMWvde/6X3F6PXpheV34JSF5JNmfbgiF+aWq0WNrT6RkqY+kiR94UiO
JHGaycxOpKFYrKPqjXicxU+jkyTx7xdbpl60LL/AzmjtMeWOHfY94OB4IqweVrV9N7YmQCUpfbsU
w9UYaLPC7YyXXig7T/6WFjIcsqzKJyaWpy1i52uIa/W1gL6hX+wS3WSyZCO0BvjoUtAhBjLnV6CK
eqFeHtmcGu1o2lxt/MWZibzVdM8hRW2gZEMKxFfVrHkJOPahc7ywWqpMoWSE7YQXvIrzA5lhA79H
8e340f8xDk00zatGZOqmDhV9PKZFFm6SKuAmI/BqO9h6biPiw2oEpU5gUxSPVdeoof2UNNc+f3x6
vBK+0av7IQHaZSw2poSRYMxzaGqmDPEuDTdBX1HIMs3UbwpVX6rMzTvvk/b++rLRNb8SJTbhSXd7
g8Su9AnwqY59Hn12+WXlnMf4JM9TfGhqrf+1kJfN05tZDdbVEtJPd9C4zzIcWGctQxHYt2kVo9r7
WC8ez16Ldas0c1WE4Z1btKjz0dxcyD3v6l0ni7Y2VWMulcvMeSxS26W0pC7FS+QYlxR5tcC5C+Cb
nNfz32J5qxn9tABtqSALveJs6TijBKOwcvrqXcC9qDcItOEfTHffmF+ELB+ZX5O2/wH5ZCg6fOwI
TaUPtLMlygzDacdj2QrIHZ60qCmDRG27A5hXwTA5mDw2lNRJ0QlFmMZiNf4l9100/bfC/bGPJPEj
3UZ3Ivzqj45EwV423wylKcQxsGso/2dXOGkET2/V4CfJT0+ES4IXR3PfIDJ2gc4B3pPam8oPG2kU
4wIGWqjusSfLDoGYV7LJdf3aBln7GcdtrgaON6KHqAZMlaIwyaqHaDYjuszLeVs7DG6wbyVzEywI
F0lNe9J5vTvzdKPBlAsi5MrayiVoM6vdZ2MtoNbbWY8+3j8o4Q3zC/CmRWPAQtajQbACX1tYzKet
Yz+Qu8dhYfCYULepIW8yKH5aN9awnMyFU/Icy/+S2tG/GE4HN1aKYoIdtkygG/JcKPfbaV3hspi4
SoqTSiq9WGaVgqdfzG7iUHqs3diWorPJV47SbyTDIHKLm56rNBP2f9HznaXpmRyfDe+FMBTBAmrv
GlEu5gNietGQllSbTsMR4OyMcDZcn7HcQZAwEj5y6ORB8Zouy6LTq5QHTjt4JkBy9HVB39nJngU6
9Gsg2vGRYz6iQjiUas67rphOQIPqo+IMGSuXLqdBOKz6Mh7Fp94MQjBxPuzVPv/6sNyBorzLk1PN
iZedsZhJaAcwVjF5ApuVoomUpKgqK1cBody0OsFwAkh9Rx+Zhadljs5Iw508p79qb3nobKZY2az5
CfAV4gzKiC/kKHGKfDOKksB1e/vHtfx0SuWmECKk0MCLwmd1aW5fedG4GeehNsL/NFYmWjDkabHI
Q5XLUDafdDUuvEsb50jUkV86YS277l2l6tvNeT4cp9SaY+GJAtzFtX0LEFj/CcGvCMmDNwZXtWiC
1WKFh0NvtjxWz2m70KexJ+zNh+dJicddj3gvdZOO1lrn7AxC4nQ3Yh6KwDZ3ih4CDEgaXIz/zmAS
f6UZgZ2v2LYmfMUycXqlTQdlLqRxQqq0kiJy8X43VdI142+Ia6+YV4zgDhpqWPjs9s2XqrjHI/cN
N4K3GGNBnqIia46ancXZF9BLIRj39PSxqMnZ4GOhWXdyE0f5eeBhgcm3IeK1rjz7TxDnLINuwBSy
hERff/4pYv/iHze4HFuYEhIRLdwx7EAGfe1KY64uUSoIiTiJ7lW2o+Igrj1DWtRXpO7FHV+k65+O
NI3z3vJuXheM3v8JcC40pJenh6aE+PTuHhDadHKU93f2mS1QmFEkshjZPAM01AbKnSoE4EztSL6P
SGUNXyreDXJFGij1k/i/nEWAqXv7m5rAyYZlpqw9JNjYbqAOOWv4PRQwk3OwVfSOUh80AGjY6sEU
TAQ4jlYS628KGB0w8uG2OrHK6J7YDB18pHkLX+OkYPEnW4jniNUdihQzpe8VM1w4o6TR/lrxGHLS
x1nXb2nX91xxnKtW6IDvPFHldIHtgbWuYhQnX594TvVibcvcaemhfzpuWQFbZe3gMbzjR1lQlV+p
EDqat9FaFrrlxZ/1UfGq/CWlnI54ceLR4g3n4AIK9u0X5vekdZD1PaeAp2TayFtHkXwlR/fEEQTp
EtO2HMCdZhAsWDUTIHvXriP2OBLB07/BZoau6I4/8SN6BeWhjMDrFczbhDeLCrXQwVpmeEr6eHT7
BnPXkaDwQg0PbxaMZndnUztg/iqC7Z3vJ5cyaGTu0b+6k+2YNVFVd7tUPKyZs6SRcCakf86Rw4NZ
okpthmcXESaWDzmMi/bPIHAzI4tJce7JQWLqyLH5qsIecgDn+W+e/BtJq3xHco8+jMIKfDp+kIFN
ws9s6XQ/+NBq25Awk4M7wX77+4dN6/tPiEG/xwGi7QzO6pIp+A6DHa/gfdCA7WgNHnvDExN0Ph6N
eqjWdceZ0Sp7l0MbTPaLHO9RlozRQRF9Bg4GoG8BJjO/JRX1c58V7zbf+KlxJ89+ivWhBGaIXgsy
472I5YokG5+Pm+eNM+/xPUCiOSjkaEXxj2h+Ds04hwj/GHAhm/YGKw4GBXdfiSmECbSrmnAyscke
GaWs6AiVRAXIPEbdu7M9PtS1Vv0JgFm4T5PgEFX9gKq0XoaTRx4UPYgWO+uK6g+csrNGhh12BX9v
jwG2m7KJ/5CGbgiMt+Hcy2GQXm4643aJtwomGkrpa0V3v8OqwqJLFTFAuFYlVpTyOyu/b6boFhzN
e39uMQNp7fdB7s312nMWaQ0nUpiTT8GsQBOVQgGS7xw+sVfn1CRDYIqlp8ePvfmIEGIkZ5yyLlZw
/3lxAbUIZdheE73EBLRIB1UZ8dObrGj5VZC1VH31vOE5RAuzTGQz38/HTeM7OiSQ+UBuICviReV+
zKI+4JPB36tlcnMqvssi1fD8GCY9uSaserMfyJwPHQmI1P3Df7RTz/62LU5g01L2nno0K1w8AW1C
eNEBsaPt8Z5yiAEzc+C7LOzQUyRwfCEKZ1xhtfvI1TtnHffGnmsiEVJ8pmtEdkRgPKbJFx9CB4uP
E6k2qWhMhhOktoTFgro0fjY5L0zCEQbBwYnOKnPV69yPS1+iZDMp21U=
`pragma protect end_protected
