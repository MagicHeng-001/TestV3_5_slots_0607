// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
D81GJJxWhAjqfjGBh5ND4731852aEmYt+9uSlHp9wBdRi3EGjETEaQkPZDruU65Ndg6ySrGzWZ9C
bKlGMai83NCZNyzlZuwARhQxc5iVfzbEfqpp9g6ddPE0C4+nfrrgnTAiZz2NaNZDRf5XsySrtgDF
iYRked44/X39vsgplki+6l8SbvFesQ188z0W9kos34laHDxTWoSwFt5eHc6Y/xyOxI5jO6a4AIM8
i6rkVYFa8dkPeWrfn1TFz+lS2zM9fnKW8gcsetB0dPgSOQEuzyMbXyd/aazH2wmI2kohs6vnKr7v
jyiNsDvpdvAtzVjwAcl/RI5223vxtZHylRGXmg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 103472)
bMX2AByhRLgg4sfpjJVQIh69c60UOZNGi1T4JazlrgIX/TOgHRUgT/j6Y4KjQ0z+wR4NVG94BoKS
n5EvetYQHxQl8JDZsOXpCigPQ5GQz5x0ZVVIizQn7/93X5fPN/+6Kk71zvuISAOlM+GeT5u0griD
GzLYQc7ycXeHCItMVev1TbaVOvXz9ufJYbQ1z+w1ic5GMlXE6ps/lKnts3KVWT9PfjzOMAhzK4q/
RpFu06wL8VdPi18EJyvmrXt5ybNakHCSjqLA7xhcAx3oEohYP0oycOcUx0nUDRRRHks/MixKUues
ABfvULa/OAYGhtF+O6QWQJF6C/ApBzi6BpnJfGQ4YL/PDwVfaFjrv3XmbXGmc9Ko7YJlHpKhWoj6
LQgNo+J1qtMrbAZcb65LIp1lyYFXhH3NnJ8vYjwIYAhHYNhlBvJXFJUzXIw6lxmdhLostKr3EMS2
4sYvvBnVvg1xTntQevv5V1jV+MiSYlldWXXd0nfC6fLlETDuaZtpy5AtUOR42E07n0ETsk/qmuzA
+pBlT2hG2HTLaRNLxpYkJO/6222V3lc88KBr0eV1E5HPjd1wcFc/IlUJZ1ysw7egAgJvn7VfNUSG
N32lMue88yJWCMzxTkjMAqPIEJ+//KeH6wwv5KxHvrbW5PdjsadwBAZwZzF018FvZ9a3iyqR4FKH
evBDw1r1Zk+5RGKObMjKxmFVr1P+BdJMl7HB1Zzc1CGiDgZBEUYc09LDavO1hnhojiCG2f8/5CSL
N4kUJQg08p5jGcyg/lMXJEcxrY6y6tj1sIcyFBa96JWB8wfSOjRC55OHobD81ZWTuC75kbO7YwWJ
e4hKURCjqDSC58REz3plNiiBpID4fYbRGyZHlTJVCInZMq2LswLxgMsyFP+tRSwiM8/0phvX0iu7
wn546Ne3iHYHthZTlvzpa+GaL6U/aTj1rdcQsnNpXvi4umREmBIulvqoCLx42U8cGbZoJDF8nCmv
gXsskj5V03f2yW7TIHu5+ojzhxOQ16HTXgnkz4vxUV0rAiNl8v/v/V+stSIs+fTAnBO2N4f3ygsk
HaVsY3P5jvRmK43l4fvvyMSAnbgMjZtCiFQZjXiEQAN83GR/QDPAPcM5KM2dIAVv2Evn0KWCD/fr
8Z8D8e5FQCeTlmqCF83JoVEH+eFL5xoZVJXK5ApNK/dtXZuSNSFGHW98QcPsmxSyNYkNsGa8m2Ub
pSi3EU+E4RJczEyNNSeq/lOzdO4CryiXO+tpj8+ELLcd+ElBAc5b+cgy4oEyGt4p6rKhLa7lSoOw
7Au+mLSLNftdpmvCHpE8vXd7mMFUEyehmCNiQ1YsqY1fVr5RaW+KE8Q0aeZ2bbdTLjPq8KqWA1ze
SFZCzTIqCslXMrvXGoBOfC3Hu7hKl8n3PHmYd9kHXTzDLZetr84b3bb2c1wibW24ZblInYfKqel+
WmNoMQQCyUP4p+5cO/bQyyuG3ptDpCYeHLnwqFs5qcg+KIp+FYDyE+CzvGmTPdiufTAh6RDHQ7+n
GcrofK3QbtxlHPfW6TYJfQsSFzEjTZToJE9HP7Rg0aSyflfkbwbHSzeXWt4DDDLl71/Jln4hfo4l
ZjTV0ilT5ZQDUDw3D9D8Ee4RknnPNExe7FXa4A139NN3X3PTGAx6M6WsulCSvwkQi3uYt2oz4MD3
4MtaQOYVQk18JeBfSI4rJ7lCiI+iktuTs1CN/JJagpmKwY3krrMFJ7N0Lfh7qbahyuJ3Z+QKmOm9
qD+CK9h+13QTM+Bs397T2KsgpLuDtfBkBI0FmFiRCeUGK2/WkGVc7DagMkgH75C0mKwy2loulAsK
XNdZCpIX+LOjseAD9ksbs52JekvVGMOmeBU+YnBcFncr4/L1febEpnwSrz3zieZviBP/nDmbvJG7
boiDkQt8I4FXBZnRmoQhXXbAiTB82/vmYyruawFOyUMZ3uhUFfoGwntYSwuMZio+GT3v6eZR03lF
VTSwvXuPIh8tsK+P7n6sWkZ5Aa9BzWOsnDQ5Yj3nL2MUJ0oz2QXCHfLGvNxP8rLD36aT/q2EN3CM
x4ZAGetLDZvKyghKcAdkmxm4wzTihnMZ4SIAidqmYUH/JivPcc5wP59owdlrdio2faFansQ810Xk
TINog9QShqitTWo6OzSq226+cGnYwXOUDFi54IFRttJn6warr/Q+KtEsWdnEMWKVxgpAywrpQk9R
yQNnF/hqHu/Ox4R9lIBPdyhM+/FRBN5wAHHiHkqGHwG5eniRAvBhY/FohitO3gcWQ0doWpOwiVui
e0bbdbToWYdtRrzfH2m/e07UML1hZOql4wO2xHIXrk3sIoY+rkh0LhWzU+jF7oJyExWG5arfgg5D
8SzfXISUu3Dz1xVpm5h+RZFqMht8inaZqSgbBd3J4n3Ch28WDW3CA5SqFkCH35V7gi00GmEWd8CB
u9nLDV1GcBB06+g5WSxDqJQ6xCp55u6fOGFvJfMHKLCfnaElxzm3aIlmTSj1tOxTryho2RIhCdbJ
LNmQRXF0FzQmC5zsWZn1ZCsdrqpA2ZIglWXLgfp+5hnvhN695bkH8QKrI51OLcqw1DQesTqroKVi
pqfwcfPssxNSynnDyAUmyUAdfuKZu3u+gR+iMic3l91nLkr0yTsYRIlbD8Dqfm0oL+hu0txr+je+
/R8eLdGf2sDRYMiGgXxGcyIBBgkRWztUE/IsmEkOXKkl78KD2EF054lOI+27SFYK+pvWoXrKiPs/
I5Nrq+ZPI8QVBkZowOzuefUamxCf/vh6pOX6Amjoh9kHa89MdSWr2Yo6a9ZA6ej7EIx49w5S7ysP
I6ILNPUh/ZnjcrKsBQZjcnIksS6NuWz6jdeDl4UMvXTTCKa0MQl0MkEPo3SPWUa3hvZzI7GSY5q3
SnpU3qXMsz7g7fyQUVoFVwyzF0oVIlCiyVwSrsn/Cv37hoRQkhf0arSUGv8K18kQGT+b0FVU7thG
zMYW4/7YVLuAUKK3V+KZ99a7ZNvgq+G99w600bKqikBX1dAE5erlZY1cce5wujzUhEDZImFsbfmc
k2ArkOrtKag7m8yJwIb4UsJ4uXTPEcf6BZ4QYUQpAEuFAX5sJb4JicBE5hnxeqjNegVnFTjFEq1y
SkAfhV5d241DNFht/EkpvWh0aIbykkuwvs6KHlGePnNa3swEHPoEsxxAH2n0MFCIrX2GJ5LWxyt4
aV0GtUOHDF6hVcXVHypwr8j7eKjWJib3nq+fOhHIFGeOpYtFtbjLAImo4LAAmIKSUlFvB6I5ke4W
WnMgWvzzQcJH4AXE0TyehwD8ZTf2cO1OMnxZ52hrJ5Rj7kn1bgDwSRwdm4pOZDtSbY4O1vvoA2Qf
8u/aCbSKUfrkeSroYb30ISI/cNrUpsgmJT/Pc4chW3GIH6SlBFA5WVU7dEiRJRBSZ5ySJvbMQ/+e
qnELwaGjbIvI/ajC7rfsz/QQWuGI/ao8PYBMdN84SH6TOxOQh9vrdlpt1cIx7wZEqeMwDOW65X29
qL07eqI41PtiFwTUoNL+tH9wwBVY9Pa69YXUy84hV0Aho2rX8SlEWClIoXKJA6kadLlx/5l7/X6I
ohc5gqIipdMxA2m+T18okXZNKocCZbFtVjcO+qsVwUYZkE/owLW+1Qp2DBuGh8GJpUKt7lBLUXph
rJJBnk2jgoaNA3UukBPfWUEh6glFQ10Z0+q2XFy/K/NY0zi+W/7AVGs8yOz2Cl44CFQY1ZaerzEa
EOvTcqs0rYAoZWnZRcE1aNX9tT+KwqgvH1/QokCyvKGcUgHCr700V2w0LcVCoVXhTJFKgXsTo+z9
ZIgtocYvZwUeTHkKmQ3N6hnaKezDGfsil9WNGC+OOcrxeTuhXqt3d3wJCUMKIE+fAwNvoqoBDkwT
s32KxmP+wGGvKXq5uU0OxoOLff4gGtzd+//nHmWMJ6GY16MhiNDDKhx8VaQlh8jUXoP//1bwvsly
7TapQcBVcAhoMH3E/L4jpxQbSRbIh0AR560kKu3Nkf3rxTvh1Tpht3YRCCwOJDx3pcJnJqoVkvRQ
HeJhNgecQ4BYvnDVca14gehoVhmecQDGcv8JbLLv1a5507m1dJeo6hzF5bJvG084CSZITxagYeQr
a2756RH3z+VgAwBcHLJSCQp6RhbJD2tFxMym8RXW16cjszQxPMGK/2Tcq/sIRh44E40LKvjmRLT7
jR5MoJkL+qCjxZpuDo+VOsH+Me/NtDLCNx/IdVCTvWyJpP2Rqk+QsNsY1L1gszC7s3fvF96GtjMi
ROz3spVmyX7YTqGYg5xtn5aSLCLx2AG57vYEdH5mUgawVExPN8D0ECSGvfSfAA7iD0TTH4a1cIKT
xTZgKP92P87/m3B5Iq4oJiOWiXPN1aeJ4nsk30wBUiaVAPKpq6qYO1pGJFfC8fP1GhRLp0RAtAce
Hp8rqqmsWJvKjSB9QhwkIA0gGvJ7AaY4dqVU0UXnEjhge0T/cxWfIy920rKz5SDWkXnMWvmb1v7E
GlhK7VujY0VJT6GKOA9lvIOF1PvMA5iMEM6Dlo/c4EUYWhTn8sP77GQcDHNAgRHp2BiRU2/oCO/Z
j41CSp9vmIkTsLkCQCfk7LRDRMBwtMOaInQM+kRDJ1b4UxX5tCMCN7h40E6OwBTKJ4pr+H9TZap8
DkbE/P81c/7gyCOWo6cWtLV/eKBjNVviKFj8AW1R3CvWBEtB883nTcMCyAb9KcnbMD+OTyu4o4mx
71PhhczK0JtLndJQ7kiSLze/NpxISVSs4sWA0Sidkj9ZxCBp926nR2x84a5jAUzpO3FgK1IYU4lm
H/FFuTWdOfKw+xV+sEJOeSj/ikBFB59aZv2miqQRmU855fIP5SMdXrbmL7DJbf6kVtm+2PDd/KUc
YXHS10zpe2h+OBEPkdAl4WXdPX4Vz9EAH1SqYniVSRJngyrEI3uMhExx7PF63uWpMRPeheiE+fUi
xOncmaC7YBGl6HPSxy2tKZ7mF3F9kXrHfl7EgHXqg8btJ/aKpoNwLMq1/+E13s4FIeBtwqB9QUBv
IhfY46eigXtAdXL9hzZVp3tpDmC2RJc6JHXj+QDv9JfrgtfCaCVuAheeOPjlOLxFfmw392GoLZo0
tQDMIIBoV4WOem4Xt3F1yi7fY9Nvwua2smqs1VGAPSEMWnQOH3QPk2YqoXpU6xhPhH0wez53w1Od
lHOluf2r0OFpHkB2C904sLc4vc/WY6pn070InpsIbcKTvXOOtv0QZVywQ0I2JQXFxapK2MkEEXhv
O68GAGVeIsL+Zk9b91wGfSvZA7RHxkwpBRP9pf8cE76IVpZQGz52zLjBq/FYIdr3w3jGl+lKAgPU
GbkFZgITx641LUr2J2S8AotqUQdCRUeoB8FRdoU30aScBXvHua93gfRYlHbHv7ipZEsUuUhaJ+Kg
8NnzZjLjYJy6FwwjEkF1C8DG9hjQKw5z8LWr0pkoLlJYcQyyOMn5q0u33PSdcEFrBjclezFdN7Rp
laNJAZgNf/fphFDCPrHjpNTSfjIQbKZJ4CakVyLjVzZLMYIWnsNllvVz+bRKxEl/mGBFZobxzOsP
gKzUfK+tyihUV8OzKyjlBKGm4GqUh3n26gZm3TVEioXSvnx+odBRITYkvHJZpbaAI00dd7mwWG/Z
wLkEDxRTbsXlwmLXbxCj+q7YmC7P2i3ii2Z98B+FMzOqqqtHKWbvt9m7I6dBsPrk/yOt4hVhv74y
sR+M1uUyNxkk97gfXeE4MG9Ujtq3pVPcLWCm+dDjlQsVMxlsnrzr9UHBmvqhn0RUWLAHyjqLVsFY
gTocNC/VjMDEHGEvnTqfRXsOHobkV+BJluZKArl1S3BDdOSZZDajqqbHShP1BcLG8apc/uI4wjU2
e7LUWv4UQlShnZjfnFPQI7+5ct+zUTHiLI5EKqJ1nT78LXKKxu/+goXob8buBimnV+3gWS/pNMuO
G0AwYsck2S76cOlfab/fXAvWyIVh7GhCpEz7FJGUX6nfEbDbWCc3TDctFGEYXmvjShRKirVnPxes
Hzsi0IJGP5ubODDK5hRlj5HJG7kFmjyBfsP1IXtNiP93V3/Tjqh4coq7wDa7Pu+5IE5R+o32wwys
rqUiOfKJn5HUAydD/eIQhDVfVxRlo3Wty3d0jP3kT7VoptXcLnfj5kHzbTlF388ttAcR3WYcpsw4
vROft6v0vYYYNjnZ28dQSOdwUB4mlqQILpNoyUmzJbSU9KIfgcIh7YJ7jQoOx0cpG7L2w9wpthga
PXoUoQmg0sgMTupPHsHev1C2NYdXCyLYZyOWQlsyokmtMShuFMBTVYVy/od6b1DWjr5GucAGQzyq
cu2rGjrGnUE58dOIpJj6i9vOGdZJ4lhy9CqIjDcTZ0U2WItn0cmh/txoF4E/8uR+03c/2xSHw2rN
qEMm1AlvRwSA1fLvjAHnYD+0k7WpZGftAfce7F54UzsJQFjjXS4R2pX+ub/xjzk72gZyoGPF9ugg
cgq53yGDNN6VEmdFIH8ZN5zIEdvQqpGdT0P28flGGGOuG6dm1wMmSUZ6Fv/G+KCLwE9rcgc+msGZ
/Hfr4yTt6vccSQwazy6qSMvyImXtQJmbDH6almH/H+bTWY4c0+x2O4VcK6+Rj1bCrp74EaTGgJ84
Pf+0AubkYiokNSJNk11ejAD/hFbg1Q3+umabJrMCmSQKYmHsQpVHMU0Wqo37YJiU/vZ3mmozP22Q
wdnpqzwTAvWBKYq4Oe1kKKSw+//401Ia+41C2r4/bW5IRApgXuhLut370x7r1oyI67UhjSx3IHbQ
sAgMlNupMJuE9TmGNOYpHLahMZ1crW7GcO73I9TLwr5Okg63ahaN/mzcVDlpuLEjCm3hNV0B91Cz
yed8gM5LvVMA11stBJ6fXY9ntklDYRFko9nXtJk6Tcu/RjrqttGLrTiwrb+TaGPy5Qk2iwd20tL/
Fxjhxiwklj20VdFenCa+uoIqTtAui+PSfoYU+UeNL77ahEek7IwC+eVG2Ipuy1cegi5Tiw9/karu
DBpNdFYsiD6nLCDREx++Cjqpt0QzNQpjm3n2rf1zZkBgWwgmBTNBHkAtrlTlVZgZVhsputmsvJ5z
qL907ujaq7mzdkNZiJIVa3T3qhtxqFJg7CldKjJOAYWTw9dBnpP/1zSNVHohO+UwoNthM5SQv15Z
kqGtQkTZNFVmv+Aa0ddgyEgRUJ7yXiQvyslEd1oEPo4LPXdSbn9Eqz+wr5JpiVxAbJY3WqClKPC5
ZgnPf8fXLc0+rKSRtfJ43TpDBCZAium0S93gU4tJdNqBqITjIjvTvqO8gbaH5/ywkJWlWY4DZ2XW
bnzuUMX0VEs1x3inTp8BsR6dHpUXQ43GT6P1sRy0WkluQt6EHX8TCFgwr8ufeEt9QjAio0vBDgDl
RpvpWyAUVwCxFZVjYdy8nR8+ciLl4OTyOltkPrNgkexH40UT7uZA7YRpUPNYyH2WLQWnpdb3iQxj
E7juPfNSIgHuKRZ0Dm8LKEUIKbnPUR5SChE8GPz26+7AtozY0sDvHc5D4M+NThsh9jpoqmfj5DLw
CEydkLpbhAUut+n60hMUJMW7YppMuQ2vXqCnSKHKatEaD7CdxfPEtmjW9KuFGUU7ttvmzkmFPmLs
04b1qs7R0XWMnfi+dAmgEsf7jO7MBQfGh8W+js1sA/4fvZ8CjGhPtVdAaJk5buZBW3xYNz5yU7eO
p0t06mkWglEeeyY937j+cEW1jS1wngjGpNcYx7oeUpIj5K3NPgmhIgfO9harN+4M8hGNAaGZCtcJ
1pAt8JM9n1qW0yNhBrMfuQ8LX4zpWex1IUwcBXlMdJaBgO8m9FlPOQTkhiXvDvpA36qvfLQtO4Xg
2hSohYRel9Do4PDlSy54ACRMv8ErJLwqkRoS3kW/3QC4c6tu4zipjifSd/L9rz8p+K20CY3feauS
s6h5phGDcj/NTIPSGIBAnhTVHlHSTaVJKNyCZcfFnDoaQpsqGEUBKN5Ikiik5udxx3U762HEIlb4
gJsBWGAuCDL9zzL0SZou2waguhb04g7Wio0uCG4hhxf6f6HaekNZPWMSCR0Gww8bsoSyFHqhnKam
4iV9ySr18uBcq1qyQodw7QfSf/1Aa7CHgs4W+wKt8aCc1RkdfgVNEZV7h6mFr0TNm1M36q92tnQ4
/plr31oto+GPwBIia45XP8aB+bsZKdQ05cqCSrfSD0tqaw615HeQ9XWOrvxd8vhAmPgK5JIjNE8H
G5qrO6fJIZD3H0sQE3yP4Ac5lKNvMTG/gObGwSQ09MjG3Xn3fYQbk6s0TTg7A+tKYzWQ40oj+ofs
11HvEIZRmtFmNKQ3G85KS5Z/JJy15todC76XzDMe+hDCy8DeBdg7NbfZjjMpQkYJFgxZJk/cdAWO
l2SwANiHswKF/AbcZe6Ug0/SdZi0B6UhU1usnONZuTx2nPg7C9DQkIXLfasbaL+T8YnWfBsp1UKq
F4PsyRHJabCfi9gndybVgIWXxDSRsTVR3OHkAjU6XROHfe+PB3Ew11KsUbtFSAwYtwC/kMbQQR58
fTNWoxuWgSJ7CbvPHGPw2OVFVhWEjx2Atm1b0wTSrAwhMVrB8BLDO8OVS6qaitb6TzNM/zOKHFZg
sYQIir4siBE2vL1YSoMahUWdyDGN0RflCp6W44okSBseioFCkjru3xFHDxyt2HqvZo2c0ZRLGDa3
y6QnAhjwqURi8w3/vdk/Ri1in5yGLvRRlIJSlzf2pr4FQ1fJ4FCZQFrCM3UOoehuSGIqGqqkyuOx
gv1C149Jb0J+Fnv700N8kSWRW7b+rmbbCRaaoKiq3Ke+cRjW4/pFsWlmnF5QftK1oFNOzO4cMOpZ
ZiUhBDcoLGaDAGaZqoH8KjX9zZ22EOkCKCNKS2tTRisU1r83WEfMUfAl5EOo0rVISD1otA1XRm6p
I1ASJDYthpNC/NFahotBkXPdH3WZSXaxi0X6yvIb2ABQy3MndmG3R1qa48QIgoT0V++qdc0gFM+4
O550PRmIsgqpUdIyXkaExRD+CKLyosbS4GTa/z+ZtAU58rfcMkczjJZig/TjS7GIOywvUYI5Udvx
xRvqKsU3RKZ2nmy+53UdqOn1J1F0mZLUHHfVwXunezg+SlcVLH7dvdtZ0VKNATHv7KkmJV44RmCp
vaxNpJKGQA/GY9tVxfCiPq5RSL3HCFfmub4M66wCNlcZVjUlCDt9kyTO1nqK/scbNfNeAIV/r9a6
61w31zsK6N8aTb1oz/gUa73MVWs+vBRok9eSWAc5CV8J0/jqGwfOGbO0VvmgsbYjwPNvkH84EoAO
Nrut83BIrpgYf98ilA998hU/A6B25mNYlzrncadp3hBz7LEwkcKGa4YRwXK3qO5qfRlAgDLp1r7D
LUV0LrvObr8BKnDpYtNkV82OOR2+Mx7tdFsbw4MiNmHo+I4aDiPQ7dunM8VqG4IS38P6hxnGtPIa
JBLezl1eKM34Nkknn1BAVOsC1yZ8DukLzAaYgi6ZjaFb/i6u0FEXmjdRJjedaeDFDfAPINi2pkBV
ERaY3Aj1jEwzFDByk9LpRQY2ijS3yTn0xtClBf+rw28zefcj5/R+vs8jLc2jP8BqaYoeVb+VXnzl
dnv31+t2dCAJUAGykYvv8Uc2QAgpqPSnGb7bGM+dtg3R35lxX0ov7ceDoZHaV88eEcCAZRnEHSFD
3xePjE7Fhbz17RcyWUIadIIAhIgRmp752Bw7ID4WAPCinXziuFnNqAc7mN+e6YzIsIpT+2eZdBkx
/nrkK4lszPFPqGc6G3bf69AYF503IvHZ3a1qV9oXdCwRDaERdBN9dPmiZ6KYsuboc36dxA4Ln+2G
ztXRtYIt7TuHf8+l42jzsJlGfeivCtQuUjax8gtEK5SWbJrvE5RaoVgDeyhLacPzhkKlIsrl7yDB
9I6MCys3b5u6VbUDHA589kaW+OpeieLEbkcMsjLSAv95a74OWysRtyBsJ5VvVh3zRHhc7GF2cImc
HcrrI9oWsJtLlpeellgl3nHkseln9YbeeOEo6fwowFRtz4l8tKAiXYLqGQJ+5vVQ7e1W6IDnF2ik
bmaNNZiT2+VKQ+nG2Z+GIEVXFvDBlui/fhw9mEeUf0Jwc2P7w8hrnTcgSKiv6Oj15x1T1sUUDmCn
CCDkBEuXLJoliiR60SOpq7qTu9UiYYmCBZYGLNmgUVWG+Xbl3XhOJUKbYM5bHHOKgo6OHdiSpVnG
xUZEducnHiWV75KUlmmO9tdcgJ6l4WlnfPmWry4RV5emZkw0kc/FP8O/MRCb/wu153gPw1LacdBu
gJY4HW760M6+gX4IFLfUu4ZisvfrsM5H5zhTkrxnGuPT2yx9jBhgJxUIRWj8ICdvDbXIejZ7+Zl9
/Kcl8ADMH1+gW4Ct5tK5IbIiI/E7SHwAaZ4Zn0Lb8gG7ZHV3usA+vR5DD4QGqzGcOAN0xfwZlA5c
wT7cLotLFbrnWV9a4J5V2nffLn4paDVVmRtoiPSl1iIDBnWcFE488kK7Zoc133Z3zprMbUViSK2I
XVL2lG2Bc2nOCoq3kcEuHVekJM0IUIyz4f+1xe6t/4k4cVrxtkI59KcB79MORjinww/hbBbPlW/l
RziGzWB5M/bsJucc5/zfnSiAzy9QpPZKfwKtCYubYO3ndVKbOayuy4tZqHDzGLzzXjB5p71LRbFq
xF9I4vvO85+OkzrRpM8utG9RthgPLlVnc6TgpI027tnj+gbcHtww2R5KkU0ooouDfXYCbEzO8rrE
YvKtYsYfopFe1GokGDvL0OLwYgGnA8zjicclkddx5HPcWzA2NDahVOp84UfI621oqsYeBoVeo7qh
lBKsvm4n4SV2Lpvwgy3xl6MVfdrhrrWxtw8GLpIDTRSJnL6K9JBwucbrtnLGMCWqFV+NbShbzdrL
ZO9DHj2aWIHMvOIzZ0LcZryhRmVNRiXurqH3MEgti96H8KcfKYdWQzXhh9Z0DR7/J6ItIRLWdzMC
h34Ow1JwGUm7/oXzyBgNvp12NDqLVd9ub6q6t8JaYkBV+y887txpSUIZyUJcTqqgnYPBepJs4Dmb
UD5FE2L7IqRKmb12Df3wrtEMmAo2isPMr7L0D3TlwpuvhUXQuSal/yKVizysUbx+QAWSThz7SYZg
3FRBD/TxUkqjvZJN41myGzI6McKA38Cay8jD9/vdu4tHEhUj/+qQk9VxETEO+98AWCiUqmEyMcOy
i0wa/ujcoNQS+zcuJ5LtV+zTwiFd7mcQG5/Ko40/0+YrHwZJ6ZktjUMejJSmFleiTffz9o0GNHz4
G/YBntQpI/Kfzza3cFQCf6262yewj5O4KHCA5e1xbYfX1ILHOaBiWfpouy58psYIBRJbdniLWqEn
X8rX3P8IISV7rjn9MwfJxPAx2GdjL59OZdm3j/j4IjYwCAmiKpcGGxKCNwX6/CjAq+1tnyBdIi0R
cbxudViTFJXb+YSoZYn54dVYiEv9OFRXDC497hUKoK1chatYAEvhfR/3TeXOxEbvrpDDSG4smaUi
fnA0X9uen7V7QLbQBfNE4lMYtMxoYsoQQEwqYPBba3aE1lkSFrvr+hjYsbt9KP1hQE0NDIOvJV5X
vzczP5tcoY8DesaZifiYXhZzWjaxvc3pvHEZFAAkliFdwN3OKZrw515bkyzDKhcGl1N0e5sDSaik
re66s9kO+rl3xBY/JnQm6zSx1ZKqiVgWH5bBlvmOk8VTCRAN/XvP8UpsHufDxRvbI2GieRW2NEsY
MeGi/mUHRBMfk2od3Hrqqm/Qmi6Ss3fwvlfmLkEM/tehgYMFiQrpLb1GzeE0ofooXCMF5NtmxTEC
55HuPLPhro2vyB/xk4KaIteDxsBof5I2C5R5MI2cnMXu2GhG5LBBv5j6M9GeANTgRR/b8odJ9Xvk
BhiFJR2toDEmwXFQ+T8BnPiC2k8IqFPcQ+bTxF+SbHNddKX4yA/NII9rhhMudLbM+zw/c0EubjFs
/rsW1aqZG2xrZxfAvGL87HQBpI5Tq1ASgfq1fPBscMm9UGlB5lTdANhYpNR6ASBnTBWOGEPuAalX
4wEwMBJrXZU8S4mMbQlUtJSs3bDFFCgrw/UBS6yEG4kQdRdzt2+aYgKgkuvddlhe8bBb2+490/Ue
RD4I4+N4fegwxrtGu1HwWqQqPub0pk0lbJL3255VDnp3FTGau4q0LQXQlQouTDsqGTDAFfljQs5v
SBXXUoV7HitSFCQQAcP/xvf5dGnIfYId3f92ItgxTM0RBnrcONIABboTlahFdewug1ZiZisbT2Kh
U1gyptLi/sMZoxvf7srLkYXw+KCEC/ZXyg9wcKlsiBoSlNbDwBxM2SAP6JporMvcCXlQnBuY8btS
o57OYJ8Cfaw+I4BNpykYvd3uZBYOaGpznIZbBUeWh3QBw2cW1gg0Iz5bkQRvWoiYupxX/3lK1RxZ
+SryDmTNSlMc0LhNGtkQt9Q7A1RuGJDJkf3stFeBz6UBe5NyKtVLTlKVzvutpjSuuPdSy3BkIaDS
7Cy4C86J4B/kvWXIYHWdAWV2xFJw7bptDZPbRqs3wg+/rujbXvALnNPLNfBbbIu9Bb9Txw0smH8x
u2KUqB/azNABXSUCCCM2Y/vHdnCuBydqVAVvNtOHOv9H6L9zUqd49dnj61MtWDQOy5K+F7G8o1TL
xgFWzVcoNY2qc68M7Aj8cksLAY4jY3ay3oSdIiCsxRLenf7fPKQTLDjmmZyKH3rqQscvgM/PJLBr
kEGZ1St3OpGjCgc19GrTXhLOZQIhdjDAKDv1uY8XEo+Yg0xsmDul+OCXFX2OMYKsxK6A8JhPtwK2
lzM9gHeI11RRruTL0Qv5J8nXQeWD6k2salB/gkO5ZLhoh2qr7Bt4efVCWMYUP/YHzpA17+P4sR6U
0QAbVai1Hq3fT23fQwlqDpEzyAbuMIbrWHlYc05GE/JE8hX85k/g38CzvzKSkmIMel7e1KHEDaFI
DG7YjfTpgZv8vRaPgRs5NAGPHHRwiOj9dB9IsT7coBaFRGKJtxCZ14cgd/u2lKq2Kfw2/pRrrDbB
1oB9vdhnRGKd3m+DVQ5ewgaX3J96br9wIy3rDYtU/AsV2hQouaO0Hfxz+vmNDtw5ONDOS6fSdM09
fLFnx8XfCrMQFwYIrd0bNXROAIKw4cWG+XdBrRJ/9DoURzqq6gv4ZofXBjN8tj3j3KI2nkRvaZJu
kjbvSJV2esRAU+8mN5ypJyUnONIDtwF9DRckhze6kzfvOiyEuv2R44m8aGeIf0WWH9tKjcIqhETz
rzkcP3bEoOPv3Eh/nYZJz1hwfM5mpvLR918mJyXMdG6EcVooPSD+MYpi6ReWzdCMu7yib5PPz95A
eEIq96ELpB7Fx6wB8tDAMnasscsWttOPNEcappHGPbhcbiuqTCsu9LZozsQ5E4YgrfZRBtAWYxDw
gRgRo2LLH8gC2I7ZYsbXX5VBR049I3uZbFEyUkni3W0h2mIrMD+3ZcCP7AWSko2Hn0/YBhPmhubp
ttMcbJRunSBctUNofFCxzupJncCoNCyjolrInvBZB3mgEu82aULW/0D0qcbiD+IBateWlsk+Ij3d
0BXhhvgqgMArp588I2UberBB1HjQTCXhhU+xdd4sFZt2/enAEkVxGsod7/zKlvqkg4Rn+jIQ52iT
ZZsip6ckuNBrbeCfk/9lpzZ3xeuiStZwJxPGIi9UvVAhjH0e2hF3L3nwcRUDMe2P86lUe/Ps96F5
7EDRiKCTRjkUUsqNVfYKQt70blc4pl1NBtB0rvAFvnY8phkKjtJN+XpEb65lCsdDPuEw5kE40szl
L1MsKUPznzfcdf/rJCBlxY8/JYOM2EuGfvOSeewaYsE1reSCz+ORw97Oejuf3g2L34vAK8ZVxvWc
vDq4zewRsgeDls+ulKgNoOR4zr2Acs+rkMW0ni563xRM/QExZi4GYCqBru9x8l+ms6EtPF/dNi1X
hm/LLAjTcmWpNpAj7uIWL1h5/ypsuw0pIGNbL05emCYsuokHos9M7DkHH5v+lRepmUuj9yXM/8wy
JbTt6eLzbYaMVzo6ehnkf5OK/f3aChwx+TkhjedIGd2BM4IIi2PzySLGmf/rx02OvQhLUfE99Uf9
C+KJwaSbXNkwr183gt69ruETpLAwxAoxdB4LjTkjiGO684keC13fohm1H0gmgVTriS4qt3Q8iIfx
KGahGiFhxB1JymkYpqNGavs4ioOEkUBHC2Jk/19jHnpx1u84OCHhVIVyX31CoVers7Iolb75FGT7
TYwJLdmUf7Xw3d8PSkSliCR9bjnjgADTmNvktcCXCFYhOW0EI21jDyg+B8wh56A7MNk0pRDOstH5
x3DxXFEdX1qdG7cTNKPCVYXHJGQ2vyKlHhlmKD4EADKnes/BOC6dcJGv7KbyY4rgiP7aBxsMi2O/
gqHP5SVfteEACkaWThBiUkX9NM9Usptokyroxibz1USl95GVmf4mZlpWt1DfcZX3kU9LTfhoPS/9
42ZFYKSEo4co9Dlb/zaM2csfUnmfZqNXf9zO5v0U+MTbeNldX0SS20ey5uuaecpASU9C5+9NE/od
PgNAh8UsrxlQZ+I6EJh72D4sQ8kEfvahiGKyf1tAsIe/t9ctMk+PEsFqYj4i8B3u9XMZeuxIMUP+
AV6V1u+QN1Ujnz25I/yAXrZcTY3kzjBdUZxAv1lg2kO9V2iXdrn2ak370HnhwFgW77c/atIBzRIu
R9IkIbEskLxQ2xJo986Qyso1tFZz3B/UqBsMhdlpTwF4BCrt4Y0Cmo34Gn0bgJD1AIergMiN8mzW
rp0M6jKxvr3/lIgeRmdwZIrsaHSDBXlmjRMAzDxo2epNwj3/6liDAB5oAcUdJrwJ930feqWQJ0Vp
BO6qPA8rPQwrwO8NUvyCLADwmSw3I9cnxmy2Z5SQfRTWmksIasX+G1mj/ZBn3EhrHoYzDXKggqdy
z1TeTVcPythtyODUuy0TV9/yUPWDBrfjlyHbJyJIoB9352TgyCzkslTELRzHqxAurKxJ15p34k5c
n1N0RR0nBIfZYPNYlEkAlGCBJYbe4TJqD/tnR/zyRmOoBx3+ZyNJux6vy/mKJ/YUOP1y5rqfKjrN
qoU96OzksK9oOTKt7vG1KzO7duxLvfXX2hATY3axeJR/PvW1vXPdfTufaz4lA7Hx49FhcKML1wjS
S2e9MB0UHKHx+UgvT4HBx5Igj1Wh571z+qVHVMQJBATfJ8rhHFaNrVR/57Sx3nwrJhgyuzYIzRP2
/bHaWE7R/j1CGS5a8gkh+jHD6jgil+IbMwxBloK3FaIjwdJvsUv75BIlbYUXQP2k9kW8053A9SDb
yoH0q8zxv73InS4SoZQlb/9YkvDF7jRPoJ0Ejz56G0XllAvB2wI/12fnqhGEm2+ucqzziQTiyhVK
kvxZeiijSA97kBcqFScKgQQnPIWd0bdxpatCjlhzbu817JKjGL0Mq6B5Xoj8Yg5+4ix7YsDzEQiG
AGB/Aw2iaDwBoJqK5ydongzgYSnK6Jz/OfkTKqzBmr99Uw1RCzhjvIIorTj4qJD+ctlRndLMNPCX
ZcpRdkmpw7J9e3+XxuPI3QUytUi1ZaEn87DtG3h3nF3b5JMb3ACFXwTmdPYZPb5sQmEzcQBwxEhM
MFxEvDdPWPVSaE+Tky61ehwJjLgoMP5q94/ABcQwaKkSxkwkyE4R8MFSXwL34+P8cGQZeVnpGAD7
KSxdoWCndzGiJ6qwjClatFVNHEZdFPqwY9cSHfpLPo4G0X1fhqhixs2WEJU1aH/knaaf0Zcle8p3
KUEKUlzI1Kd4+BOsyU4oZC5Km72jxPvom6XxzkG9hTjrwGswNSsa0U7xRRQrhchQF5gO1KjxqF88
o7IuMr7J5s2v4fQEuUeJ96TO2JVarneZqsVzqy3sRRfiHBfxZPLRpqW5iCOcKniUYmCJugJk1+qZ
Dtpfro58nUqkF19RkrWdxlp5Cux528ZrmeMNJ8i8sdkvIHXEJ3ysEPvPi1ZA2LjXRXyw1k1k6y9/
/LGC4ZzWc69RwGw4zEuOLs6tS2H1mUP9zAIVWBNB+/fezU7Sjj5Zb5P9zrELyyoWHQ4Ye8AardY5
Fd5OasSC7eGDLLZdp2/wF8BDThWQ1RfQty4dGAwB+JyqhC1aTbUPyFGI7Clv292zMFHWSelGyha+
lt6EjL5eQb2TX0x0EcY4TEaFkWO05vWUEvRMKtpn+FruJKFbH0oWu+dtYYF13u37TaqGNnQQ8WNq
wQBRTjVXqyR+tALKslfSuirVpQlXQFxH8PUZiCjDMGhwtV0DvrAS/0vCGB5Lv2lIGCO3tJiyVl6Y
lozelmgjIvRAnDrXA+dGLf5hXcYmptx8UYf1GCjycLEz7tY9W0HTxdjZRRMvfQQfGSUDZay5Fjay
ddL4lxwRgkww29PJaRj8jrMMrIpKjq5xZRQ4wDVzjYCv/vN1Nw2D2LlZT6EZKV41uC6iUW8C3mV+
BP0BFCe5Cu84VF2tBfoN+SxI19vIircYLZ4ezJ4ckVVOi+WC2FVOf9b6f/pkeLxLhlI95qbUVY5M
poiIDRetHqJAlMawrXFkNCrr3ULYM4FrmlaRBNaEkmx8FEDa13Z3P+HerY7yngdnT5jTmYmzMdxf
KVYTrDizS1j7uNyord5B8ZZNVHsixprylWUXAwnP7hLk28MGHe5FV8gtwClGDk23zrcf3iSb3h5C
+pdjTph+SepYn2MsyB9WWGFjBBb1AaIrw9oicioKMriwAlGTvXu+ADg43xWhotPvunYRoq+l3+nO
eb5Ed+vt/On/X9LWojfq+Y7NeX+dn9rERXoV6f5KDA0ZZh+5GTwRr/ErA2rRbtRJNqSFYtiBsZdW
h4oSbhjYbBNzw9PaGpfegDUryogbTWLSbjnufBmhPIj40N1RwhSTlwjOx1mQhMqPodLnT841CxcB
Q3vzXZWd425t1CM+y34DJjtrqMeBRm0fTJkCpMQbR3bxS9lbq3uTjm4dsk5wz4NKR3hQcIcGnG7M
7BDA3BFOc6DZbKYDG5waenfJVBWrUmqwStnDT/yeIlxFUWjqsZNzexfgDVPgIejRpkXmDDmAyzFs
OgAahiV1dajwMCo4X4g+q7DHetrRLkMVWXvUJKDSe3WvkoaivLlQJwhH8YvPAYZ3bBKOftjSFObo
xgRjiavLvhA81zvfNXThM9sC5rTH/NnmqAUxuXaXd2dh8NWygx8AcnSRCdqHNHXuskMCeAYO9iKo
LIcLlrNlffWlHTkbkqAjQHtqqlKQ/Zjxuao4tkp+605aYwDIqZj+lOtrzWRBGZPY6ZQH9hNHB/g/
FYv6B79E4GTWJE2YziV6wLzJR9jVD2jsN0Uvsxe9OYs6ktcBBwlrqxcORX7kr8BVpoyQhVOXg0MS
AEG2u4LJrKI1iaWWKIlwjo+Z0IxFy5/Mp+IidUOHk3BznPCIQsc0UuGBiQzqVma70VL1g0wlbfVn
dhReASg5DWEqNuzrwe+5ryVu0XjnDmqYProOt8zweNm0MIOb/vq21QdxbNjDo98hEfQ7cFpcp79k
IDAyNmqhL2JmiauO1euK3uK/2rtcnabuSrXcGi08VFrIELNpmcfoHRZocpavw4n2+BNNA/E7kygi
/0fZXOffYPU4aUf+HLXsMKfLIAUyNGp9hAB/SY7z8R8bKiiV6bazNQjLvRlW7O0GpNHnndTbWPh9
yB36BlsnBSVwme14vIBzR4bWRte1c3NbKD2ekpTAgbdtweB04q/osPa0SF2cV4nxZbcEjc0hJ5Lt
wsBrKoj2R7/TogL2P2uZBqvnFM0q/vCqpLRnRIwQxgEI6iGvbbgyHksk5nL+7EaV5J7o0MXYcuCp
aJBTlLt0VZdGX/OcVPkvFyCius1EsVXubCACERhn1Jq4EtG7znIxylmc7DlAhlm9eP3bXsjCkMTO
zzA3d0Gpjvc0583CSbk+qidqgyK+06xh6QxGms3OYqV/yYJk7E4C1lNQAm72UgfqJG5teKjDU6ug
UuRv6OWxxwc0OJS2YniwiDIhzxwJz85qRmf5WfYmTJUjKg2ae1JR2/6cVD+5htBzQVJIo92MifKw
oz2JRLrKz/N8BodUAWp3Gihm+KQEF+FIOFmiQq5EN75+u0WNGKGVhbmDYOJ1mJ6aYBroAZ+RCs6u
pe4Hxe4xbShZYiUUQD0B4k+IbAeGPUTU4P8pPANRv414Nkm6HdClGVXTEE12D1gY4+bit00Jz+Cw
q3snkH74CLALD8fJox4tyHOJyrJjoZiVg7TQKN6QMFpM+cNzL2F9/FdR58reXSLtvvDJjXUukvwP
t0sWgwU1YZ03k4IsB0jEvbA8xcfzBjIMRk2dXzJHs3YcIYhZNuRkZgwu9kD8fJUo0wsIXbD1K89V
F9KjKTFyd6Muumvak7P+IeVyR2rRuL/GJ0kjGtsiryLkL0+B5C3QsMAxUrqJpQRTdt3IeLSa62xy
w8I7yHYJCmRNuVRm4xsPJZ4J59k8N3eobpO3hFcK7giFlydBW/Rb7oLftSlHtHbdaqDy40mJ6+Wl
AOM9MFLaz2cM3k+nawlTODVzHVj9ZcdmMYlg3e2DZ8m4HWKD9rE1cAMKEQg+KXcLHdOIo2aoWQvq
9ue3PzuqX/UGhMo53vLeI8/6kXltsPHeLR1JW00pIkWpdd/YzG9NjEWL1IVaO+Pg+sduGjLHefUW
Uyh4oXmHDuqJ7m5y38ydmqGbBCydUYQlcyBgimBfLY8Nai8im3Vw9fPerEp4JcOHsM9JfbZkYE63
Yr0QXVOvUj9ncBs/degx3KETRm3pAXJK9LrJ8oo/jnyUf+swWn7r07qM8oOZ91vuREU77Uql/3WX
AQzCqZ3V2P+UepT45t4dJfAaRxsjAqGB/DGmhLFhumsY69a3znxj0wgepPXKicYWG2WaaDLPGqyL
UQ/DYrGoLQsVtjqPFzngsSARzWlSlP14PLSEm0zFduZTeqewJU+VFBIcaP8WRRLhWj5D6bM34y1Q
Q21pvaqWBVksPcFFOO9H5055urAlPUcEApBXQ9D/lps2Pn3Nv7FknpcS6uqb32DfwlfAla2jwLcx
VmJWD6mnUyQ+Z8lvxv5Ma/yFmq4Ys0HPX5QNGkwPUXMK/yF4G3bG0fx9JLVvsD/HgbtBGddBxirj
4Za4rMDHFuxktSI4fuoYi5KT2SV6miDYneafXMqZK4RNnG4zUzsk7z6I4oiQkCmH9rrVhmBt3mZJ
s34sJs/dmAlpiuJKvPNnryln/emDQfcKIot/vGzJSALI8uiKCgVjJEibtf3pje5/A4tWcO9F0jeN
mvY/nk1w3zWsdtEUsx3804jZsxk3O8WawSmaMVoAB5SEfvpmrC8yN9h1Z+HW1mLDVNC60E/PvQ3Y
R5KJmcRwg9F+IGhz2nDZEPPUjuWmtiBtnECmvn8BeLrez0+jkI9VagFer9XRkAK4pvAZSCApycGt
IzlJ7n6KP2ejovEOoyWK1F+LeKr13VL/AuoeLZvx/O4KIUGJZwoAvKgIoAKOqy3PGCyOsP+HPs4T
RTeKHk+4K0DZ/2+HqQ592bjb9WN7hj0n1evVc+W9qHZ4GTuk46xZUdDNfrVKghAiy522hfog3ph/
6f002/nZGv5Oj1PZqLCCnt1p1rTaTG78X5bBDPml+6lw5NFW0KKVxHqIN9TerdsofSNJ2pobuK79
5TmxA/+aNSJp914ffiGGuPlloFDglsCcyZkQhcyEklpdYUxvpGhVc9/QsDNtYEODNw/jnWgv/s8B
2WAkYartpYDHNo8Q2t9IprWFkysbkuIWUaWKU7avX7aWrfsD7/AkD6ij6/jAyLtg0iqCWQ2Cse+4
Um6hy/3yssnKTY8cgEYRtqRQOTwYbAgokTOa9C0Dg1XfT7PDroHI7IdeqxBWYR9K05MXSZt8Ht2l
Sd38qUM6LCkcSQktrnheG4Ce68ropJCjlYRulfD+ArYM5qkA4yDKF4R+fAQWDoAFakd3UtsvYlBs
G6DuAQSEtzxdTiedHL/O1lGjDwnRL7WltMp3RdX07xUtOJ/ev6WNF0OxQRy3dLtsXdVdyYAeLV7+
gtewPzOE6fRDUBNxwyWnQfujthsa3alap3ElnYmVy5EysDX+cTlrkUcBIY9UERl5p1zXNzKDGcLJ
eq8/miiAwJO+QZsehkdNVXmln0omO5GAOUtVcRX9JsjurxkzJJwDrXjG+uMtQMw/BGDgfRqI/S6o
QFNoafaCeobnEr7yMiYYtONlIS0UIl2f6D9rYU+mPpWazxDi2lWRzmzyedFXQJYrTEnVVinI1DOL
QUpl+ObInGkvHcLzvHjDbTjjv9YuIumUqGPEpB+pj7tc938g0W3mhYrpLSwiQ1Sqowa+QgQtukKl
gvtvx7XQ9SJwbLghx7W6cwafKYOCc1krTvvYgSY0J429NyjMxwQhuX+c6mQRXmVtOtQMOpQmcWgn
WxBCZ6HIUG41mdexfTxAwqjDZF6jONCBWHhAS9SU+IrudhcDnrYNBsaqCwGkZnK2QD/Kidf5ej4I
qOS8XZ46JVk6RnN3RFbucI+DnsdTDKUN1WNHoRtBm2heCMPVXcmnPtyqCwm1EQ0L+hspQLYNIoTA
VTxarxyNm1o8xbK4C5G4qwnLbGv+jvb/PM4BPzU0jVLhHDyqeqGN2gU0Z/mkg2Ji/HmYIAZg8bzL
tVDvzvVUbwU+nrMV+vjL4kOByYJmsu6BZDcm9ZIbKswXrxzWRSWtCjCFjAOvlt36cOyeR6lA9QuD
x+BFcvoA+5rcFgP/l5wxF4ySxR1jSdPRkXDfsPDCoP5S/QVJZexNtCzhmoTgbZFU3hjMY3jSZ1OY
XCWgJcPdDmzOaFEo9SBa/cuY+mfVM46w/xo1PrWPEiUgw97QMB13EcCWP0PKoNjlrPUGgILx8OI+
ak8f45AkLlyNPJlpLaYOdEBFfj6BoQj0gIQzNS3xdXGqJKaVA+vRYP6fWJJb9b2lFsA7slEARSRX
ZNL859/uwhut6A3qsRNPVyLVjapDnGp054RS+8MhpvId4hIAE6Jb5ZBlck6Nwupc5vsiZ0ApysjT
7XgEAWmEqltXpShSz3XjyDXOTXbsn/hbeBIi6OJ9yPWNZihDU39NNb9UaGwVxp+NRYw+pPArCOWd
LbQn71HBUoRRHAWPg9W5tvTtQ3Q+wCdAZOKMgSaShZmvf7oNwlbymLpye4cmXN5SM86ru1Fgxqyk
UUDqEX5P3PXWUDI4QZY6GF4ongoPI36R56CXatBUp51YlbiQfhR9shEFWlbyVZ6q9+3rv3zkNuhI
aYBClNxNNr+4eIL12yZ0pMgp9Vmt4ceejP/EdtbUb6w+4uFlWaOUDGLnVYreOw79wHDR+hgIyP6v
uvp/9zYYWtkMndBNIP4oI5Lt22hQpbAu4rbaQBiWH/cGP6H0MazJNjMRINn8+DwVAi5Ebw0QAJMe
Qt6FBRSUTo/Z8Tfgds0YT6MHQ+z8mZQCKKFPgmQyNGGY7vSWwgPQs6m9fhyC8oIftnyubSgg3lSz
Zj03gTGBAeVKmsPpUQJier7beDBQ+FbV1UQKV/hrf0hYKf1URiQFj6yGgO+0IbLbEm5UGVWnR3wA
r/r+NWGOj3m1CDNrIXOVYyqJ5Ug8vyJ8rW3HAFi/oexB9JLI5ox4sLDCW4TRuUbMfzg3xF8HVfzZ
PTrIvJe7nguA8tU55foy26NkZbIY2aNrHTLt0pvDzko+52mZi748PIiA0sC+7EHvo0cQYCYeSEAm
XclKMcc9O2I9Pt1mmmZjQoWVCFS2B557gxja3aP/L6Vd927n0xtMzXOTE50XMNBaWkHukMmZBbwS
x7dFXRuQ/NBwdxvhrZp7KitSk9thDpmo2WugUKKJmcb4piiIoh50lLT9RTmOG4TljnugleUQRE01
oLUGf7qKnMue16XssRFrmyEe7A2CLgzee2a57As2PM3ag2Fu+V7hLbwBNTZuOIT6IfyNyKR2QkcH
U1Ppr7xa0fPm4/S2wVT8GCVcbHCdxeNn/GyOjnGEZ7LX7oe9moOIpbZSAn9NSB6SG+nyCZdpJPsj
vNG+pm4N7QjZ2ZB6Q7x1UadvG93yUgly8cH3DDTbSHirNWwT8HgKzgJEmhlFpV7zbHmTKOku0icN
OKw6WYO0DryJXwYaykQ6hzMX08Xzz3kIt9hkWLHUC5WTaSJlJBQLiv5rh4vVB5TAuH75KB+jH32J
JGYarWkcp1pojgoxDouAoecqVLA3RYnchheZm7dd8322PQwTE8ndxE5rroyVnfl7hlQLpYb8dc82
qdsjs/aChom2nU/OA43IIpo70MVkF6W+UM9JsEq0DLA9YJSjtos0Idfk70p1qnCblw7y2VhBr4HK
StOc3CAKf4YmBZEij+0woaopeQwJgyV+25ztBAob+vNC+CuDfi9XMzF6LZv5M4XbYlajnJ09Zaoe
/hlOIZoR/FUgwHek5SSz/CaWKXMrVsMsPRpz9S62zxa8uLGUrDEiaeZuPCtA4DtDSETJmu/THJz2
h2JxU2P0a4lTiCO46CxAd9wi7LkAE+sxXKMvluFNd7jSlysadhpkEjlCSoFnUPZ/2qwMfDYNRGxc
mNehWp8/vsRCIjtSopBgYnPKDwWJnfFNcjBcpVpV5AjcWYqzyaGovWWIqrpyQV4RVpcUiWAbWFxn
yHgGhT5Z/jUWurJanyq+FqPP8pDDVp+CHtJLKP6ND9rTsM7pUyWLClaTwiTjkGTu0VerwBUQzIju
HwrhsNA38m46YrqegTeytGA+5ew4/FlgAQAk+yg94IsI0c2AD6FNT1TRvfsrVZzv1m0uV/9Pb4ap
wA5V/SZiTWFrWj/R+y2H+sGnWS8MiY9yehXCB3z7sLBZpz0zP/56jlBxAaipZYY2oJgJdEVLHgS9
vM/2h4aoUbJHidrC/vfGtHTuQpDdY9aDy++/Ozve1jWudBRb4+N+FwPyCiUFpDlTKPAN9rAew5Sa
HBLRRe695PtqZPgPzpLukO9yoqhdCLOH+NPWiCY4R43vZZeBkLERm04jnpj0CimzxOaGTZFMlDDN
JsMlTelxA9POV+QvdLgVtVgfv5iLGL9poq764SzTNoO83NID4mtRaKxhDv1tH3XneCj9jdtJbs9Y
L/SRbS58W8ioZEo1oJeatmADsFUho5iC3YBtDNQmWShw03JrdWnWv5epMAfK4V0XErq/qEmMTzHa
E48kL6bXB8JT/tVHR72xbKHVqioLb0uD7jBkZU9sxHnKhjhPPc3q6chjIfsJjdBhWJTZFN2oNmJH
eK3o2HPP+DtrEoYl92sHCXvDP+xAQl1eMExDEUC8BBdRKRc+zAUF4mkgVYQ5VT2FNBvrJxl6uW4G
WS5dizk0pBLqY0fmPoesOFDHXgGy6pyiKgEDBGZz0r6JhSv3QsZ06J48IVABTXK5xawYmYneEBV5
rTi94jBWAFULjWY2HEliRmJ10useXWvYboAqoy1s+aXIWDF51vc4USc1Mm9T0UVqUv43QYx29Qyy
j1v+D+QJ1NEl4YUColpXLCsBCVuaHgbPYFL1pSuoao3QTC4YPrmOdbN32vNt920XPZphzteK/kwo
9/M0CcuM9jFm50E7wqNpP8rjDbDaOo4qLPWGehlcsYs7JKK1JVzPHg1F8R2wljKexCWxmlqLdoCI
tX6+oqNrNndf7EWmVeUsiDI7vokUbqZ+MbQwFTRbc4WJykhzsHn/SO6L2WuUFPFTg8TJ6ACl1dro
LB8BWRpQyw+6Bi9mp6i75ctpXiEb8yU8Xp/4BDvq2l96KG88d4QIJjWI1xAQUt/PHzqqojktX3I4
TDSjj0hhXbnB0i/wWiLAXD9x/Kj8x5bpA2rIXn/kMJgc/aCoDNfK3+wB5q3HQK+4uwgr3x8nbopN
p8NSr9hDClUu2EbZtC6O3L06H2BEYakp2EYFclJXVRVUvNlALG2HrhRzsrccPP9EuhoT4ag04Zlg
RHrdn6qHIDdDIuNrQY4aXfJ1oyVm8rfii/eP4EYq9Q8cR0fd78ib46Yv3wZCMUcEOXG8FheQtSfj
zGWCIP7qMleiMzcFAU2yjrgkXuhgz3/O2RT5SEsFYawJ6cR5X3HRt3YBw2EgKpuIzvYmva3ou/7g
rFoG0oBJkL3qONEEhM4cNGV4IFEIgqle2uHPwjoI05zlrEV+mxmsCoge3olZf2oaeuwgK4LwAUUH
Ws1LqUJMCH42CMyaaq6STGFF1OZ0CPocONkEp9IGIuNSsZKG2XTYdJ1vkLt16lICzF586Q17c/l0
ZhiVngAXFuCN4WlRKZdiKFyJDKnHbB+2rzPalQI11AMzGfqZSCoiSyhRuCXKhunhrmJ8x3u+oogU
PiFTXPGB8EYNGKqhf/dVFfYQepDocZ9ZsCva/dlLXWxAfzmQARGEsmvQRhdqEWYUzJD+/OWW6K48
QFh53PTPl0SV9zznhDai5JCJkSpVvKnTdn097kUwuYVPZn2igo3BDAQHeQqxOWnycVxUvyc0a5ky
V7P8vB2gp+GoeIhLOgLmxPkwGMAzH/HGqQ8FIO6+P1PtG9SVjF4HQkDl7jRVFTNEYELoETl1VssE
UyJuE4koKf1ikqRqpZsyP/EdKH4J0IuIktu6MptmcMtXIboh4x6ZYA3COtRqZu0RIwAgsPFYUS7v
Opf00PTBGyGSNB+bUCPrZcZhzSv/ulsv8XPIUie0bTp0PXPFL7xVKehauzi3UkAtTSwwQv/zjeAQ
QJ9yZvT8GexcMJof7QbqfJ6CRtKSeNyQ0X9TMH335igIpl6kwMhgR89LrHeClS9vjb9VqfHwaLUG
a6+tqA0Bci/0lfxmWqlgpKxX1PU4RYTYzALzJPcz7sqN+vc81PP1HBOrcwrrD6bOOpRPilG+kE8D
1UOE6SE7oe1LoOpjnXglPXCSZKzJWvMVMgFP5H01W5bTeIljfTY8LOAGWz2VlvJxmE2M8Q4T9H5G
G4AIQsi7cV9I5j4q0n0MxsR5qb9czy0iLkgDPNsYJ9mlFblGpT4PwqDrYbgZtyAoccjY9B0W0MSq
stbT5hhpfMnyC2kcU0eOHm/S5Sz0XfdUUeBWILHH+Y+fUR1uKmV/EjEK7GSCNc4c3rVQCaKs7zg9
31PC25OJCqof7d4LTUhQiJn0Oe9m88eBT1gHbyAIEOWctsIlI66xTAiEWZgODNh4C4aQFpxHCise
tHa2DkU9/YUSfsbVQh2X67KQyOiuCqGF0RLnMYFFtyNu21Y7Vn52BZ516WVtvZs+mk5LTX8nx6ju
XyUCa+xgLiYAGXBQ/SX9qZ700fCkp3Gn8sP0uKluQHe71BoZX6fdtvOGHgH4raQ3Rp2yG4YXkymX
IIRtb+ZKAdz8TACe9N7DwE0KNijUwXO1eiGUroXGCeEKqqtPFvNejL+qhcJM0xLTY0/X2IwsEcPN
DY9XNtLl+qZih9U9p8caRqIXWHCbvA6qH5MtGLaYX9ovR8E53wjz0a8tJ+RZ8eLojEaqCumkLP/G
F38BPYq1hXrzkcF5s/48/lAVbgdhsq6hVu1Qy99OhEBQIrkqBHa7WKgos7H8ZwAOW5EtTcDKN+e0
ToNewLbzJ+yD+PRZ4H1FbRdNc26fKOoXsyV4N3xdoJ7VRAyAEk6v2aw79kBQ4wAylFEVD7Pq98nZ
+PhE6/8TMQvmKqNEMRaeAcfv7uTh4w8rAWEfw+mVgC6sayKjqc/WhpV8Ufj0StM/GRM6y8JZ4cTR
k7rOaeB4e0Pv9p29MNJaB7AORECLLhH/VaRDiyZmXOQb95l+E9dAt0F/G2wr47T/P0iSViA1R4h2
CbZzWt+QY/3tOhnysxqu0QUUDr+UlG6+HeIxj9NMTdyhYlWFvTMa4GQJ5Kx1e88vZdwWlaFFQrYe
9SGLXrCgVcDXkFi2A8d3xu+VZFXxv4XxsIdlThCT28V0utnaWEgewELVoQR8arwPsmCrl39i8/17
N2eTn5/thiHx4PTAvy+XifshZIZh7hsr9vaiIecKvgiDhDdgWUOSM9VHUkeiL+c7DY2VHZ5MI1ba
Y8CJjw5Q2KumS9AMlGN0WphXZ37qf3ntgyBUbyd3GfPuEf24gNVbRdM7Fuk2sPlmwvLjyVB7WnOs
N4dlga2HIGpMbm/ZHYyWXOrclhcALsvVn+vgenoFssY0vbHzo+6fBlsWxwapB9RYyxtoGXz1dRg+
hVikGBHz+rUKQxmvaIk2kE626QqxUszy64ryrBI5d2sPNLJUXq14fu7PLH/QRR60ccm82NSV0SLW
flTrtSvWpiUrJ0smgHeV8G4W4saE06wS1TUhwDsFDdRy2TuVEokfEU58NfUZ0BfDYwZSLbQ9mQw0
LgHdf3/H6HLCe4Y86Ia+mudAvX4OnyOoPMncqDVkPIiPb94CcbOrAkXMCxOxv5lJ7sHK0BTlLq5K
XC3AlH7RDFWsEIHM9oYylPdr3O5Z1DsiPEemqE1tMYShItMeC6NRxgd2gtIWzw5xFUjPBmmPgIVM
35r+FWfA6GdkQV/yn6WfRsbPuHLhTHaqyEmlua53aJ+NQYY/ovefXN3NoF9RKfM0n5pKywYqJjIM
DdDZZ0gjgxL4VAH9mxsMoXKht1mSGqn8GYoHN5A6qHOxao3/+D5K1KhG88g3/avFxJ/7mPASe2Aq
5coSMGcUEivp0cjT78mjLcu/MvFRYrydWeHo8/wXWWJ0QBr5SS5WeYLVUdxrEpYmqsVR8ctRpPny
HoriMdge/qFHfgas1BBzXyeMiLnynrV1tnukBVEmDY8ekD5/eelIKw2b/G+mOAT1zJaB3FEm8//p
fiM/u/mSEcdTz9uk/kJJRuUz/O6/KI8yNc6D0s6C4/uK3IIKR123TL0UmbctZQe2NRMb3ySuIwWb
qGm3n0wN/fnOJrZec68mgxu/jJ593UuCx2Ex3a7LwhslKhkxro7trqq6eMhL7T+T02u1z8Wla5L1
QP3ECxcKODkwvWrPg90QSube3XpbJCjso7fNXJxSJHd41vogtV3oAE74HzmG7okz6Wl9rmWzRozd
y5q5QDYDNERUWYovMjbF0cjjdNFnWJ0mhIFfOagCGwVA8snYkzjFJ9sNMP4xKH7fiAoSzZNVgGoa
S+uT4/R4NUjEl6w+5vkfjcVleMYAAxCWJHwh76uKZ0ir5eAJ7nsXEHQ4OI1udQAuVh6zsRb113aI
33eLiDWI5gWLBCTNjYfjFRdzvwAkkzOHfodAb83xGgAHngfiE9FWQtvwfGwr9SCoj2DGtNsOc3TU
zod8NRerQdN1XqCBcCmuW0t9shzAAwdXI8+NPSgKahIbNqKghY0TOo1lRp1L5CN+fKYIWyvurwsj
Va06JzR9ImXqZ+E4jmC19TeW13aBRzQGnE4ibwx2HiQ9Qu5PWglNBNsDbPIECP86LJBt1NkjBvZm
bJRvil4cdsJSOmudoyPTQX5bHzNMVPk0s01OTGpukGQvAWhJu7d1NX/RkTmQKIJwqS3tPwno8dm7
8hSeNdin0hTGVAYjx4BPk3Zi7Ri5gm/naPLkQfWdvizPEWV43QEK7EjBpmeQEPxUD3gvwq2/03db
fzIIZbn7/Ei2x3JK/1IgcLJqG9o2uk+nN9n7AUMGgV6YxTQ939iPfZAO1TJR5qTrfudVYKDhc6Bj
i3FaD6NPtstKbnMnDiZcQ5uK0snn6gUJelQSTl8MFPt9xAdwdY5XApD79OUKSISWIVrtNwUyiIBc
KHF4NyvtzzE4enDb1kj+mp5tmLFmU8KNDp2PNbYLzvTXOKm6QanuLkqw+2t5Pv1+cGvHRBC4cwOs
cNM3yj8JtsqjNo+x5hKlxesBFpAWhDeXY3L78ntZoeX1vGi9MWx4lntSGWP0VyLCIork6Psy0uTq
6qhkLkE9/TEoM9xz8S69jxTXuJaZ2+bbqsUC2EImgmxTcPNhrjB/gyOdm8iS44szhV9CHTkoXMDs
TXEQ2KQ0NcLEypMJRPyrSP2GNigwYGvDgyRroROzH2mmmK2td7XOWPlpwDJL22NJFglAFZ4Zv1GM
O+SubvPbxvf/2FgBX8ZpnitcBzgzg1weJ5HWgV5OFozBTKhX/TlKdf4KtJReBfSXJhq9NHd5uc1p
5glrIKyFKjtsaLqYNETEEiBuuo8IGPELKA22/38m5w5kCa3PqdLas2gv397p4+3pZBmae4U/VNQ7
OJSu4FyuA3LGlleJREpjzpA5KJsOfPzDMgvXwFQaz+0dJ1YcH+puO3J95+aJa11I1yCSMZ3aJjqf
VAnkxiZZmCZXwoNU+V0F2HikuXyIhovN7O96QCq32clojDJWLMgn74CjtOdctcZCa5SNVMlfA3M7
yFwyTmNybF2ylQeUY8LZ3sey45azu3DYUp3WlSq3tFhvkLF8963x2F7tlzliSvHKW0G7A+VodLi+
smHo+vkadS2fYwuU+EYSVLk+zYa2OCRVEUMKwy8JsobOiZAoeA6dshM7J51NI8c7XI8hno8V6Fjp
eXpUm6D7JzD+KyhDL8CcFahKmAy0x8ydCMT5ZlqQtQfwz7rI+eqowvcXqTh+Oe02IfqF8LE7+103
L05isUg1mNeWmGd6ZKmVwHmqrSRYVLEYl8RTOya8t9bU/RHyXc8QiZaitaWT311XeCjmWZZE1lDX
NPSa2A6yYYuhJQaITPXLMB7vhIs3pF6KfDGJkQ3yVxBNnl0cxIgJgMMEFu4GU7KI2L8m07n8x7EN
s+UadwcM8xCzEGMBqQOLmOpb1dNuDTfxSl5AKfkAvNCEwXVE6PXu/9LnBjHkbi90j0EWVDD8sdtN
01O64VTTqjT7ewbXefNWVACSchTiGPMNmhU3wCOBOHMEmH9sSsLFXHq6uyEZoWWF4fiUJfnw+yAC
RCzlOfNp82XiIWqbDaqVM9l2AzCk9d5RFt+kHYanDEaRFh45pBZ7kAzSYjfVnfc0SqcLxd/iUrJE
qnyr1oEGSXtRiDd9R4MoVo7I2mbNnE9TRbcdZICr0eRU6agSgKUU4v0APti14gWP/RiU84oPpiQ8
0Yebiarx5dyxNnVJ8nCRD0Ncpc3CbKQHPC789DFskurNKAe1sxTEmc6mk3ufGfWqPoZqpVa+Dmjq
nAgwhrZirhzQZRB3VApV9IGFs8Z3qJO938cCDOgAs1dz5CWN7aDLdWRcTxIVoLFN00ohhpJ2HXdd
jfL11JAhXgg2nrymZAEUkSppDy5BTiC9iQJIvBPxpXuya5hAVr++bc3NghawzUoHJCcw7Y4C6jiC
WQ4J+fkvL7+gjdtOhD4hdfeTcyJLgc0LL2xeLBU+5mb9icggPoorqVU5l9m5R6byy6mSbzxxrn5T
KB1VROvKUUMq53ExFb1LnWpos4aI1ui2bE9B+TmoHeRA20SxgtK9lxgILaYkbmwd0QJA0FAw771v
Him8zTemBDb3FsXvAKF35hRYpVg9NKXmLxYTGbL1iNwYj1kWB7+Bka7i5J21N6xkeOwtefF0V1t3
308VXdY3T9D1ZXBwpuyZVlkFBmlMUen9ZMPAbbgGycQPkA4JaVzQTXQDiz1JVzAcgAnZdnol11Wb
dNl5nowTzs/wHdJ+sjJZmtjWpIJW9OtRQFaRWPYKfffc7NYW3dDuR3ZY5+a/yh/TwEFT92iSv3L9
kuuAwGN++0+8zaWfAO8mWnv16te/p3kbmbAeiRLMI+4d5TIURjgcMV3LZDTod0znneB9FWVwbdmy
ZPtD5D9az18+Zp/5lXbH8gjW+2EBtRW84Ov/yb6WEDCkz+rEkPb23e9AkEsU6T5V25erMb6YfF0P
UuNsyZY2UaJgYfvLs4aNYQrZYK1/1dySoXCwV2tyl2RKp3sryzOLqL/Sw4mAU3Q7GpZ9ufk2Twui
FNHnDYX1vW/6KTahufw9MOCyuGmBdS0zjGYhfuoDWkIhnx3GGI74wfuP3Al0aTYTrNrWJ8xG0y2a
SXqCR5W+dIiHr0JVFBouhCa0hDw3SrpwClJgCtOVeV3sIZ7Qr2hs6lZxV/uomxiehHwGEJ3ywje7
900YMdXkEyDKOuy4JLMZprRuHsIvezZ9oyeA4cR/QsZNYx/p7XSWHpTgfyahFND5eLVDywsRccNo
Pyocpsv2EFSD1ek6zYImydjmPEJi5xT/5BdXdol0vgpQDdlcgC2FYbXOMU1C0P8BdXok1Y4VWHuv
zUYoqP2CYOmr748xk252ohaCn9m50Y94ykcQGQcthek+skns4cY66nR8EiFkd0PE9+oeW47xwA73
sniIhFDphp2KvJ98R6S14aGcOUUedOztSk4xrTkbDMd+M3toz6lIXoBcPyk/xNF/gg3UzKKkUwD6
HhqAh1ppr+8/x21WcLi7UDicQRp5c6gWooYHid1A0ImFXxkP3ZvTdMUikbqM3JDceblGuw4SZR1w
JGwcaFE+5GpX/iqvVZPw5PK2TL2F/f54srJ9Jr8YtCJJj5jJSIy4Q8SYlRWd8l7fErUUzVzNnxeC
Vb0VN7r8rEPwINnl6sDICCU7O8p5Tw/dxIuW/BOS8DfXn+V7Gi/SpvfAeY6VKudN9a8D8i3j/bjH
FBR9ZuktMf3glOTb3O/+97wdwZ4NIsrQtdtmCu3slOZu004T16xC6SsRzYynx+J7difeTfInV4JW
C15mJgdjCbVoZdaob5Fhx54SnpxEqk6g41bE6Y8mRBV5te6E/+9x2tzYFq3anmX1lqKymBLKOdMR
p/qniAuJeQspEzxiSGZIAcM5jNoCc8/oG7TH2DQu4fsiL6wwLoUa8FFhSJyOSygn/27AHvfGb2Qg
b6z6GviLhNZ9yBcoHqa5pgWUzL1n1FipRlhwt1M8hCNZj6v9n3Ogy5gybQd4g+UetOqqRYMbID37
v5kGnylCTUT8y2c3PQ/WspFtzKU5oYEqqiWmqrEgeXomnbp6w2Q7QJ3LpcY71uaZsPCYFgqE7GB7
2alELEqLP5g9xnAA3c6w3OYvGzJAT/pwcSKrrl/4DWYmV0R6QRS+EHw2sOoaIcdiAFAENg708gjM
fq/lSdRZM/zySBqEpxesr4ETxlaJA6eCmVgtFgzo8RowVUaok+X9GyUurmHtEXVQv77ruMO+9lRW
Y6HgIbdHwYsd29xRsVHgHfHncrcx6QSr8KHJ5cOXNDjBDoUWVaXvqvEIDZckUKJK7I9Co4BxxzrR
N9pzDkJrl2+1M6NpCL4HtYViecnyHY2exhczPaFq0pLhYyDi5pEHESwa3nOTnZKYa+N+zMWVo38r
PBW0ZYMMELoNbVXnsRFYu6v7gH++BWeizTAtjYO7E4cm/voeM6FUWuW7Zm6mC1wSJAZLjUj9ujhU
W2ooKGIWTFxusCkAZf1f8xJ5xUtwRF9+iyoTNgJYPvWV9I8qVB+oS3S/CqLSc0zEPaacAOJBEFpn
po14/lKz5wBDYDuP6Z5bzCPFfDF9NQOOXUC/fLpVTAYt3HktgfDuCUbubRguChXpanegyTxdr4Fu
3ZnegdowUE2HOdZOWqKfeGmYPrJYtqtehvVG4hle5miDi2qIpyj2aCMo5m3xhNKeljlKCa3vwqiH
B9SWvaWyUTBGGVY/J4lWs+aoHgvnQCCio8z4FHoCA3Ti4QHMfKPtVoMSRUArx6t4jIEG2RCLlmtT
/G1JDF9Rmx2BSoDhrov+G4fRVGDoKV/Wqcnr60ASklTMuDTPG8DSv+Buun5dWLu7Kwxke11X/k5W
8igmcoFWMMm5YPaPlsCMaE1L5IFaE8QefYO1fVST0z5MqriTfQsBfYNABUUNdEjEjFMgR2R/FQaj
QisVlkM9LZA/LwJ7HR+B/EgYxABYaQuZw5b3UlcWTR2EatcbTw2vcfh1Y5w+XOFN/MdF2YXn1/Aw
7+0lWZ0prUFUPy+XclI2gW6MbAvjlW9JG4hBFcD8fVlIti63hCAW8v8guEzcA9LmL2cE5IowjspA
/QBBxNckveNDv022GiY/tXGTGtsnb35zUjU91ZiW29JIvY6GiAeS1VzUTwUMwrm8yi0g4uZexRaC
33RoTyzUJUPBpGnKCxfdqLvnDiBVf4EFDJ9AfgnYJksKJVlCcpBctXyR/mj/yeUxdxpofDjjroqQ
RzGl7pLjll/csdMSlJa5JsXa1npVqBXEfqrcPvz7RXsvpj8dHZoMbyoGoyz2v6PneBnNPTFytKXQ
UBcOiVt4cLOZ5KXbr6HC0NgGOo06sZtVy+iZMQhSnYXlWp/8GCDHUYS8Xzhnh/j2BM7Xb5/RL6al
+a+UQD6yweMgsECAehzeKU2uKlPgAxAUZI2WflYx9PHKJqSwB8joN9WtyPBPeP6x0GT369S+E9Y/
ZlLRtXHr8IxWoUlphfc0Vz+B/ySt4wiXMaltXF1ja7fA16mEbR4cP5hyoqZPq5P+9RPvzslB8UwH
HV4h0k06Kwr+Ksb/hb+aKxQ78L3wukp8i7yWu1zwiwwRXJXnF9XTrlonWyP/m8FXw9GKLyV2J88p
ZhSoNCiJ0ycAZ1Wum43ttsHf7dqtWdgH4Mcy0Xiho+dLdcpS5An+gJL0w7xPW2kfQNX0XySDsrL9
omgPXhr3iiq4UqmfrsFI9Uu+uYkxuJqWRmtz8tZohj4V840Rhi5E8bZvnfGjojPRtGsB32K7Dykt
0vOXBigcboVQFljEx/cZn+5uumDBA5uimDpjh7V8hK6sLNhvVCFju1dp+bzDEtEppjK6gLSo/8Sz
SABupB/h/YqJKXX9P89TFWkXPNCIVKPdjBPjJKNsoLBQDJITHwWcArVmUTok4eHc4JhEMaXHFlcP
iFF4wLdPsxeE13G23BZzbCk2e77X+zgiqizBZR5yoyIsOYT8aI2EpO1mpwIhstQgU/8iclvKWAqn
Nm2ElxL7fmJY9Tn6/1h5EeJsNz9VUjrEbA5t5EN6EnotxrOole0Ok0zVSg10FKahyk3C6z3CMe6t
970skIV3Ouagoqgeec7sD5/0UtkRV6H+GLdpP7+fEv5st2eix4hGIwhfHkpV3QBbYP1r4lsBmpt7
JtWkuX8SpgHkJIOxRfq3jlz92YK5MvbGoxHMzSh4PWAi7T3Obm7rW+MVaZpMFlr/dGAxb+JAXw0H
00lixoo8j1GYQF2ugAHJuPwmd+FMNJYcMYRihjUkdDNgtPkL+TSe+UMLbd2wFuwPABqV0hwfQ/C4
Dyi4GZuhUStRXassflgYdhkE/DERW7lvfJUkHj5//gcNc3bycW46KFt9feMHstxXNXwWZekFF3r0
FkekCS5GwkP1CTjwHLoy1IxSB3W+V2ZvC8z5Y5zGqd0VkGvnTBYlglpjJgKJJWY764FTgM3U2N63
HipBRvIilUvB/cNku+Da3SfbhYnEgt5+Kb0IMbkW1yMpoEizAfYJWGocHlewGN3FevWrktTrOzMB
uDXw4joVP7eS/TCReGXmOJyNn0TaFNV5iOHRgIbXgD3PLmtFlTAmlbx50KQ1BoMxSfMDJ8lkYeCR
98T2wqWvyVuJ5/VqHOGKyS4QC3YQE8QU5CK5EX8SN1Hx1VQJtLkebQHboOACjZAfDN/ABe8zreC5
ow6MFxVtSuBH8TeyQc2C9ccBKz8QH/4U1xsv/1t6LIa+G9Ltpf3eLEh7hhSYpHeDHewMAKuzEvGK
TfpNudrJFMpDpBuQozEcwBmtv8j7EcR/LBN4kGdtPdR+Ytup47lNb7XNgiIv6ayA0L1Ki3YnsG9F
lWQQfZYTeCUt/vyd8dEDosuslhK3u4dBD8NL5V+d3bdMCCn/nRNu/8COyFt13q+1Ql2/JVj2bH0Y
YsPQin0ddKBSoz3/zTnzvuCtBacSQLJY/7DfoWqGGBt0b2xXbBK259+654lu8+UFkFbbLFI85Cyv
4l8hBMwZvfa/YmcChcTcgu01vc4RQVdhdux7I3v9VBfSkmnpl4vZWfgXDuGRB+YAsHgSLPJtJoHE
ylPApyv6JLSQalvSZC/zfcyYYg5kv+UkQqkjufmF90eTtBfl7Uoj76sdPKJ86vMtz0l1vQqnV69+
oG7LaZ1lDcNpo8Qw7zSq6sNIe7u5ukWmikw5tpXK7lfboMwCkdr6Ojy31lI2geS3QNWFtlYKBEnu
3/ONFxCgo64fplHLv6Myhu2Efv5/G3gxpBw3zaGNC/CZ52zZ1WxeE+z9JPm51R05gf75fKnw5v7v
/UfvQht4M8J/wEQrn3IOVfdmZa1BfQYaCDwIhbh55baK8E+3IZxKly4Y5oopL3uSPikZmEMNHbfB
SToD8YErsaS2Go9eDvBfjN2vb5IMBp6m+K/Cmr3kJaBv6z3eAnqyA7aJum5We1P+xH5hPpb/UMk7
ZxbC/BYVrEw5+EE9LR5eddRy5yeazwcDprIm/p6bq1UfBMhWa8AA8JyOfHLVZPHC+X5dPt2X2so2
Pr1Adk7+J0Icy2FUvDU4y80aBgsJ5rPM2/JMl4yM6CX3mdhanZyMg76E16ymN9Yy9fnORUQnS/si
vjaQRdWHrVPfr2qSt0sv7pF3t3ZXrSVH0ajvv/0a+3IuvGQ+SRItRpttWi23ZKEHAdY5sd/x8rht
5ZCL5HBkHSlai1PrTmRXs7v8v2a+EqRUujzKRn+fNUxZVGjHgIyxvn4lPcR0FMA516RJ68CQQUCW
LzSrMgTHXvitDH4LYADF9GIDjwZjL31g7QMJk8OS2xSOEQn/Y7oBOi/3gUi2AFc6ZnLLR2A2X5lf
uFcakRSUEDFQdy/NEaHrbJNOvpjydPIaudWDPcqqYAWlaQDaaB3a4YQsCbWgv886Z4iyvpOn+hPX
YVZbVq2ka/T2dMMGCfyEOelWsFPLLuIP43WwzXXYPmmD2z64MZcn2nNL38tDzZwb0RIgFYtd01NA
6SFmUgJMkGGL5ptEUfiKmpTcz3FEfe/kHIUeJlYHb73mSFzPX0VH64NsvuxcqKSvTNXedP13n/cH
w2SVOPw3HJSpNTqia/APtDPwjhmaaMadks6GOHs6DsquOSD3NJjXhv7NMnh7yeBM6RIKh0j+hlmL
gxhlLcVL8A4OsEF8g7XKLSSP4M4ImDg8ICG37ry7J1MzM5IT95QpvYqatABiWVMTWULiXoKWxlOC
YtYR8ozTcbJSlMh1WkhA9Wnw3qI668j9JJn1yGj2cW0WRWAlHkHaH9z/uGXMAs4qKaaT8+QLMRIp
6VvQs1+saNYl9PwGan7dDrHK0a1s13iYYA6WyiP+PnDySvfCUXqVWXBayEcQnFPfAiynXRiVXi4A
nddV5EkEhciiIUKBQGOHtu4n7VYtvyI4F9lv2rS0kKyKevOdh4vYlFMgQm3K8xl8dJfa9tA/8O3B
pAJMvRpOcQgRRxl3M/MHkjqzd5t1HU7z1vk9pER57PenhLXutSrEtH0Y8eV7PS3Q4eb+Rqbr60ff
z9VYZn+ytO9Y/6uy/2WVyD7KKwi4sfTAzyA25LcXeGrbYt94kfP0d7v1skzQ0/7PXIEzqqaOuFGC
37/ialKXAL+fLnmFFDW7g4mItZWz8nbyYG0JdKoJVUFHwTEJopmWxwhP9mKpfZVDUCAn4ipfsfr+
khcOUm5ojtVFykGe9Epe/1ZutPUM9VBktZeUlFPOcOQ55CIHgTEveVoIXmHjQVHvhRH66nTHG9N7
VNyPAtvjc7lvy8HCRkEghow1eGcS8wAwdJ+dRtKS1anCSwMlhoyDwZOEMLLrfBrH6zMmdUZAGz8i
Hr3RrlcWXh5NjDnBnKEAM7oUXFuXtwUCke5ItLOrDcmytVMvOtHoI6Rlh2LvvRzyo/MbVbCE4mHP
egB95T3t7RMLSsNrFaSLcYhi25+6QKwIGy1DqHHylqzQ+JvGvgAg4G+KFM9RskaRaYK2gIQ000Qe
Aj4MqMuhoFe3Ldgjy/GzkrhPZ6AWs0RSLDjtioJR1GS42KJCKhEHb1/G+Y7zyH35eNIaBjcgBCDL
yx2lHJlAFGytxDJwMvhw7R2TOLPTk9IBWylH8J7hvYifC8hcp5FxjU74gCI2vWVW3f8xxd7ZxWGU
hI244uScyceaU1DAnLxdYhoS4aoRuguYmuylCQWYOsAaRxg1Y/n8oX3KvilvSkoVnfIwcQ4tdprn
62GHbDwfkH7QlhXSBdNoFnos+0CsaNKRpZiSFASMoek49H5w/OJk79JS3anlungX9uTrNDgTQY+d
kzYbveZI/C/KIbtdoI+7FYZNGEBJRWDAuUIJ8B2KS5anPToUrfuaUlJaLWeRIiQ5mRL2NdPD2Xxp
kVcx1sIjB8a+RyTWkgAexGhxgwZoD4Z9jxB3affQU0JCA/KdUL9EohtcGH5If1qVXK96bU9rs6zY
Sj+55GScdhJLFKFwwQrBxLDHSF0R3fbFX0t9ZZZ5iZLNClY6mHwfshCwqyaeN26c8+XeUWSr9baV
Syxi3K+Fo54uW4yuGvBCCZJ62oeTb4GOmlS30lFTkRdAEO0I1R1kUPn7Drwr/FaWIodWo5eFb19G
vqnQi3aPHUfkN2AVBOp6et0Z57sRKcEh7NoUcZsqA4kU66qn9mN50iQLwKPB2XefhXPz4WUqoQ3p
858LIohRdpMaA9bL0X3yZEyhG/4pbIXHMcdmGuc+P1QcY6j6JL9yDqSCv2H/0tc4EByqkmF9fltt
HOgC4EyJuXvANIuRTv3HT4/RtmdNNwhnUZwuLpK/P13G2Ec4IZniRjGY7q7z0L9FMlMekg8XY27w
Tv/V3+sEHDgAjaYtWMRTY2ymdSekjT6hrDRa+0EUmari6Hj3mrQO+PRLOJ/8s3RLdJY6+i21+O+R
GT2ooxZ1ivbd9eqWP8KfIZ+38p2dBfRjWem7STMfx1+HVva6PfGRyzzLdAGHCnFmJkl/sigS/h3k
2tth3/AInxTpKNGXIA9GzbX4SojZ8c7kWKWCvOw06WHy+pAiOCQs3dN/fryA2xHP+QEiIKhoFrHl
SXF3Op0nrLtGCfnVQdeO2v0iNN858Ru/wsVxVlP0qtbTQaD2mQsiJ1bUMqcy/XzNhWAdSf1A+fv3
Y5MbhCqJf5gvzrE3ZXa99lEx4JEwLEZffCTvFtUpHS47rioElIcuDT4Fg9ZHrGvYUL/xxyZhQUxh
RU5YwCl+af0MWIO54Zjh88X/0EoFK/dijaNMtkaU0j2dEVjxgudvFYtFDNv+z40sum7GA2BuJNA4
dZCooRDvyH/sotw0R/kzOS1H5pVMmHhiENPWW0PNeN1zy4FAxIS3On1sp2uUpb0Bywss6KGIFKRc
Cuklk2Gt0U9opduJmrlh55DYYSsV/tS74M7+C+BAnpa5nsKV4TXPeAcya/xnUdexYvBwaBB25ko4
1lXgAS6HyIxfjh2Y1Lw6FyRxOBvrgW9dpNT8Q1Oyaqq3Zdp46+mSIFyjvkXoa0DbwLItnPaP4eKk
7isugekVhT4IPvN8Fo/Kvv+X1VadSMr52bZsII7YHQEvwSZHynIdkB21RhAv7BnM0aCd8Or57sU3
3VjHSnIENZ0dt6uANQfENbCYynZLtNgdmqQJGdOrTSyC8pLcDOh3PPp9rP3dJMN1y6FOxSuIt5No
lpN8C5yFiMyFqdzrOrO744ah1Bj85BO66C69QDIRw62zCm+P3kbMKVh30Zmcsz8g/3gJm+mgzuhe
qw5yy22fQPDdcUgdm0XUGHc0/md/n2bZot8l5+vvQL7orMRsl0XaUo54wXAQfVyT+f8gtEA2bzQV
paEa+JbsV/z4kFKY2/t9vCgA0QqDB9hLNFt4XMvfHm75oPsVFaoY3svPGFuMOaE82j1jdn+IAxNv
k+HlZhJKT1t1rXfSp2cS7f/zcZfh1d2QzLJcxrR3FkYeLebRxvUcROLgJALTfSOFswBalBhdHrgU
jZ8G9fYRyylBGV7FqS1WbK4VoEBvsn8oCXkTHo5UEYzqMJwhLM9JBTNGrOcUl+tEbmj23WF57hfb
GTrEFHW/1vT0keKeb2qQv1mrIcL55afi4OE4pq2l1ExY5uP5ddP8CKJ+OecYX4PFH9mDdCxNFnkP
CVjbhg4GEe23GVh+VvGPNdUuG+dVvP81kk5QD2bQR/fR/1DItbtBRklZwxqrKdgJC9RqgFLYwCZz
rK21RJiRNDnR8h1WVmo7B7IVgwmTqmHVqFr5xYNy4zOw0XvhDejQCSJxXE7U8gu1tT8eDzFmxmaJ
h8KFakoUh1nWz0VMPOFgUAxamTDEdKzPbjhfXbrkvLsUsAMbybdWQE1jTqYzyjPX/glYwoukXRs4
n8Ssd/+B1eX3X8O/wQD52PrY4x5uG7McjBdEdDEPcWdVWeui8F2eDdqKjW1BMkju36+j9j32a5a7
GO7O3UQjysrSv1MlZrSeTrnbl9f7nyrKQB6Lz0VPnQfwch/KHkIdKVd+mANyl8D/NAiNPPqqwuOq
Mt3TVH85yvrLIIj1MYkA1hGKusGye48zLQ1FV2jRtWx2SQ5Q9oIk1dmneFRYjgEJCMG8ndlgA+/m
4VWOCJOUcGfyYciOpPf78u3/N8JFSBIkYXFg0o3euNbDtHWy+HoseYbTa10z/D+E7CR8wWQkA5A2
9e+Ev/GXTh0uqTwoqHYVENzevrpyzU17mbw6VOtt47Z616298GnCvUCvUP95CsIEOGEOASGWTqkU
kPULEh00hxHPnARms77QEPO7WVGG6GPz9YQHiuU0IUYrouRYnXzEgLuA/8MED4zdqm9qICOEc0Jz
dqPNnmYV6ms/G4XuwU0d2gspdm8ToJg5tB1ZEDUxSgBnwGcvhHveJv8uRXaX1IQHVdDMT05R0pMd
pGdasVCX1jfUbrzFfvMBibZ7P+mPl7+/MB2C1sx/wSmOWUpNRir+tcuul7Ap9VyPuqnO+KnnOobm
YCQ0BSF4+b6hEy2bLuSOtNGWCgZw8GVs+CuNZuEMkoKi33v3EZZa4yGJ0zpVYs6qS/W7vQJYgrwB
VLdHA0kzn9NG9x6in8/ctr2CX8R3shCy9CmcL8boJPw4mrhic78FTKdXqs9zDONFam5dyfEqZevt
1qelXMJoI8Kat9vnzl8czen8sGg9Wryds2fgbBOKyG41piTq2W+FvNZbpO2JYAS27cEAuIQBXkI6
WGcoyIRe3ydN+u3NMI08bG2RYqQMyyrpVezAVTqIvF9ulnEvPww3rI/JpDvPlplNgG3FMqBTVvG+
JSEX5CwQTxYIMcvV9vlqLpgW6KOKlGV+wiMvKY/DUKM1ELW93gUriJiuJWXDMJ+cLRlpYKTjcsdV
bJWlPZN+h+JES/XAmN7mXJEIHq5hDOLt5+bMo+VwCabCOLOZxnXeYqv4r8wz6rrc8d8mGgImID2b
X1nALWA+yAcHYjY5oynHNUF9CqoEQAuEVy2A3BsmnyGG4oGb9wx6u8uvHdOw/PfDvFaOIgZicenF
0VxxWr8/WR79ZL1LHUDCrLmrPgt7aw5Z8ZImFItq3u8AtvnMEs5ALKg9en72u5wUP5vzUyje/2OF
wZ+M9luwaUez3sjZt46IyXlqhHLDVE3BJhvHRsiS6NpqAPv6pc4nzJ3XVROC+n/+X21SMiLWKzkW
YVtnLJ+mnBuaTFyG/dyPyvrrdsuDk1CnHp2s4QEH5x7OXtLKc+mh0xDmrlPrwfiGF3k7ybcINmn6
SH7CPz4e8YOE4lCF+OAr6xB8Z5hLD1uoGFyhD0Y3ChXgZ48iVEWOKVk7LzXxjzmUgP/YQJAGsHAC
C9zmwklSf2OfUcayb/O0eKXvIAqvk0n5kxrEEG4G8rdnf3xDeLw12HMmi2+NP6n6gVCuaDmScLWv
4imFtxg07G2/tQuwzWOGxvOKSORLeu1WXhpTzvj6UAhuSTdTDjdQqVQjtoMfkLkmPRo5HjTO5fMt
Sx17XDhBD/7zaAobAgsXSVwmXtdMkCBlQFd0uYfhBW3ZOm2Lc5pktDz7X4c55jUCyWOLw2qFK66d
bXpSJ1N9AnneVLnF52tFf1BU8twfmnmMzhHkABzcTe7CXI1c8vcKH0Xcbm+rkBtC06jx+ZAppJr+
7wFWcguJiBT5lO4gFjol+f4zCxns0oBvLtRcxJqnbK8rLky/Mrs5oIAH2e83n90z7yqdCjTRqpcl
B2HdxhOgCdNA5ecgT6ubW2jDxHfHzjVOAN9jjK8LdgU+subuD0WTSq5xJK42aRBB/vilzDTQy4iu
baar3i65hihdL0l3wdof96gbpT1p5BYh6GfKDSl0pC8auM44bjzGcWpNcsKJVBgE1bfvhkpPp9/z
4RfKhly8eG6xHeLtshtgxejiLz0tGPlsrBI1OxqDRbTgI6e2M2amFqgU577p333oxoRt5gd6U4ig
kSsGZJ9XCLQBjtPTB3l4cCNoO9XuOF0PKckZnRMe09HQ9gMUaFp8tKsFfLOuqjjFHzQehri0xdFc
U/8eq4XdSZqVJCJ+wiZkGLb0sHf1bpDXHOvQA+Jr2MuvB6cLcAlWka/MruvQPWv7MnbHE/1vUWCO
lvHwhQzGo2HazE5Vurk8pFxxOOUDFjfJ7Nbey/7WOGbqmgpfDUJSKs7veJ/+++Z1EMuFPDzuukT6
21mbsCRrPSczbH1TxOtHxOdqW0EtHWPqkOF/EZzi2yHQoDfD2ijaT3IaE5BEGc9ak0udANe6tzNO
I6IDC7vhC4pxOYrUtahtutWTxMQ5meoZreLYUv0zFewuDoH+nFiSe/FO/663Ln0Rk03v3TyRbB/L
oFAucYAtqvGR4c4XNkep90qAphEMZ7JiEqKh1sUQzV8+tFCUQefmqMWgLVT6h+1hr8gd2y42905y
eriX7slM0Bxagxb0jxSgCV/+E8qtncoVebd191tgL5S4afV/YKIBdJ4DqHXbpDpw3yhC0b0FVCwJ
NX1rIIEmZqcPlMZecmZqtkvrc8Us+aVBCUWcnUV8SY6tP15pRDamAfH5+5P5UP46HmXzNd/f+K1W
vzUN8l+Q7IdXh31lkYUjWB2gBIKVnp7VnsENQzaAR1NC9o2P0V/KeLuAhtAbRFBuhP4b0d1IzmqO
nlAYFB3aMj1AfnHW16sn+UBJiR+yts0JUto2OkZLJafEbGZILqNV2xEqIfE/o+R66EK0fMAJOQJW
V2ZzLgsEaGCckwtKzP5DIGFBfUDCt5U6wRjLOLb8FUjE8is6ScPUcYlAegK43X4BlD3imkxueZ3i
mw3TBdiVvHFII4lsllIiXrpx8RaQu8FV6DPbDAPHiQpuforRBGZjwz0nonfT7vEafMriT/LLhKCI
okqFc7A6TA6Gp+HxaZT8aiHGobYSBA879iDqD2v8X9ZTjWj71AEabaHzBLzi9uwNnVYQ2EIaX75f
2VRtuJM7oSSC/l84/mOnZ11xEkhMRp8biAOcZwxlmrhruJj/zNosQZlHLUAzyPJHk7l75H10Xd35
Jz7FQ66bR0C/YvjNIBFSP03h6Siib73wuXsWCriUNj7no3nTbMO10wFXgt+vpil4J7BS2TBBxYXq
pMafO7JZVD4Fv7CcSu5cSKUcBj1k1eSNj5LRUBA/s7QAsYHQZPG9b0noUSLgTxRqnX9VfCQT1DEu
1A3FDJi+NNUl0VXiUPW+yncwzMIV/ow701t2BjLgc0yAjG7wangyITNiFdJrfpiKaApAu45SZ1Ag
h4c0XGJ904dDHxX1+1u5O6UuS1RIzJozgfZpU3n4Xv/c9hDMjVrtXQXNWNTgGAevpFcbnjO9CTef
zvsy98vAneaVEP+vpw9wZ528eORWKgfYW2rbWpu6cydnSonb9BuWBEt0PzG15n1C/uEh6INl4pDX
tsQWKWcfxoo+KQAxV4/HdJB3J3PiW5lFsPXOJUYil26zB/YLKSGN9wgkbRnrBJ/hrhyyFGqchWfB
VXB9qtyA8RWVEraWpEFH5jjoUvPtKuhtNuAwl6C2WDJbvlX2SgyyXkZqetPyIzN528GqPKcvI3ML
ps5obuV5n7qb+knLeIUi3/ASqszFeWAdNanh7deLG0w0L+AHzy8Rl9YbDcGvBEXpQPyiH2SNxIIV
ZCsAaAf5ttsXktdh/fAyFgW0WuZOKGgguxNoKIULsE8z8GXUDMq4Rxj2Eoysdg5P3Y4VkJ9AvYBW
+5Zep/gUWqryZkrImNwvGrQlTck6cMmJWMmfbqjHMARGtNw1nfae/UVw663Fqo7fBvSo4z/yLGxr
bW2MqTDrx/Kpuj0UkChraoRxJ+fyJyqtTLU4bLokQQ+rrEwDU3bEsy93Vo2FGok//VBC2L7tkQYd
7AzwP13d+7ZKIfleOZPtC7RAImpYkuVprsd41nv2kfJsMMJ3MB8oIaZyO3OxSqzqcHKy0dhQ/nIF
ZlvkFrCrIFWo6gA5Dq4VWAuxjlnqfOpGnGf35iRj83JagEYreaOf6t0rYb+QwPH9KCwmukscYsas
sjoxiKpOAIqNAX+E3NJfTEdcej5Kk6fGEKWfDEPcFL3xgImSAXtvvJA+t/iEaEBjGmM6bySA9pTw
pi1f0YTIrS5IYDYtdqrvKZZTcFMqWrilJv2DcTbrX+CGPT9+B1R7UT1uROWu+/C7PBcktwqplgZm
0LJgOjLyyroV3+mcubJxaN9J/UrnUczU1hRfIb+XeOjo7nYC2esvMFKI7zXkAd0pemc9FPls2JKc
HMwtsB8+lPCHh2onvpHytCYaz3apWEoYmJkHZQ319EXQhWt3EeM3mp6aE1FMG/kID47lwGJ+LFwB
s63lbKcWGgVmd29OJLUiSkVy+xxdxhiQRwtuwkN7dRcijq5lE1U6gTiGz27SG/Dwy5A3QV+i+o8X
gj3PBEpDWdCChmKWhjGh8pMLKFnLwf20Z23G6j0BP/LkxI8oVTYJDsfuWujVwuAw7U1IVa9LI35v
C4DWdDuRmo7tQ3cCIBVWDMTJkD6ASTgIuHLOIn3Y0VLhn4tXogbCW+BcW55JP2xMHTkKUbXZdSQU
w4d0RShXMYoZknQg5OJr4NJWEI8hE0FHfVEtLlUd5xgUKviwXYhV5RGNgZKbHeg9jvO05pyJmFf8
5gYP1HWuoASUEGccQAu8OX/VWeE4+hb/iEpQHuQKzkWMzV1YtYDOK6av1Ob6YYm9L6i62cuVp+Dp
VLWq1FE1ZuMuu89f1WJSHP+OSnp9/thku6o7w3Co19B4snomTB/hEVtPKc31JaWzE1ys2ijDlgRe
anBrlCcvvcZOsQCJZp7AcxcEbxM5otVrnI9mf1aDPgwW9uDMaF/xVc3n8mtrDhgZyKlxaiaLrrwE
eg7QrXNhuYDKp9DfquhL3J2Vcyoj7jO+x3Q83/e1VlvvO3zpG8/7faEf+i9M2M88ZaWzr+lOMmwZ
Sqs5VOs5pqWWfweClQVgDfb55tegZMzf8WNK9eD8/vSmb3hPTexcd+D7NjnHkG2A4vQuFx6dN8i6
4xisE0ZFVKk7rMDy+u6DRMVbut5spUbM+uyzV7Z0wtZ8X4YhyJnvLAL+Mvx8TN9ROqOUWW8BPt/I
yFELZPrCa52Ie+gLtQkN2Hr9PZ1YpzQIl1u7fDKOpjZObcenbsqo1nfeX8UgABdsnEO1avJl1tNM
X2uh1sga6powpFpGW8LCUeh7kgR8+PD3ivV3ZXP/EcGUfvesbxhZhaxKc1jmS7olNOkh15cZmAAg
hCHbO6g6xAYiQZUqDbbglFg9KojpOXcCYLivW6e0fiTMqekMEO2WILsJtpd5880Lb6bsmKUeJ9vl
5Mp73s+PgHCRvGcfiEfyNnDeSE7Qc3VbscYog7gAmiDd5PfrPpPkOoU3ggbuOFard+pcMuhCBKPN
IYOvvgmuYzo6DJyycJk63ueGZRy7CYTruemaVALzawx/FnzT7Ioxqj/llDVZKlREmu8am5tW7D1g
OmjRh55v8eWM9BLn7ssgA8MnGtJUuj9peiHh5mtHvsRQOEHgdhUZrUFBn2LZKHUfPIpRAtjzm+uz
xQe7SVkXPH1GWZ5dVzQUeOP+Nn4jVcOn8Cc3Kr038kJfXIhuNvAIjkb2g2Ujys1VESyFaF0gJHPP
LG8vbqXE5N1RI05zE5MrKE08C7VKzFW/vPgIhPLfP7JhMYPMpMnGQ7gOGSNGN3Maxn5OwC8A4I+r
R+rnU40bRJhqKoO1+ftxj0eNfhkVGdG4+lJBnbVnVaUy9wmi5dWkcDiVXO0uLpi0QIUpW1ZTBXUq
WBdiNgM5m+8rI8KcfTi4PNbEiiLBCPOMumAozvjKX7hbMZo1ICIklnRRymlG6Uohn9Rinsov0+Sc
3+KKe26RA8NLjlrVvp3RdS15khPYPotsdMBJy7YINPNLRR3YeTiJxzKoho91Z9DdNnRsr0DnQz1L
Tu7A7kGaSO3T1AbU5BM2zZUUN6u03Y4DZrmYw25W0nrA6R37/nojuqdCVrt0+c/DB+X1tdt2LWQk
KDdpKATVSC2DVWRJFcOCcsGvDXwEBlIMF+i6BXGSEpexJCCS77DQTtSWoh0EOkQWoawJLK3deNdb
1v2rZXssidp+maoga54+GnIo9utCEG4pEKjb7VAisa9Yl3iRBnEMSMuDffDaz756G1Jhz2mKv34P
LNh9WIy/YbKhUgyZgbV0Djjxsdlacgkyyqeld6jbYuiND6NiiBJwzCmQYs/iKhx/Di8SpWwTVTx9
aq05pVDKT+9s4cu1g50YhYlJ0OgJ93bB5e2ZvSyNVQitiOXWqjvl+392aNBjgjVaDZ+koH/6G6QP
A4jRiaCkwIJMi8VGO2xxyApu/yxIjixK1KMtaE0+vdJOPE9ON4afq5KVzOT8JQrOmSgFZyYtPJTQ
ftWaMtRlsKmWsfhccaJ0I2SlCfO0FePGvOUqvfJfO4/qcc0Z8S3OFdfhXNDN+vxLzHTnogHrdQL3
V813QptT+4otTNM5JINw/gauxvA1YBDcwuc79TlCLGPMMt2jkyeXjGQVHl/tE4NEhIPFG84rtTVA
UI8iKjSqTswNPUaEhVo7HjHR3TuUcTXRli82cbJ4DUgdrklx7Vi5Oh8LSoe+A0ehvdZieYXFpH0U
Qm+y/P3gZLA0/2MJaZfQ/+czQh/tfpANrcYEYcjuzaFCCFNof8n0fH+czDTMGMPadvHDwV0LW2RV
2Iz5qBYeVWifbqXTVlbVMkcAOn2UwrYfHi+c/XBflkfxxQJTN4sPC8n9bCLrUPJbuZsXi3g7c+UY
FgXuYJckIvXolyxS+Foay92zemy2//3uvxnmG0NhHeWQlFziXervGm4eo0bGx089fBE80RLluMYa
Z40mek/1M0EjvKSMcsyB1yBq7MGjs6YIieX3D5q7m7x8Fpnzebzp6LrPkU58mypZwgzvXOL0illY
HdDafHmahBUDyzmSJDe5wVcMXD6A1rlWFkC/X3v+t1Azw+3vMNTLCwlfa22PTHYeDlZ8OQfk/EfA
I8Xn0iO18B+4e1yrvgFbm1qdTQKOHnuFGiY2B2aRCef3H3TVZdTNZK/19yJPYOpm51NgjUfeJp4P
NMd5aMl9KP5de2XHMszqUvSIVTXHZSeQMthSQF1I/JeDaRj815HDvesflks0UM+V6F1G5XQ9grO7
cjT1bd3ItPfIAeyNLhHh3uiCnAtQHlFC5ykacNChqKH1tO71jLOACf3vU3qA6KDZOJMXqu9LlXw+
muMTE9RyXSsTD0HMzx7aTbwEIcJCkDcXuTH8WgvBBt6mvnhJuCtdP/gE8m8DALTdl2YpOQ/3YKxf
5bEbkUBGvv7foWNFSFYihc/F28tX3qfzKGyUNlmlPZvS28cFaHDy+ACdygc2L4yBo1htPwS8b+A3
NMK7Kp2RhwIV9e24+7YCh7mkUxhb+nSAED9WAc08i4wOSjEuViZsCTL7KwWn+quLmI1swGVHPcOF
xIpuDyiT9g2VBqM9zToBHaBq95Mm3wRwbxdiDI81JgJuBmNs90fI/Ek57k99/DB2FdifhPbJsqUY
xWRGSjqxwBFkO7TAQJ8vtLb9EIRZ1V4+xY1Q/WD8lQqVe56hprKP8W7Pv8Z5Dm0xYDczQMHTQxz8
peOP944ghcClHn8USrdG8+GD/cLVgqwoHq5IozNbdVWYrSfFAgxz8oVXNfgHXDEneg3GHHA4G1bv
Id0fqiL1+mpMDf6nbvzh9oSmFTCNPSyDGZJi+KOMKUJFo/ChZBfEgSVazy7hRJYGuhUeZmE6uDvS
8MiI4zuT+w1XkXod365Rh3prSsUJcSGGcbnlPAu1wmbYj/F4MQrGalk/BRpBsLMS2xHbnhgAH8La
oolhtqLgCXIOMvbIC8AFoO8aVvACac2VysemRu/fo3OyryByUy1/OtN8TWxu1YmOCfN7lLMUwbks
ISSdxBung5M8Cq2cF4TB51+4CPEf3ZJikpc9HHkIbuXsGCaQ5Ya/xpjv2V+Twy87Rfp/0f+r56L7
UUURbw8LVCOrmzF079s6CS3CJ92XJdmCUs6dkZd4A86ZoJs1yhTMmzcNr3Sm/89OEjPp9RR7sWy3
tYb7k8n3eQk3JtRGt0ni8djrWhQyeEg5bowDvVX9uQyzOcKDJ+AdZXqRtZlF++Ux6pmY4riqRJAl
MpY2dZmws7cSjbwmlMqMofwn2OhvvLBmoTU5LsdvtU1rz/KO9NAFQYXjS5KRtDJOX3dO14hV4jyK
ombNALyYcRaYUp8rVLHZXzHFlDOixZSM6mx2hZjvQZW66N9f0iluQfmOHB13TRcYet2pOmTdvb6j
QBmypaXQdKT07lL+XpunJdFvS4Xub+sjl4tERJZY9PZDZeYFw2mohOMn866wYywpZ8aSRLuKqO2s
J4JzuQ72NDp4qEs8/l3ia6NGnmIrq6CCWfND4SMeErzLP0DE+9zxKxuJuop8tQaG6WIkdmHQaj9w
dRSQRwQgJ4Cv9xnrQN9jleSjBUxKsW9ZQrxfxvkW3WROtncN+3+87keJVJtBNsQ0tvOWglN1VrmF
PJ4VHUgiu5G8i+M86fzM7Ihk4KxoYYkQq3xq7SGVvPT3G0l8tddEW2wk2waDTHt1i+4tlgn203cS
KW8FG0bOdlIJggGDJCfv7+r/N3w0pMQsCXZGmIaY7iP5Ps95HL7luSsRkxms3eBBu1FmppunNO+S
F8p0hPUxkhut2Gyivstsu/zpoHriO6zNWwuUPorLRlqgcknncfhJTCspLyPJbIRwH5X63ByXZzbn
EhCSf5A6HenzwTbjdDOdGex3v1vsssFRFU9d9wCFNZztyXHHDFr3DC51Fh5zaUIP8fg7xUewLXKn
knI5zPi6NljzNxv3s40dDWe5NiBvV33oVh3DoeswJ4Idw9c14yYPAgeSBt55KWRxZhFLi3G8BTyC
9xeaHhlzoaTkWtMGKfWkC8wnM4VBa8HyowuXNsx6u5+zeU5Zx5o+f/RhB10gJyRYQ1qWY+0G5rDV
h4H8Qqnlx/VVNWKICuoJ01bIvd0rx0VK6E318EZgKl1ihvq9aV5a45/Lf6rnFrvOMy0cYJYOPaN0
JVN3nbD8XcpaaDzicgFjSYGQpPGHLgzLm/HS/WZLbbGuuCccC293TTvoEisiVmibB2Y00RQMBv4M
rMLXzBKIpRgt0CFrPVWYvdgD1kCgzXTQ3WClWGQPG4AFqdOecxPwgYKXQr6OkkqyAVIAa4eKpeS/
apjl/cnZYuiuVGcBiNvLYwrSHM1lWp4ReNAppEXZUbe1YRD2iEbaLuoiQ+13aJlPkoHEaBTYgCpq
/Y6XqJNjEJF1bjJVASOzf+5qujQkfkyZqKj4MbHdi38MGofygYHDCqQd2qGazF7y1rEuteKzfmCh
qUGizCpRrUu0YcPAHd320BFhAHBq5ulxiQ+PffR+caPWu+srWRPLaZm19M2NQ7X5WNKdXU29f1ne
mrygnYM/5pS3fTnqg5upxeziFgtK5zypTgkmtV0nC+HT8I+veS9GwKFVGzf4jXdBMYTQp+NVYT1B
GZTDBT2uaHvt9sHVKh47Z5iou8fGFAx+p6scYkMh2klLp28K++wExXunM20ZNjkC0hJ5avLXcfF7
1TOGo0tZxzrVPoJybJm2PdpRLgytXWnNLQq4N0RU77JOIrXkizD+kzsFkJdtOLzZAbOyKowVds9x
n6AfrToY17bX+16RUNOE8inBUT5x4DaO71wiev7gn3FavkHz489fX9KPG8kGWN/fpVMWzqrMykGG
CDTqV5ID06w3QZRsewbOgDXxveDjxuaZewCXjlksBI0aWTxgNKL2jZi4bKETQ5V3k3/PhjmRIiu+
3ThlgEMJJ5d4eHhbdVp4NqXlIFB36oRoxukWXlcWlaWf2fArhmiqg8UYEdeh/XIHVlLw/GuF2lbl
REvDC9xHn4PAbT6Jk8MZepu2eKuwZHILzyJtB73v4rpcWMnOfppNdbhEzjj7PTkTpSY0fq4FN664
hQInyofHSPCK2OZJO143OcuXGhdP1x9syuwPaFuO6fcjrsrMV2f4L0Naid+moAcH98NlwasjBfGd
x6b9xjn8bUokrKViiNjKv4kPw8kbFnxFPBrJ0XQYHSnC5qYjd19KW10xTpHRsP3m626bTfrTYJ6Q
ezoL/3+Hery+IExdxop19zyWxQHmX7LLfdwWzP6vQIbCHSNZoVoTq6fiX4ey3OzuNG+2I6Vrd9ia
28NMsMMgKrdZFOYvK3vhs7p8nA5Ko83lmaNb1EC5UiaYYdKj69XUP81q0mJneLiTnbplUK6VWR9k
ZKaG/4T2ei/FuFQXV7v3DAtklldPPUovmdqWyXPAyYgEqiNEgbGciXzvuNOO+i2o+JoV0N2/ZqwJ
YLqyxyG0HmqFLq/9g93eVxtrhGYaPdMqa1mNQclab09RO3mN8bCXpWZH2X58bU32ZI7sSLeJZaDm
AGHgpxgpUftxPX+wnKl6blNtMdYYgdJpArbVerVRB/D4jcopBqJDIDRnWd04pA6HFg/rhD8xD8pF
PpxoXAORjJIei3DJLw1GmQC2F22j37dgyBeffTjgQ8Dces+J4zYUkVdSEj0C5uWVTKgidqrhKWar
Cfxuv8KSbNlor73gu/BdxlB+3Fe01k60X0hZcM4WfrdfUoykH5w7+f3I4+46poWoUPgS/Ez41GRp
SxnoqvEIwqE1B0VxHOVu/uFuELGa2FpMLJOQXRyKNqOLlSlVtccUHqvEKlkBdqujmz0n/y3hjLFe
UrMvZNXNVRT0hwmRpJss6CHkf0wPL4iNPNqrN1EMPuiudTZ92ijTeaVAPN3ErK5J3Svw5AIhdoEn
kv6F2j1l4IhuonP/3zEChXfi83gMzCfnCeAQjx0CeYdfu5lP7p0HR9ZyHBqoOyy1s/VJmHrEXNdw
Wl4JBj1FKBYOrEp7WFIOiyQySq8YUdiaYZCkscRxymD1mB844kkFWHThycvSU8iimTyz08w9KN4E
Utk4S2X1kAlczKPjfBj7LC1s5orlQZcILAU8C1UQdw3Oh4yGjF1jDh1NYdxTiceW1oTv4UnIfDoB
MBna0h2bV7A1XxiiLAwpvzKg45nvlG1tSoda9LrI6ItjEsvo7W7rCalwNCtJjVpRRcvhxjoRpLxB
hoiPHTjT6Rq1CTcxd4R7j54Cwjmwq5FY/OztCRDYV6xrMG86UKKXUpg4mbWu8eB5Iezej+huFu0F
6fAUo+QxbvivYaPB97Upaf8n9+YztKXZIO0aVvXAXHxhVMDUJfSxSYmitpaSA/ENoBqW/LZcYXj6
AZF5l8KcGPaYGceoo+grSsCpLwdwzNslZ7h+vRndn+2852wBIkgPCe/Kp7jw1e/0hHcztijFYoXt
O72Bt4J1IJ3WSenOPsLoPOofjzDWwcxjOIiR5aaocJ2yjFsbXc5/vomp6Q30P0yn5mw8r78G+uWm
sWk9cXg2VCzAJBH/Q40VK7GouS6IypOWgYGyYFgKaIB5PL/6fs77gEMFgEIbAL8EZ7Nc0LGm1It2
YueM74kNtRcgvPqHUtWzwIYmo/V88JyOoL/bmh4mXacVXXOoMREncejmEyyor9H+bl0EnmpcI8jL
Kv8Aoy2MZ4vNGTsaMDi8/e1PAGCZSdRbfE8yKnFDolnp0rG5LLNZvEwnV+GiwRgDWyqWOQaqOsAs
PxZxKX3ErC3IyGXpLFFXdQOwAbRYnsLMdL1btjkCTmbkjn+c8Ek8dhtvemqLit0QjYCclU6ERfZ5
ml+/6Rz5cVlx+5Ok6GjGyKSskXIQ3pEzIwsa7/haSDhgnOeqVbgFIAsAYJQiHzCeO2rXL5zp08KJ
4XI+EXndc1c00sfJofUSTX/wThGS/cjuLeuWTadyomeSfmahzKHch0SKPDkTvs21Z9mf6Xc2W82a
T1qipyB4eVvMyuYm/8tYYiBJd3oJilbkMlKdD0KblJM2KpByOVR7DmwYRh5EpGItmeQP8H90D06D
ZtrCMB/6kLKhH65zgncEZPAnQ4peNTUGrzXOW99AxZIr/eweDCpOTc5lu/kQG2hB/2M1UNp/5b1j
6eShtFAfaUfQKPVKSHhqb7/sPt5HpDlCyS6J9oGyUNdIJEl0mnVhraPmW0D5YjcocBg3U6YCkU0I
E6TZTr7BKCILw2hz0aKnsyiWnV+9Ksl6e57hsVmKD3PDWKYJj51c443e6s6jfq7pk0yYT8Ps2BMU
cu3f+L4gO/vTddDs8qHgF2kgtuPrVyNkoCC0/pfaH2QMPMNf3Rk5Hn4rTGlYPuzT0HvbeEo6b5PI
J5G03W3s0+hkBkWyElkpdquuoYq4IPA81kXoCf9XhCD832UlSc2gABlV2yTvXlewOOU21rXJTGrt
yRB6EShHgM2uxLdSVwN50Mp4gg0OClmlX5c4f+17318ajE9a2Iy6CJBaz8ljAybjJSPHzWb4U5kA
iJyUd6BwszgFoofHnb7Ziip0uyplq0CLIgtCLrvcZVp6Fneu2va69uwdINR+xmgaClLBvyGdSMC4
Vs7b+JsWOgP0KHVR3Cl/uNZS33Wwv6znTHnmuGPlBumtGCdOMpd6waWVsXasMKT9rh4BLyVFfBRl
yy3P6eMPzwxGydnk9HaHtsCy0XLeUw2BvdzBq/XWZGoTnRu34ZneanGweh4IFE7XFNRquO7GgYEc
QyRC1obkAhmqi9p+RiheLa/r7VpSqM3Wp39QkcRBIi05B6DNMefFrCURhlJh2PgQ0F89kUEtfIpm
meNZpG7VTSx2ltBn58iroitz6kpUIY/nZVMo1Qu+FF0ftp5fOKgakDcvq3GR3MZjTDNGwTUdVvJ0
y8DqCIbjdnkK2COuOayXeLSeDuH8TPkTtMAMMyEwAJLo/2DAqdxDVB4At4F6kIraJT9EgD+0NSzO
QtOLV+COmByaOVTCVJ1R2xR3+p5nlBg3Ezdq4fkPpX0t+rpTIcrpr3XZ7dqVryWVl1gz2nR7lQ5Y
kCXkreBQnnbPfNkaPGbmQRndJSWo3Kb04MTceYMX6d7Y8hedCveVFvtyia7qZ3/uoNJFpdxWavsY
yx6p9MbZ2zOHoNGzUQVW/PTZSLAtm/QN08Lar7RUyQMTT06YYZjgbK9fTaunHsK2KYgIK+k92Sv2
NassDuCuh/vuBlBht+VWgQbzTwrPV1/G0jEu2lBL5LZH1FY0nAr4pqGFd0Oob4jCeoBXSxM2JWS5
V4PmdGOajP6PVOgiTyuDTMwZzIdAlmuGY1LzHh38aAXieYrLdMYClOjgWlV4IyLJl0JGu92AWgXK
Igxayny/xpHEJkt2OZh3hvNEw3vM/G0P+8yjFhFWgjpD8gRPclpOUfc1VWsUU0Y4V1agA+p8t+tU
XObpsuuHfMCzHKDTWPm042zs1xeqhOeiWESYK/VTdJh81MQAwuTfSIi4L22DADrnkTMp/AWKKR/s
Edo9b/n8VL4dpmphv7uETuMOzSSmi/7Gz+1Rh9/2dLlmUzNuPkvwJ19jlknCX8ZoD8IwOaHdmoFf
77/nKpOaWfFh1KInHAJEpfKAbkcbTHp4aP68wwRK51rcIrTBmMelluPLttDQ4aPXPMOig8ieujJ7
h7MHMlydODOSppRa8W79aWD94Hvs2ReV30uxshPP1fcKBvaiXFXALSSXJOm9nRa6kw1PEc/1ALKX
oTvVZVKHvVlN2prPy6L9IEvf/MsqfbMU+psCmw1t4iP6sOUpwnSg4gVJMbymJF1UdwfJO5bDWhwV
RH5kOgdzLeq5vYYtea8dBceNATkFg8mGBmh7Hhfkj+u+h7Lo0mnb+tSZuKu+MYGa5MUgj9jxxx7S
zC0jWGnrCA096ukir/idrPTBRmDPw/8nSIyLxyT01kQ7o67XzGkLEXtZLOwH8ZM0HRNR5vd9aYAk
TB1JLfM3uzbZ6af7DW3va2dxx9qLyoKi4JgEa2fTpcaS2qvRVVgf1vyp36CBi5aDS1EstaTaXei9
5HxWnrCLLeZNJbLZ+DPol4v4AT6kl7YG8bERjOjOaHe6jccUC827pG9h0HehzZbLpyAP2vrQlexc
5PYXqGwZJgYgtMKtIKhcNvdCcOyZd+JlhMwW/omYzTk0hDVzHhxUMHEradQsJtT+cKiTIshJfu+f
TE0gFRq23fs4vdoHRGPmM63rgyqZLoAHDAfW3NY9AKaedTAAJEBBJdi8MkS+/8nFWs1okIdtjbtg
OeH+oUEZk8oqYzpymktzKDGOYu/aU5rXe5nBbqBPYwIfdoZ7vxjIt6VC9/MGEdDqqPwp8l2bml2A
Oa1jYlhHejv5OS1c1ic5CWWfLJzo8BTZWz3u5gpI/I1E7uFUBHosAn/CEt1PLSiTvmWHSXNOTt75
vFwkg2kyUT91amCKDlP77z5Smf0M5mKHRcoLytVkuUzchwtjh/v7ZC3CoEjTJZqmxscL/fn2uZJY
DarjpghkXxSJyYfczrYa/a79V7xpKnawIZ4cZQ6FcQyoyBnym/cejjxbeHY8OZpxP6jDiMCDHJIe
/j8Tf4O+qb43UYyaue5Wg6VkC7JKKD+2flAP4z0O8QKYMgDLV0g354DpmpPMTvB0l2WK4lkky1GY
dHuMtsmghiVXOVNIbIfJ/oTGUCKjMwID/VvuPMCW6b5jYIKCHLk+wOMqBK6jK/9u9MOuowT7ea0R
PRR5lf1kLLyDwv4QQBy/LDpS2NgksiydwWHCSH+SYfDsC1GCawBga3JtBVaahN4qVQyCqJbH3caU
1YSKaPHv3rHeN1wtkS5Ty2Plgvt9s/VsLvPgkxStnRhy3pS4UGD56wf7SexIN1uWb+q5ZELw+FsE
D/VRNT+zoOnOpDTPfZ7iAulR4P79HNgn4jV3hyQBCz7zRmg/JgYNbAGQPjSwEO6MDKJah/biVJn6
/2mPdo+v8EJ4rISbwGn5CCvljMVU6Ml3hXzJzBbgvbl2lOp/L1/nGSWKWmlse0EP+b13BYX/K3RK
DoTlxL+qUIUhYnJvw+La2rCuGPlU1wKG7gpbdpG7MZmEqK4lkb8VajbT+CA2bi5zSEmY+HVnT+o6
fRHmzcL9cSVoMARvQOMtNxi5dTYJ8RveZ3Gl2J/dTXrtkfyQD81ivPVdNttjamS/Tt1W4b0YvUZR
KLeLbFY35Nxgct01DHkUuYzHlSKC3sGdrPZ+SF1jIsrMREpsyqBJMW65z9kEktJcLFXxVeA8oGLJ
dlmoXouiaTajO3TP3clVXGJyB3HY+7q6XDZbvMTPa8jSMZRm0mp475wm2wiTX9dwIGddLDwQXXt8
RPQ5UogmYECUJ9kEY/DamRePYxuiMhptlGpcJXqO2dwyeNgpuv1tl7Oet+cwwWp0aUWq+l8otGOn
325tFh1NIfS2t3R3gV0/Uu0OIVOqoPo1bWHt10eYihcNubERsnIxN+npww26gP1zntLQw5t9vnyo
/vlcUbIBux5VvZ2JcbHn+zTVCYbH3O1dLS7nFZ6zEK0l0FQ1Au8dArZDhXIStotahBcWRJagA9Fo
iHzP6e1EOWV3DAidPU+nIed6QoQeJuzfI4Ypfsw6UPeR91XJgzgNWsOUz47IknAEzyIG4sih0Osu
2t6HS9Pd+dmY0arjIZulayvWZt31LKkmK2akeEGUQ1yMEHD9hf8+/HF2oxO+8yuNmhFbEYnH3aAJ
Jnrl7h/r8gOGqyPWUBwaTYfLEdBrFJuio4oDw7vVTPR0dKIDIXoN3BzqZMHmA6YeAOkUkkq67bJt
7RWFe/ZZNTqe4mFhBm9MuR8cfEJsEVgvRzskC2SaqgJ/N2QgYO3F6snSql+l3w29B6WY/l95mfwt
DSihLCVSQO6Plox+6CAugiVWndJZUS/KkQbnfGIwJLDGJehFTXPqlsJkrYWD5TTLOETWbf5GyRmV
CJDZx5qHqL0zP+8ltgSqjuOgTBnnU8TSXT9UNMZgXwtMeWIH6uy4AdPZlKO4OLFkRefoLYNSxq0v
QWHpWMFQ7PTX+9wwWlFExBgXEvk1D32Udb7VCDIkx1LVgfb+0tfPi90tYmRs2u4KHoYMMXqX+qvC
RKG1jCNl6xjNGzvlHTf3KXBdNYBfjlCW8TkBJ3srVt4cm7dxYHxAfHGlHBMYrzcFNJMa+6tCZpsJ
G5+DVAT7N6YE7WhrjX2PSJPEu+koyWdhjjVYDmHUAtGidRSuNQkWo57QcrR0igGikghxbklfXzry
6XUMqjrOmoXFEEMUAWGScF8/h9t3tkAHXTtw/jTFqVEy+rjqQ2j9HwmbfxhRFknO0xTwj3LOv+zX
A6MeCoGnL4ckpNgOu/xqgT39Tn2WtITuaph+ZOAhps2xwbWh7Q3w2GzT3gLIIkNlaiDuMXMcJFeJ
sBuJxrJ1ucufbj0yeBuu6kf6K2891bDfUQ9SLrjEzGbRJGrWmv/2+Jd0COMfjHxl+c7wS2rSJmiV
RuvCHQ59MraaOQ0UYBbVxg06QmelrE60ruczQZA4HkN7XgmRPeLdFlmngYp320Zc8UE/CLFKApAc
gF2SGLllJxMsGOVCLT6MZzSpwTZikQYeOMfn8KHoI5kh0gnF7txOyk+sjxqimrkBaEubhGaS9GFo
beknMfNghexe146EsT+MBaupp02CAg7oPwl6J1C68AYQErjSsxx1x3+ni9aT6EmJ1bftBMqBGJ2U
ICM/njv4Ehva96q9p5c+peYu5+UIQzH3Te2U0XbVLOTslZ5KFl1I+Sdq/TAchLjQQ2PPm+4D3yPB
1Io6XCBhXFFr3rry+qfb9mPO2cco+DScy3bk+I+UGHSR2RmW/mQ69W2P6wXf9xPjgAEf/qfPIgtP
yd114mBr0LKwG02aSCsTu+JFpKnckKD0IztvmXCveiYiVBl8i46pnMnAhciUBKcjWfbtTPscmxOS
nmWmWXKdR8SvZD47jg3p78027aiiMHd8y1j8+083TfQkgVNi9KGyAjEUguDXQgmyyCc6xjA5FwMM
LVC6/YJ6mMjUpOIgaeehuyvqvPsN4T0VuacpU9NCjb2SPkEmIKg0xEcDWj1VBQMWo2SleuL3rP6N
e2kCRU9TPh2dahAUqjx0Mgs5T+jFeH3oCPk//ztH+iJ+mFgTQhpDAX4Z9zpnrUR2R+cigCU9s6tU
0FGr0x0WPRGaBX0JFqkvTjyJFJnis1IolSjSUHWiuN0eBabK992prEfu/kbtdNlHjZ2f5e0Hprjh
P5JTgwj6HQxnk5K8nEgW3P2GaKWStP9g2c95kw4yHd8cIrJaOjZOB4IAlJloEjisUbwK3oRXvqLD
7D5SvuwN5mW6X39UP6DYm2MNTTdAOGQMqzM5R3pNPBkEe2OFLkXQBccpqrh/UkR3dRZjQHp3Hd8v
5W+HBMEoZ7apgHzjz1ZPvXGXMcgQmEXEVDLuwiKTBKvsermiQcrl+BjopOQrsLRHLjrfmSZ7HLPz
acI4g+W/ZjRrBAl5FixLT5p30qXja5SMIVknVZD/JN2vBZK6hghPSgWNthSM1zGpZlJMg5j/DDux
aNh0q32OQpFV3JRUwUPgxHBr9NkBvBjNhojQp5BwWHbGBFOcqzOdadcPuuigqNd5aI4X4kkYy/Qz
v6V9Zinly14Jd31QYDX7jZRnohFm70MBe1KrFXH8cgR3AHRrYKSCNtn6YFlSyEAxj9Wy3ODZZZbT
ghPYzJHWIULe1ZDU95nsB0RXq5n2CLx9ZKrjoXdQwb/7zGAbdL20yZ51ljPt4Gv+cA4RyCZK4frh
XoVYoGK+eaPtZjcuIlYRytBR3nUJdbKjBrAU51GChtxO6rv2u0vwjNiITvHc1ebHc0BzXDEkWmyh
PtELOZCftJvnjg/6uGKbgsWvsrrNEuI9ESb74SG/SyIEab20OqIbJ2MDt0f2ezAdj8IgYSIw3W9+
SN9aJWHnXaGh/3X7RLSQ1cnm8qDF1H+gl7QiRQsC6/sJnUDhKJqum7YydLhGGrH3PNSxv6Y+pj3d
J7Hd7g3ClOg9L/OATcPotPGxGQ6wGsAbwclheHg5GvL8zsKAYU/JS/zgXk426XFax0tcB/9JuK5G
K8bxqMn9bAzts1ayBLIeVSMvo8WG02jN0qcTdB663iDoPdsukmPaZi2phYgXrz0nXpYC2KeABvwp
ikVI69uDYFU2MySMockC+p88NigvuwyLSiZzckYNQWr8USq1/KGyixcmmjInGi60qGSG3DXLgwRp
neHKqT7owXwp9QyBXa9mQelUwxurp5y7uXYRYWF8P1aICIkUPYm1i5THoS34LHetzLSXZWoetDXK
lpJj/AMMsynsHsIvSBlnPfABCP4fLrEkxhhc8c+jqbH6iADlPPNXKBkV/JB4eHcfZBflPBT7cCUu
09nmH4nYqxZJ30p0hWikm4H5KouFVgKzj5TTtsr2u5iOFZdlaxJi1gKqeuWRWR9t2wIGiSvTsEXa
LhHFF41j+3gEa1QApUz5QjCE87p4xfKCo7RcLrY7z5Yw4a/XFa9k+wPxP7IXg5ySIIRlifTt9uD5
7NHzskxAG7OmWz/9pKhO1xQiD/6x88W7DeduMSJfpwP4pQaMfHIcw4R5RzvcEEG05wu8O5ENdcX3
qCfupq6maDOgp65ENSoqvBQg8hrt4fmOg0w5m8WKNTssZSIDxUMvQOx03vFI422XSpse9t4doUfa
Gr824UVoA3o6vbgCONWlVG3dooO3Tb9hxVMl43Q7yBvApj2iLyTFet4zeTEtQ+neCLE8JXwOjP6W
w+itN3IGGvNpYM6EJx3npFXRySd0yq2ArPdpQ5/UW536Bii4jxQv9PIONZgLBNFtL1sSuedhf3vW
/r7LS5CTIXnOMeLfNae2MlJ8ZgEqzagdTX2krqVClLoT1EA368HawtD7VDmMHOQvKp8p25ESrE5i
UvZizqMd7lzxuK+d/u6gIepE/VnVJ/OfLAGBneNghXZb/q6RHPvsow3xC0OxnjbmThFfzM6U+rAT
rvE2fnyS7inI6z/ueMceG5KmYtHH/M8XbDT3KotLYulfsslMQ6Sjne3ctugXKKd7GDpXc737Ntdl
gSOVR4oEzAKUxvbbQq2kGYyD7B6SU9ya+iTQvmely9NnIzXoRbswpzpCzfOLYWGu1C4PXn9Hp/XV
ZMACZ/N3wu/epyTMEa0BXB2MHqKS9tHhRqkH/Dz7hLuoaAFuWbeK2Qu6m5i1JxMDFstpKgfW3+1l
yjDtKYOovJ9g69VlyUVNp7cJcJ+P74qytDm7L6gZqnFG19j5ubq+KbDs9GjyaltQMEoKpH7PqgfA
miSmZzEIKnagfK01L85ajwAdrprbPpAfsZisF2p4oxcSMdgfpsSZEdHW/xFSYB1LB0bCbchqg1Ps
XECXX15l8ZNa+c+YNAybNGaTXLTjQKFUTr80NKWGcdfsb1RRknwlPR3HPiEFLWJplvQSH/89MzaX
WP8q6kg+YpgOwkhyV8A7pZILW/X/YKdPfTafM/TBAhqRuYBReJE0pTJSzfKkxi52NKnPi9iZR5KC
MWPTPspGFegIY7CH4w6+Xanz548lmA627Hv2eCNLhFttrqYVgi22K5TJwa1ZzLqrvtK9BEj8gDC+
s8y/3ZkgJdbNiTo3HtF8OrXCeXZO7CGuAvRRb1Ga6wgWjTMGG1wPpOXijfNgpI4oLC+21J/NKD7K
BPnaLzFmZQvaxsmMOMLLRdetXik4I4U3iob3sOO98hzJ3Yjp6joZ25X+vIPeTzroi0foo6ozv3Za
FGEdK3aZalTxH9esNqP6IePmhPp3JlQ4VKbSEWCsRnr3QOM1uOD/qvomLyE6x5fwEaTc575IrCZ0
Blp9b6tseNOMGeCHtX75peqdUpwHvlRkYTV3uvg5ImaaDMr0ANI92iWc/7Jm0/HirnHKt4Y/MeIA
SPvSzMxBRUhrSh26urXj60nhJRR8Y/svaVEDrwVs+CexgECm+Mg2Q3gDb71JCkmcccDB6Oj9/VJj
hYOyoU86lhPY8MzVBpskIvmnTZ3fl0DV3r81K3Rp2dOhoqNlkejZEWaW+1q3Y3Y7fAsZ8Kfn8C4g
kFSp3QwhMyIyDlrqFKP7BKDwlr1nOznxHUZWwIyIAviyt/0LNRRqD81SmJ+kl4HKL6mS7+4g5W69
3Cyl1eW+slPQQNRYGGCE26eqiuqbDp/VrCfQlRNdt/VaZBbbyJSrpLMOk+xDC0mYE8gRTL9CWFWw
jTnSNvJSSJAekOwRoSVnx1AhIDtBhPVSLOZZHH2n4Y3uL1qRPyeRNTJo+CZ0G8OCs1gCVAH7vuoP
2l8MpRyGcu9LaXUxT3DxaCc8WDmxqM20HouRdltCQbKM4ej0aarLus2Z0YgDooh6Ai6qymz2l5Yo
McDT3X0Hjl2NtH8PRl3UUV/UwvdKMVsxiGOkqr2ArlGdYGrSU7aJ6NJifH/Px/HiO5xc3VUWP5W8
pyJhl3yAczpaM5xjwPn2fp6wmSwWEhppawDQBgt5GYFUYOn/Cn41p7X/bygDZIspE3Q2SjAuMR9M
G6HbUTl5h6MoYDGDALo6+nYitn2jxBNiiTvQV5m4+W040n+mm0gYtyi+6R0cyOc7Q3H+ByTtKH09
cAHxZiA3mFwkbmINXWdy0QkB4zK01ZjLgFpGDyuVp6YQItpYnt/4H5QpPwpH0qOIzUB7kd0MHWYn
S4utaXPeGTwtP22Jfjcmf3S46NIQsP8z2V98PXJ+gct4JHpqyikYwD2NfsF+ORjAbxzYfHm/7O2o
pXCUbDM558/X/NcyscUPkMjOL19qgj0insSnOkb6adLTuB3zdKweMf2FFdHJYNYIGAAJScQcawPZ
z82+Z0qIvnLLdHyT5ITNlbzCT8nAQaOmLbS/7Bp20FgCa+MDVUZ/rRtTgw7f+reqHrTefjQ49KVH
LBUHdLrfcFeQncSdudYOMMOkrF3J8SMyruf4dhLA/idmOFfjEXAGm4K8abtKlRK5MPSoLVEyTsSf
dTBN+IIj8OcZdJV1sDcoqva8AtYVPIHJ4zxcitkiBG48fj1WyZDJHhTk7pl+dl9TdMUGjehasGRA
KT34aD7J4G9+I5s5VzAPYVR+bYEB/gTf2RsU4TUWOyGhEjHX1g4/Wdw5f2yJyRJIvb5O07CNcw3l
635voMY3X6eS4WhBNKIyC1IJTIVYnVxfArOV+KojffASWOr44/MqgqNcGols3Fdn7oiwN6u5DWGv
jVxfKTWh+67f2N0CiAXet/bzhogPyXRYSha13YQCHVxi9ikfBhcwdpHMuA8SMmKztGLg9Wi7jjHn
5V3f6I4xPvDKB753Lb7dY7zJBRrJ+fNWMkVpcXf1ZvWVg3BOfSF0396sr/eppqmRdZyfmC/C2Mm4
W25rJsbU64QctYMrs0GtdFKR1Nk2uAMsBEU1AuV0IQ4o7csmeQUrc1j+GE8eXKMKKpH0TWFyZzVf
lqK9m8V7xBSTlnJ48UEip8h3ptRCJfgB32XKnbAbYZaR/KLAPqK67AQ4wbZr8NygolZy2DA8dCD6
1k1WuOfqP7fVAJnkCB9xNERKSIGasyN4sMW82m8Qe/Ht8d0B+KlZm7JafW4y+ilFOORcQld0IbzW
7+cMLifgyANht5ux651Xl/w6dEGtByrvw/0V5rO8uzwW0sexe5BIdOYm7XR2TPKKiFY68a/PVdFN
p8Z+F7PTp4B8x26KYY2cq7Ae2WAATrECfreCscOhrRTRvJfUKQrzS7dpw4kBfbOVAayQUCfoHSES
wX4W7Io0iY+Ts2AtbClYlYWkw7fERAodrOm35PP4fFXVQPe64GZfFRsVBheEQK7Dg3uBH0RO80xY
kzwn8GGD41eZ90sBslOmzQHq3Vylhk88+cBa3B4BKACkk5LeeublrMpalhwTbYibEOCvXrO9VPVe
12BUUs7NUZeWGbXTn/Clq2kmoY89hd5WXU96X9aZkkgdihIHHdAg66KgunxMI2MuZ0RUZRDFgqhk
/WymVp9QxDvYV0rkA64B8LVBdKPKJVR2RxfGcWPNizN15Z1tERSayJ33KYewiE/ayOBTwHoYsjNK
tkzNbdFWjMnNVaGLzXeEr+4ia40OGNw6katQuhoX4wjfAOWJ2beGahen4neS+r3kvEvkLHHyqsBl
Ol0y7bPIcMpFNRV/7QHm3sh4jVRc0u8fdWoL9A8mqKBeptem6A8l9BhExSWBva1NjizTCVQGiFGs
DLdDGiLLSEYgXID7kS8F+09X2QE3EJUZw6PzIwHzWenMJdkOpUGPHpaH1j+gKVQpio3x0Txg2q4y
9jzLh8J4vxoFiKt5gObQ2vbzLLhYHURC8IXPdMI5DRh68ccwYsxrny4NUgT/+8YpszlwBIiXNwib
CZpPEhU4SmnTkQQPQ4S3z822epHxWtAuBTAXMKtSnxHgUAq3naDMEHOYzg8sRCUA3nP4l/Gcvugt
20iGIPgorJ/ulzLUdiDYh2/9b1YWrhIjn+bfnWCrDtOdnUt6vj/7HYHvgx1zoCq4wwQS/CoBjLbD
0IPvS5NAXAiMfx5ndcJz0Ly19Ek0BAY3Vp0yQ/PwQVwBra9udOk9e2/EzcB42aRqgAynl3d35uDR
LynAemafEECFfGRxO3Pt8vd5IWKUlH1DDcUk0P3xzd9I0VyFw2tyMqxD8ZAzJR2qgTiaKNqr/jlr
h1KrZBMGKWvnOZ9I5fRAyFav5bSTT+mf4Vw6I5SVOPLgvW1bfDAdhfIxc2qZ0Xa5GYypIexSzseK
rc2JSp/qJuDgMhsHwm9rUDoybafzAEdmlAdR+5pfoqEdVg9BdD5v585djUrRdkVm8P7dZ14zgzKB
NRK6RYVG5/pSE6ITz6hlqmP1DmF5Ns5EJ8aj22aN3A8s5jA1EoRB6CGf641dPZOucM5P1SurrDIo
ofo42pBN942/birLagxN63tIDry44rGkdHpeh5P/a7u6QGNBhGynpouty6hlTmgG2l81frdUNifV
+1Gs3zTQY+fEHQmLSH65QcOP4PgiVqdzVKCK5xhpJCIT5X7S4BRt3pTiNV4fzt/8UTkV9boKquH2
i/v+TXwjL5+sZsm+W4YLEXr9NblxA9ClSTXFZfDHWbcL0YGS/O46RstPblQpQdfHtZAHak6F11JY
EIvBkyZPq/M9GpshboCVYAol4RX48qnJ2F1MqJxyegBJ9TIYLnYUk5IfHlrXodhZJhl0R0rWIeme
h+DwqE9QjQeqJ7yPue2pQfaJupMr4o1F/arbZBbSrVAaAVy97h9r613lmuVotH69IRqqFRxXmwQ4
FKKEffI+febwKdHlfz9YK0zU47Bv767aWqvxaigInxn8T3RlyD01eJR/lOKhCxL9vJmFxWunlUz8
K2uOayCjYQafnXJ9bzbp1NrO2em4vQmN7r4lIaUh6RFFtru7IUASnWVQPscotBGHoZProQNOHRq2
LmdEmO93nGi7XbGHFY3IFjHm1mLV7GN3WGn/nWrfnAUJI21b+qf2Mz33mMwHCJTd9A+b6v/rEGFa
fefxQjczmZeS0Wl8SihwHn55e5NodrPvzFXqa/+i0POTygtEkd5+AjrtGocQrUmO+i+JT5fBA6nL
nb3fNgSNmyQTH39qqE7PhOnJdeR7aZWiPpkcLRYrpJntCA+NcTEWd+YpxaINe3QxjdffJ/bnjPte
GXA2UT/Zc+6wUEYGeCWGulohwEQ03lZj4h7NrwGudzlWJ6ENDZ480Tr3C9wEfqyEytbICTLRWBhr
XX5ULilqRH4w0nqILbsBz0yrbVTpMx1E9fKWMB/bfjER8ZdTHoKRvClI1b0i8HUf9Sr8g90LTYc9
KpAn0s7OiMx0e/EQCrQkpXr01wdzMeLCUMFwYAIcryybN/vUJtWCrWULwUudxQ6WmFDNXzdtHDjK
oht/bbOoJYsOza5YA1gQIMscpfCmkoG+s/b5FUjG61qLFF3TjJv/ONl+dKHQdOdDpXbDDQdyJy5f
DctgO6JPGP0vLsoZQWGx4tZuypOApJ26JsupFujmI12jYEWBGhu+44pu1jzyKGA/FHozjbEjUvR/
7Q8MATylX3uitiDMO5EXPlADlfG8I7GNWpHCZRtPvejCBbb9mkjxlq/ov14HyVCsfHkRHSi6oavk
eyKOENjErP+C76g+qA018lPt8/bRajkRCdFW65eVjfL7Qe2UVJJLLOyNORRuSdSU9Ov+h8jyBlCU
NJTMQdB97FMrDGopnIi5Pa5ZyprTXwIq+TEHwHSi4Gu478o92XQ+H7WumYBBjbNSEeoFI5NfYPzJ
0sXcFW7xSGrmGh2VrPcHgS4/04Ws5+K2/lxHscrl/XLl9UwRsKFAccXkl5im067KKMVfmdZUor2X
Juh5/SsrBLnVr/G1UyJv9fjbpzS2q0kBcv2t8/WWyBSihqZqnZ4h8XIAliwmyZaL46ONY0iIvomp
3agvHDH8aP9b+t85jsgTAEWnBOi6CwM9CNTrpp9RRMLZr8poyjCkubs+QxV4kHi/UB6vfXUJYKdo
hPHoj2KHEQ+DZEknIXzx+i+4cxBjzHN7mvkoteOxanWQISfJPHruhC0/NjhTtC2ok9dAOgE7tWnS
sERk4AdaiSjg8q31k3Vw4k3l6BFJjIddzx6WcXcGy5bs/mcp9AHzFXdqGEgU4I/imMvXL50f5lQD
VzLz9NTYRDmeW2GrPYq8hNAj3mIiiIxqfFx9gKF1YBU0T1CHt5ZHYwNXPCl0odFzkmQ8PSGTWNmT
LD1+VOYEuFP5ToWGkZO5Yz0k7oJxITsOzbdxQPQfAjKDAIOheYyr7vmUcJcBW8YXYTjh6gZP+DwY
A4xBIu3v/iqZZ1ii7eTR3aAJPpm5pHZeoDHN1bB7TKWu/G8TjlFHYtUeuU75vQwh8NiWzBR4j+6k
F3z8MDinIde9XvljBYvs6wLXhLk4TMj4IKcChVLm663z66ZGXSl/2Qy/SZ6ip0/rBfAv6wewEdig
RbxjSCn48Z2X5x2E9JBNU8tdp4agpkn4qehN22IjO3/XeNdpAFF9cAuLcy6QVtuf+3b+IRhnxMbq
H7oytQRsszY5qm8l2JY0V10em3N2ME/opKx74GoS/CazPgWYTSnhXsssgrNZN0bfG7k0d9resybT
WAV/yuGKfB4z0dVLYRwdgxqkE2UGgAsKiWoGJDAB99dMTdaV/OjwUuS/zTVKiaIU20bOqGawqUdu
lZUhO4PTv2aUl7ymejelkZ2iCCavqud9W3jBScbxC5jhwokD+UUEPsJk0x8URn+XOJjOJEplaiDK
7sD7Wat7e+ir+PpzLsA7ga0FRAx61xOc5pgqhLy1fqyIogyv4sRACxTphNuElslQKpoVnBGBzGx3
VRGOUFItUcAITe+YDnh9imtt0SZ3Te22cjUkU3W31/oAQWQrtRIewbGHo5DjVmLxI4L1+1RcyqlJ
hteolr5fkwSEajJT41X4BsLPXEuEpOZvmO6dUZiS/XVG2PfnE1gKCitaHFD8uWUpqVbksQDRfoI6
Xf/N03xNlIrRth38C0yRG4mEpUUorEeeFH4uH+Gz35LOQ7BJYo0DUVGz+fqPFYpDlmtcdXhLKhpr
LQWJ/3DZOkoM6aPHqPaJDOWP4m2HGYBjYvZ0zrA0pyAZBT+T8IxqIMFYI7p2t6OpqnmJ9TG2Hg2T
1PXvio1/SNG39scuK13MJ2a9l7NloQW2EoIFxxRXv8hWz8/JkLTT40RU7gVoiWaUBwr/1rVIQPWi
qUNztkYScu/15WbItd12D7Gti5z/7bSguH10Q1IMTHvJbzm/fzl7eGY5qdgIrtGFRvUZcD/c60NG
KaaIn3lSEqVmk4vIq/cdRvywh5pUZlM3eJgWDR/pdHxpfYfh/zMOp0ZfMA+q6/y/pYW2yyUoHots
+ro9GQO6WIWO4LMfeVLOEduTi7Frrw4DCACY4qZ38VZXqv4bjTjmbSt0hrKe3IGRTIYp9mfo4lVr
A91ZH2tiYowqRJpO8tT6txkM5q26c2saC02/AZDV0p6ilKHVftP1K1li1nkL4Oa/ofLvJxKNgD8m
oZqn2u4H7MqIpOBw1bd5ucaT1GZ0Z+Jl/U805xjdMHsFC/uYs5lTGnMhh6osGrUf9cCU5NShhjkW
7Rf/KpDM1Ak5ar+ZTVe8JpulbW04XrTK/LBloC6hxDg1SSSSL471Fb+S3bHwOCGGQDodz/O2mnuV
ryF2WqzpBHRMXPKyXYIMNSA11YiviLfaxpJ8PmrmdzfuIt2fsSH3ngrabhQe1zJI86RNEML4BCc5
+F6Pauk1E85SLrjmrA/AzjpfHfqqYnazv5xb4Y8PyJ4Qr1aAckL8rZQhX8hpuYf6Okzn8SS+31Wa
6HLLdgcUx9rJUIymeGnWfH/gz89bz1dRtbNHGf27w3yzQWyIe/3IcrzzStnDI+7QY4293UmeAOGx
P5/g90Qy99pzstxKqAzuJox+Q2S5B/zTcd/TXjbZYlMThWZCg9bGZ3m19hYDnSQCPVOLvwo3NtuF
pd7+DDK5PcXqn3AJsXDhQVxuVANmgy44adXZQNtR5UaEAbJQJWxsYMZfkXlgRp/1FmLxCntz/X3D
vpZCD6xYie/yuu7qzlVN+0PFjBeZjfXMPIRpyt261+JzFed8F4/XXWuJOTtGNPuUc35irqEhZcVk
jszQuLcGU5uulWdPLRPEx9LYnz/AVVMcS8FRQOZkmv6wKmgti2y81MM06wOV5ieXpUra0VDWDS5e
ttEwT5Eu7Yp4Rgo3jDRkGsBv0/MKHa9Eq+mFM9B67pKW+/Exi1oZRAkWnx6oNi01iufcSUkRM7wF
/rEfnLzoR2BJjLdofXMt8LUzdyLPZovMPSKrAUjOJIMblQjBuZ+Y3koJZKSBpg2Bjg1+DMvv/zNa
uvykvt9OOyAKS15C4kHjcYbVnqbS1i9papewqOR8Zz6TVFKQbYwknlh8cnnwNHxV7p1Ze8pdHFs7
/8iELJEFHUGaKQ/c5SIdPV3Kv7OQ8zbBYOBdZzEa8m5of6DV4+IJkx94CmWh1hj8SiQwYIrqJdfQ
1Eb2VodGgqQq27vt+oUU8gsbMERUFO/24uJLBfTVG7LcMH8HDEoLofGDIiEy/FnI4COD5iSBTW16
MDKDwks11ubVVbLk/u12IPLojg/0eaHHZT/H3kIEsZ2vw1ZauxCvOlyUjXAUq5vvSo82PhwPNkJm
rDSweiZJtXXHIJw0zvAouEB2ArsJsa5LrQ4mib0RX1kpY1MGcmzJgvoyBiwxY+D3K42VKVMM2brm
/n7rQk3Ks/LWDgydUdWKSkdgfMFkV2W4WRg/YhQoRZfaeIlpZkR8H1zdAO94ez9HtcLUIsjt7RF5
Q7DVVW6bdVMvI5QsUbSvk+N78xhx4Acse5hz8UAl/1d+7SBWF7qW148v6XX6y7/UVOKfQkx6trMf
5rb5+vWWtv4KdzN4ud86n0N+2pIvB0ProJ0L2jU6zCnkZFLuOAjmaMzfqtnT/UhipcCnurd1WvEJ
Nc7iZMJc3Bz30M6axCgFPRIl6v6EFHI7/djuaDNcKObPW80ehBo7gr18uDkPXm0gh/ifQB24I3RY
cYCWDgz5OVTA7ZdE2ccgxqNkEAkpuUfXwOQo90eNCbAiVrEo8/uZ1wruLmz4T1AIec3MCvO1Y0Jx
tVvi7YEtD4n+BaogVLpezfXs8W4Cw5FOi7dWHgqS9D5SctRB9JPCs4LdLFRmGkCMh8dAnTktm3r/
sW98+AsEN9KFDie3jZm0Vqk5/PI/IMY76fArMg36cUiRjk9nt3LyvhHZ5ZWFbrOX9vxYJ56qVb86
4awcjwH9eEIUoFFsxkYhF1Ot8l1K1DUVmI5GHM/lChMUdymhAn/7LcyPOwAah43DBCAP4luiKaVc
Uzc2UcxXUKS4jfGH58VF11WONmFrnzMfOKjykc7bVOqli4yJ1fWIfukX3HaVMSdhBXhneqJtW9jg
DjkgQ59TQSFnGtPHOfFNkC3JSIqxvyv6d1Z9fEyAMFsSwSP6ZAg4aTCZwhYRW/DFEyeUkcOPd8Xf
tV+RrdmytqCsWWKCj8q4vpebmhCJQorjdRucmwiaCKUAQiRZA7efhAT+IPb/oaaE91kc7WHd2rZ2
Ea4M8wD008O6XmFlns3QM3UD0mQZIG6DLbrVOQEkn4MyPL2fBaDBNSGfjWtD33iKmmbp3dBKVVHE
7Dnd+DCho3IV9HhfSzgdfNNh4Htpa/JayGMjdasFAO4kB98t/uDQlPi5cGeZ4xqhHhyOyL91hvQ0
685sVXtZ6WhP05xgD6PHOkxjit9FtSlxfo9KNMP75dzysRBfU2FjCL5mDsaGaRKjFZtoXpfsMILA
LRLqnOZfSmnN8UGpxKSTwtORwzF5Rh/zh4jqZqjiGBYgueHirdkJkX0pLp/ZwVxAjnwO6lJ4e6Zq
ID2e1QAn4L6zMW6rb+JyBfRhC1M5EgMj35/cy1YyZHUq5za+rgm3/uuW6CqviCGoOV73v6OLpDPY
C1zAYaENNSureTfipO9BBE+zCb4GfgqLzJLIL+4FuxEGoPn2cpZiGOqFwd4+ymnjlTNGfol1RjAB
rEOTuqWWFBqxvup9i5FRyZhvlU8fh1GUy/Ctn0EupgzKDqE5qaDOw+zLEe1+xUgjFamQYgw4WTyO
7lGAZLYrsgDpMuid+FP2+s3EkWIsCF2KuhbjkY6HbfWjY4q5PdiNvmFhQ/PChADesL557R3pDqpE
+sYFB2yMVLAhdAdfITbtbSw8lz0EKzOv5XpdFVwIjrOChHaj1te9C7OC6QqVFVdosCORXEEpriGb
GouKnOBLC3IuuWGWRwC4u1rqjsgI+abZrQOQzDWLFdjPC/QTFDc304hokdvLtvbreSQ18GrHLJlz
KfbOvKiRDUuQiJf71Y/O8HkoT85oDf/pC3Sg/2XGz3eb0MayY8fBHAl8olC/1hAfh3xmNwddX6oQ
W1q574zMAGEzKoE490jaGSt1G3PJTIR3uApBhpNlnE727GvthS5MxYLdnJQy2Ge+HllOIkylISRP
cSYfyfldROyum7sNSM2qAiyzBW9BBdW1TZpW8uh14+mHrUpFdd3AMrHNb37EocNepaU1r4Jet9yF
xFkQrVWPZqeeeeqnenVfAs6G6pJD6w0mLdm2tQ9sOla0fpCVCZYtmHINctcKcO3fp7fkYVqSy4f4
0OtRJE7eMqehp90mt3vRPoingD9/8hT93ZEOtl1UdErAt0Qe+/YNxfu3wr6eNpIxk3bCPHB6pOJz
GwkBluTo8ipNMgzqURXl+1t2NN8CJcCPsYmpFF1lh8drADVxAWob59vXaIJgwUEhILUVz8pzkcjZ
UUKlzmh2PpabrIalKq41Yxae+7YsvVssT2pBhmytioufsEbSnmSeVRfDLuv5vlCAKir2k5a6LShp
QrdQ0by/GYOJs04F5/SsVVrCqdcn/R7iGWN3f5imRO9DNEPIPMrNKKQnfxjDFo8ob353xPFhSzTR
XujW5Nx1ZuGS4k6d+iAmSJNyfTJjXiXzM6LyZG5Plc1Omia6fGUorAk1vF2EG2u1pd4BmWCyI872
2pM2Isa6D+s16yWtOUWfGK+5MZASMovler7uyuQYzfl4WvoO5wWdiNTJ5bRJzLSne4C38TBRXEuX
iPtVv8hW+Ascwost5O3+lwjwTmBa+3gAwfuKjx3QLAxTxmv3p1fKn5uXgdaZGmtTmkZDqS+vz9nq
rNzqL9a/+6BDGt0QWMPMvnugidCpzUGFvzfi5wbQ5Z2K6w7CEVouQvRCRh+hiqhHNnwEjf+BfIec
j7XqT0GDgOtoJGHzs2Y9gm/wykGc1wdTes2eouhD/so3oH4NfnDsTD2KUys1VcsR4xN3tXdizXMm
ao2kF/vWzwNZ+XveS6AqEqB89aJcK1o/EAJFXfSTRmbJToujsD9s63FN/EHCpXQlWJSGiieMYnkk
hrOhbZrNfPhi6v9etRcRmY5GuzcoIgY4UEldpLq5rng0AWtkKCpS14kc9CforyKk3aw+1CM4sXCb
gJ2YVNHOIJEIOk7xdkcmnSNeQHYjwqmKQQ2f8sCE1jtgpySACRuXZhQaWFkfroFlrFR5jXL4uSw1
Wu2zFgTGEFBkXdXGnyhNS2jGpc+MCApIjd6qY59wUA4Nuhkv0Ku/Ya4iOtAytryPmB35OKm1Ud//
fnWkC1qGr4piVMZ/y1piXpKf5t0lXf09EAQiVaMGc4+m7MLaUhvuw0IhtImjxk6ssQBbdsJGNN+t
LepTGBdycGk2eN3lziP1Z7A4ocpSuiQAvc+J6Yhr1qdtQbvP+Pj7OQGJ7ram6LMCPni1VQcLz5wT
oval6jn0Si67EFSh8lvFY4+RLrdGaV+SKKpLi5B36XwhNJ5WuVmIwRawN6eaIi6Fa12sCuEoqhCp
3vs/EwlW4NlvE5Ud47hD2rtfcwPGeRO1Ep+j9PXx11gL3oVIWQrMhnbICLQztTgh7lTmlaw3Wevu
ppPrFlsZf+lxF+2pEPvP0v0dUCWBY9c/BzEX8qwzbaFYnqSIBVjE9VCExcpjxpdJOuWjGwKWttdk
Ur/oGi28coiStIUFxqECdA64pn6VJjBxttmPhy7ySTgNe9GpD07uU4hnaGZfQfwEzsduaH8Qm1Gz
WzDYe2ounVlXOucNLtI+CXPbzRZribzzHivruULeFlK56ra70+wS7PFxOipItqbrdkDaZMTKtOaX
DmoJt3v4aecOZjRBTqrJCeKqbcUb9sulFe2ckZ0YohxYinxlrD2diRBNwcIW2f9+Hv1/vCEAihi7
b49dXzK0HECyA2jj78VKimzmF7s4hZyp6k6wkw5TtpjWq8qbfP1McT9N8CTvIfroc4ZZrkdDxYoc
ND4/PKCATHfuBt+AYEFhPjYlQ6SVQjOJMLNAh/4bZE8GOH/FonSdrVJJIMNmEFkn6w8kqSyjAaa3
M3+G79JfvrmDGGiOrKtj0M/bMVXJR+baUUUcBT5PPzhSJzgEttykez3lhaNtKjnKHkSXbzNA8A+n
793vwZMxt8iaNXGIh+OqEHFTwX9bdR+azKWG7tKu0pe5H8XlS0QU9xo4UTIBQnhRv5yOvFfPold4
pt5/9NXLi+8puDYAlXgnahP4MDDsuhdP+bg1mQ1qlaaOR2pB2QdTjAbMaT3xFZg1dcMGEuM+GNlj
h0boEQUL3c3uds0hkOiIjntzcJNKdDASW2WvgKmeAUGQoh5bLtsBQ1Lzp9EFmAiwHCzJ7argRMcO
4NxDES7NxeXDI/y2B0yp2E2M8t46/BTcW5WUVYGoE4hvKRNWnhuibsVRQGRObnU/ZvwlkUZ+9UGK
NEU0UY+lqo26O9880v05NWxG7CFvEa6/hHR2D7qYuASCGH0khRB45afp57kLh09DBOiq2B0IEy0s
8JUA4PKjXvQmCTBKzg3jxZ5f3a//o6C9l7Jq2m2qlmbBr+tsIXB/MTwiIy8KKtFmnlCJx5+ODWN4
76s6DwE2cP7X6VP7jwwXFrl/5palPcmiq0n+jrkhQCAwSkt3GVCWcUIVRFG8RTBJXfVVweEk8RLw
NpGTi/K1fL5ejjvcdv81f9sprUYdT7GhhmYFzNy03HicAF2713MhFOWjQxo6sTr3GyHHpvAa1XJT
VSZTJa0gliT/EOZnC0T/QNNKnS1ZYxPgZ4AqxPO2UjVSiEdLout13qTSd66yAEMLCRz70B2EZveN
QncoXLUgWswDAAAcJ/YM+ZKuud/lisCH61BxkWHpsxr6XjOVmxtiRsktqzQP857hOuqqxgCThXK/
EyUqEjXkwHAmGXJQnaTn/cufD/E2UvUtwf6AnaLm2Gm05/s2lktZ2QbrU0KIw7sJ5HZh20RSW7w4
p2se4G29NBAB8XOm3QYBUZeDBIjqhWsGjjnn7Xy4RLnfzUSYikaC6M1KWgBQVxGWVRMrF9tSDFfo
u34CXyctPI2s447RHi+wIZGytGLCZVvc1X4X2+aGy/+Dv6qwIt3hjIYWElmtnH7AdTytmv//1DR1
vFdW4fNml4nhPQqxeNnHdR2H4dMx71lWQ2HD0mIyIVK40ZJ39KXuIm3t8KBRj/CyCH8Rj2jbe9tN
Bgy/YbTlkmO09kIKLVLrT+ZCvYinl8aP8N4aDDgIsekjP9XMbp6qxTHEgoqnQk+gwxq4BUEADvWM
qb2epr4RTeBaLE+UsCkj4KApWJS/Gc1RrdeKBF30A8G9uD9owQ3d9ZEc2jMOa9Iy0dIeOfcMqKFm
fNvy9hGDDQjK/tKwd5IT90tNC6Lrwqpz2WpGCZ+c9HrWFzNHF4+gcTDlj+NBZonm6RtjVsdkjD0j
Wl9BXJRPFfvD8+2k4HrWJkUy34P49JuVBjcHP93FdOn6oX7DNx/sIL+97D4KkvTUzTZ1F95JN5a6
A+l1S98wkDJjfdThxgdhP5MpGxrTz+nf9ogo20r3ipac75mg7olaEf2NDNdhXiJRxE+haxcDH1t0
4zhWzT2ldFx/irxO1Xk/s72g7B0Irq1K9slfBVADZwSjLWeg8eje0oxei9XqFmDuJ76bUf5OO7No
BMN71x+Xjz6aNbYObDXLOuIQGXe3bb9hMB4eA0iyU18UvkSVKuVNyWyIxu+KxfjzsMPNK9ML3FkH
G1gRtzKU0pPzYe8qt6MVFWAqFb4iFfLYMXf3EHot1cY+4oGWagXIZsuCwSLanEZJmBqCtZ4i6pl9
npJtHoeLbLFkO9WVJi7mUD0EGfp3jyViSie+k75N0VvD2ijP4lt50Lfs+0Pa/WlbRgF3Cbd6SrWR
j1wJqv/XdJbl8uSxkW0hjXEvpvl0LpGRgULV0tfZLaV16tcPmF0i1Qs1Nnh++QKWv0s0/Gw7d/Ag
RjNJ5XhpjpwWKUfIXYOnBVHwzT7H3I6ea7mSy5LhLTp1kSCIOVRF5l9ApJCrqQIGvFCSUHTFnHhd
GWbw4yYDQINTdHcMffgs+9/D+6n96WPcsr6cyzSEqWgAZsJozSVvtavaiptQ6BhbaI3dEMww0F3U
cZh+aontOnHfA1NNKfbJq5OCJOviKUhUdfrlsJbsk5tZzSShASBlodg4P132bifB+AaWTHj09eF2
GpFrkHRQzpHDF6FxeE1kVtCDXfINWs1Z0ZZ7wIVhKt4Cdx5It8V9dy8xKscPYC2GAqEGb3Kc5wO5
9a5OLtbbQowwOCKZ7DlhS1KbXETGEtH5wOVzoGCDxDPR4CIoXUsceC0g+HWyunxCaa+eaBvhNAbN
IOB4WcKe4aJxYIOsVvkAi6YMXjrqS84yBJHCVHw7eCRIw+C/qoaeCy+RNX/dMNQ7fbSTFbr1H7UI
XWnVZztdW9OSPBKJN+D2QmIiSPxXm4o5EYcMWACpmOxYKUB4bar8slIGu+hWnBpCPf1dmJWP9agQ
x58r+0BLoCsqDXJqrkyWBWR1Or2fNKPqGwicljU/9GrUsPrHVRWoKmXJMwggdHxtXkPD8FY0x36O
tUvLth06JuNP97s43BbL3DUtfaqMSMboYDTHCrQb0gWes571iDe7cGSMnSgZ1X1WQ358/j3uB1I4
2ug6WkBhdhoTNDwX5nwvt+l4zqHrrtyWb7U6EHWIJT2QO413HfNwDiXnLF9PzjbSpqixNdTliDiD
2yRaAm1lsIsdl5Hv9fcPAePPjxnf/YQH89fb2DUPmjJkTVGY98yBjN2XNzc6Lo7bSj3s+Eo3q9+b
axNSX0ivoiohM0MRnhj+dLr6nh1z44KEPq8ufJ/Tms4LQlL59lVZWbRyZuwpK2/UbpQ0hy/yTCJP
2e9H6ja/ywgyW1xCEYID3+FY+dHsusn9tWlM7tf0DqnymsWoz3cMu/G5aOYKXPAZ5IfO1tAjRPBG
fyFXI+bWSdOgtyhohKk5JfibfgukKbjRmMEjo4Yh8Ap0S+gIz3NbAlzN5zAkrCrle49AsxTFuL90
yRSsB7OnsL8IEBCoZDUJKbwrkzHic9Az1dGgPkWkU4HEe+HQUNApyBHPDemp9BT/F6e22MDk8CHP
7G11dFrp3Gl51I082GbjuiXrS6mzWo89iohLr0BUJ/WR+zTnlv4mwwsGb9YArngzTUuEsadnKOvs
T8s+5+lwNJjNjr6Crdljd8P4NXziSA9Lc/c7oRRe8X/ZSrYy587A5ClTt7tEIaPEb+ZRaG1zZKql
7P7VR8BQKiRmkt1094SEqbtMoYB62dLyiR5fAnGvpWKfe78RNOfgdEKdOvn5eoRh7uiqEqvF/VNs
koGCdyDCoIVToIQlL8X7kzBgt7eTiWzb7x5rDv8gco06unPRJ6bSV7QMM9xxouxLO+me/qNMocqz
EhOxR6ZBAzd0Uun98W1ZXTP7g47OvVg4vlqpa3gMkfQZ6SENPUryKkjOZhq+8bdYPimHddve4Gj+
F+Wypyo3fnfb3E5TfOKUbBE1E2UgO5C9sLu9E3Axc8LJO3eRQlQ2WXRQ5y5hQnF1GzEQlPc3SM7z
X+DacOpUfJHkAJwgOE4dc3kPxyhy4lfBMfJOLROEVOzwqagxmDyaS3ixFnXPbWJt06z1pXr578s/
9AdD/CHSOa1KJtUF/RDxKVgpd5FHU97r+S/3nTokGIfawpXj4qynvCkR/67jijEMKvlFF9iYnLdP
NpS+9eYMHD5uuBi+EEgmTMT80t3cCqp1+VWyDgB6gNqVbmZTIBi8J+HZPDKvsXWsALX3bjYzjCmq
ZUWW/pLMI+sqkVmD4Hd8aDSenD0QbhR0brAQxMPEg1/Tr/3V6XOj14SgZNZbgbP274aNcjFldcG9
LmkZu/H4Y+lNRO+2fQ5YBdZ5p767SZP7mPSzEAVM9YzTE5k4syZV/eYCz78ikOl0MXGTlrK1d2ZZ
+GMoWwlidjP/qCq3UzJwRjHNNFV4Y0CYHgupOdPTt+Uxf5E2I67SDKpK6JuE7T+BZ4oMRSYVMKnY
Lx/fY3cpplG+1G1L/i1X3pOk8x0ibxvZvNJEKG2qWFydHzI8s+fhtCUGBqq7P52/KZUkAkpmo7j8
c1fRCvLsXjUlff4RF7F7s6Gr6LOVmiNgsEtQvP5n5F9hsCAA+Iuf28xLr6+A7tooLZJScfxlffDG
RHQEQfDPbITC0GBNlkTg+4RKgOLqnc4bz6TUQY8mddnrZYCe6+A8lLxfqdZt0AKn51UmixiPPC8l
SpZrt7DFNzoGkyTGoTqMV8Wh3R4uZos75FJ/0iAZX7Zgkioxxspl9/xqANsiun+0kb1FOgELsBAD
nr9gk+xFcPMoK6uDZ5PUe8lkbxTWwtpqNsVTzS3sQ7SpWwaOIzwLtnfyfjmWInn2g6DiyRcQvSlT
m5SBWqJ1tciN84M7/S1UtLmgsm3BPZGFAdaTDQPRGyT0f8pd5iI9+mnb8Ez6ViiczruuNp31TEVx
tYj71gPzCuVNgD2Uj2P4B485V2qQ4zsst1ka6cLeiHTqTP39an1PXNwLmeF680plbPhotVJ4+12G
IloNBLEbFURN2EHU6AEN4ft9vdc2ooQIF+KoEuEW/2Ze6kz1uT5S5kbDmFWnMeO4Pg53AqFh8moZ
qAVnNAzlM0bMtJ0TPoHoC4QuJRJQMTi/Jq0A0RJaZ+10t9EqiFrSUanTCbX8opaAg4RLZel9V7Ul
SivbYeGA2uWSa8P22/oCxRMsft8x2hGV0xq7eWMzg0CFBCm6UQ2jRwyZzdSEIbV2FaSvQa2bpV60
B/zM0FYzIMBdq69LqdtyOyBwGC52eE+Mp2ChsVrz4Vi36neNa4M15sUcVySnQlPGxsGzB8XOjZlH
obbBBi4uITOCuH3JWt8hPGTEBL2CAe9BUirmONGcEXzLweD+B7iZLNkn7D6lYIcXr/EoSzK2Ox8z
wuDevId6fNGQK18O6LYUa3ANwh225HWvkwZiAoL4w2tWmyf5LoOJiDZULB/0mjjSZoaCTzFXYwGW
KXR/tLUCGNhUwQzC7rGFs+amUOeCUub22P3zmxn7RZ976UAe29oKAYB76K0nX6dHRTAlG7gUmvXx
oqOc4/XoNo7c64Ru8PO5HJaobEfrtMUMi5/y5LCTBlmkxAhZ0ezIOXY2qMJsIwmQW4jH49mLoSGk
OqGIYnxMLoyDNmYK14OvR/5/80292hqSrEJxb/+yOAKZnmEwPRPxTLWp5Z/at2Q+p0+SSUal/iru
Wk4+wuZ5aRWlTIOpqURLi85wxBfr4JNkk7JuPV213oxumKiSM15EhDwLN0eFseXfmgn3u19e2sqG
mksqkXLNZG5GJCNjtaSVa42VyCYU+kUmVQzuMq7ks3OPYrtclD0ttFKR79kRjMyKVfejXo6H7x+V
Va7QoafzpRDQnWRxOhNI5z1Ql/H/7GonG5rrWgFJ9zwm4BPfgSTjCL5bJ7xG+5KiR42fFPAvcOcD
Seh4QbGjdIVBk1Abz9lzduuelE2GRA4YhrJXnMqf8BqKuewVDsWNWCotlcIeQ4HQmcpgmrmtfSy7
Jk/TOsaWZSTAAR+wYchk1FrIFGMRSFkIjABBxpuNVL5KS5UZNy/Zfsp1wZgEG7FRBL9qOI0vf+K1
0dn1/u00R9CwUseqCBsvvhbl9iOuDRxaTRDuf43uKdfENSYKpYlHJlXmy52+3TaSEko1lNlOnzMS
+6imCCGF8tBdKOTHGk79HXPg7jNg9p0vDoQmPYtaH2uZOYeqXPuDPi/384qkpteRpKdL2ecvpNzA
HZoeCUrKIMpYgiIs729m9qnAqIMLnwWGSWCeEs25/lLwAUEROCs1/4yAYOBrzNTAQVQ7hD4eiSHx
2NGvr0TLeKgIdznOu5sFKBH925KlDz6/7KT7QbvG2+nJzpgOeY53uU3brOWNxDL5n1gH9Ihqi+f/
aY0gnvzJ4uoSJL6P0BQ20RNuIzWpLbLcJvaxp+3Xe4mjrOlW2srR7+FRsYgJ51zqkcwUIOc0XCau
7ZmwHbXt3N0lkl36QQcou4GXFPtPCuk772ooDowOZnh10t9HVDR5aGcwn8tnOpOK7wmqK3xHhYsX
53EcqV9mBwnflddSYG5zP1khVDQo0KLGRBWO9PW/M6Y01WvefTWDxDL3c7qM/Kyce0dMwH33LxcC
wIPoOd+8PHg+n7zWZc8z9AvMubpaiKbYf2UtLYWb7KzWp9V+oHwG76suGObKbWZLM7b5XVoIXols
mQCmN6qREaF1WACIS9LIyhlvfuGG7ADrPM0rqRk8igleX795SRBPn8lVK+jxXyTJRJB8wYLVlciQ
jVlpvpodPD6xgZFcSu5zR6fqynTo1eozn9iOIv7ZsT1CZ3E1Gpb1kf4t+Rt8B/iZD7+w4+bEUkK0
l2+GaXFKVkxR375We1rW9866QeY35UViaLAlPJGR7hE2qWkTUas7rC/t90u4jyOT09/YTv8nC5y9
FHhKEl6yPwii0DL/7ghUeMK4pJcvkgVTvVPIMkRsCxATQ8Xb7MAoaUlf1YAE2TTJrfouYxXY6OEj
1UGHAtbyJRkEPu6TWefpw1ge6+72U15K1XjMBBZAkd9ZyBR1qQKTO86cQBNYz2s6RHxyeE7f46X5
uQ2cBZW/rjK9vDX1cSisHP+SXMiCppr+7lLWF1t8nI3J6LOqDRN+ktDshu9lieBkoKdu4PXrpAH1
Ps17jsy6cIO3ZRWVefoinG73PY21/AnAlMUAGtQGVHmvAN4uOyk99kKwTylszfmD66qKddiwzipa
hYgKIkHJpGyfax4kSGtZVjre4ZfV7m5CtxmtPMDF6DXhkdRJpA9TY8hFrSSJgfgDyo8zpmbBdVBA
csHNzP5eT91KLD/fyvwR7JEPCDvb4Z+GWUHr2Q/vZPqauVIVGjxN03XHckEATW042CgTJ/P5sH8D
tXYbwroYBbsRJ7CUOagHRC2p5/IavOBmaXghwE+faC4rPrsDoeu3WjTHSaL1pPkWKSgY+DtscG2K
6LCU7joJDSjGUMIJBxeT93XcvnRbNpb8qr4P+8zJEf7QLX3JJx3oTloUvXgxrmQJoEfcvOKxE0u+
4jEzFJ7YIwYwXs8khsZM0Psgp0Q44ERs4mzk+TAGpYalg/AdjwoqxnW5OawzSHm9s8aNdZ3Ty53c
12phANagUcU3LoaR7CT7vIOA4ErxGL8g6Hor8teaDua4c4Txbun7PGOPuNkKNq/tgexlLXfrjN8k
NDfgJEUWzVizynNGel1y4o13Z/Krpgq9VTbG6e+LQQlqb76crKVVoBGIUcjzCqHP3eW0WBcu8ZH2
1s4RUEf2mxbyuV3pQltiMmisyIhfCAPSBMFjmaJGY1Z4zZrU6UuebJnr1lznjVAvZra5beuRD/m9
BX19IZyFq+nENHCz4vgVuKHRd+KC4OOVHT1DtnmCDHM2DmR+i6N07RRpm1zcxtjPqkhs25aXTVJh
OgxICPHpd5ARhjfc/onH2In6aRikrkH8CQB4sWeVQNAFk+Dwnhnpb1gFn46cHULMEyKRSIDRHRLG
6p8AwTHTbks0IjnBQmczj7A1u5OhgG26CIw1WmhiY/TvfAPB45UYb7DM8cIpEXfyGt1nQxffWmXY
82+BIIfaLWZ8KCbwOcG4M5Mtqa2tikWSgAZ/yHkTzbjIm3wcZG6jx7fUGZx0Hd9jLJ/FdYCM10mJ
h/C5my443pvrTiRixgTv0V1UJtxLgujRB5x08KP02xq8e6Vy744shdHmhkADqp2Q43JCAh6iyHg+
syDlu5vWok2+ioCs/yh3gEaeD06zYiRazKPUvnZR9DFuqrm1OpIiEoT6P1vxr8Uu5tX3i84QGECY
C+sgrER3v8J3dhUpNdkgpALGqpBiZqsa6vuRvtodkdVNcX4aejHN7t2oP1ikNFLDvmkKExeULvSm
ZJ10wjxFRw5gauoF/CyK6jKm+PV2RScfGlsCquCTav8MILqV9wYDcSPcl5qRz68xKcNz7MiLDWz1
vQMaxi+uTLpyBBwH6bbBFaJvUsnXgfChZ+zZlpILGWUk/YT5i/zmrPu3RornGcYHwak7VK4amWEh
vunXTfjbGmmLs96drcmEnZjVZg0zYtEgAoRzgG8njXNUf4ajunfCQ55R2hiTew37oEDvlPL//hFI
sbPKh/onFWFdLXEqWnJTUDoBmRP3oadBS5iHSqM6IeqKB8jgqneAjEf9wZT6/Di8tafl/wI5YdcU
diZGnUC6a0NYZaLdmyohGLww4Zikg4SuRzLaMqK9NLoFUOz7vhtz7g78Wx3fktHAMGV1DjsTjT10
ElJS7i7e3gmPTAD3dTY3bK/Z9i7VxsIvbdBjos7C5euHtPwCkNkSPD4IybPGDV8BuPUunsSGHRFu
5r1JimrH79T0Veen0QiN5SRmiZS9Y0P5M3X8ACuRlM4Cp52bc3/7DHpSpcQfi9qn1K1ivzjAMozE
TDt+o6E+cBlsjijK+Udd4z+qOq9uJmrypdEJciibfr9CBSp5kmcPsAB3nMFzkYwFH2sYJnU9/P7T
QdjPyYz3KMJRiXCTqof4sjhDYrPelySOB5KpbFp1yaRmBYXr1TA7OtUcDdnjoK3zSUysHRK9W5WH
zcKPfsTxyGOL2JA0h1zsv5f9mo8+xYK+FpEyM1qo1JCpZu163amdix0ozW4tUvuGnUHLVk0d9vZw
r6wfa2JP+bWANURNgxX4KzYATnvIF6pQ73Bk2ITAxHX32ZoM1eyv9Vmhfu0BDz190eGHj4AYCZRV
XoFokcHeXylk7aPxCp8v1dE378EOPPQ3kEmea3/UegMuNDS4IyjJ2Wz4cepdyLmAe3fw+n3ZrVrM
qCEZAJT9m8WIuagfr/GWoK67xTcfEFkUADqbmG3x84Mb7tXhQLFCL2oNjaD/6pKkxbwQXaUtmFSk
cf/VoUPHt4lwcRSqnnHEKw7lZEmTLSJoMEZ5wof4YW5E55XGTu+yKMtOxaYiinktPOqd9X56NrjU
Q/kaxnO5spmQz3POJceH8pCLX7wdUmwOjRjjrn71dZfXNtBPkMpJq22/3yMKZFaUIMSvd8zkg6Bd
fVSvRkPfxsH+YQtDysUI/Z28r2VVOVuHDj4GV9OJzv7JpywBYnoyW3sG3qFS66EwWJ+wm/BMBmLY
YWZw/BYLq2wI66sHwOix8/nuqn2dypumcepGY+098s5/ylYDFQd0GdTH6jnlp+J99sw3RKN6KDfh
x3QZQrhjDpX+lMLmG+ru8Xay4BJf9Q5re+L2GdgV8jpia0Q/CGltqFW5RO8KWrokmRFZCL0GKqLM
srKSF9ezDqjJb+PiLeo4sWbeg8B3ep6Csoj9J3w01WFjudSaozz1UzE7roLsT3Tc8E/zJFIYUM5N
pZ4ty7aaqsE0mhHHZV5zPYoDl+hRAtQr9yGtJI+pidCIjp7EqOVZW31o8frcPLokT/MfWU7j7jp7
hH+DhcioLL9FbhjhQxDTBPwweGsxbS4nuIXihQOEsPp8QCeyYTwtKVUCDIJyhjxTg2/rbcKRPh0H
eJse9Bx3gBqEJLfPdR0tdzzzP/gnjEESrBJe8L5x6bzQ8WMYKWZTHqPKyY0OAVSDtUfsR6/vWt7k
7rF95h4wp4H4W7iISDc88KNvfD+5wsgG0BgoeWw1Gp8QjNpeDm2TMAjwl0hh7/8gbS0GtjTmfiWv
YPgWwzjNGjpysXeRTKmhR19813sruXGh9iQKPk8eKfCPqUBRp4zWZixVKzNzVga8vIqkIVBYSgRb
LdDyqf4/o2WWOvurFMUlmhl+7DvSgcIZsGw3KZKUNwnW10fh0EevorWg7tQ3MGHQhLDMQ0/zZrNA
XhxM4sqQDGZtFBQgNE+MqXdIU0zkKJGNsfc6/2SDrsht/2kKbNp5fZWzfA7KXyY1MmAi5or9+dqz
gIETvT13YUdhh8zpwrosKZn53MBbh8uYv7+y2mxwOYnFdtTPDujT5dE4C3/FhbymnuNpAIGtz5pk
/ODLHxt+zOrDmfeiS4RkO2VXsYkq5V/7NOMsf5ZQ/CzDrsc2XQHDcxHrrePGxwRXVTKrXoBPrYsO
zjkQFV2Cwxbh5GtYNlaWjQS6u0u55DbimvI625uxkVJk6kvBPOCwU5yqp4+zahjOAU9oKESQo1aZ
Xxn9tM72z2qwE55M5fyMWTOGzBgbxKGgtJGZtN6bP+qSXMlCoWq79Se1J5sOTX815wXqU24ya2a4
RK/itHzkbHqK/6/deZlpLLP6RFQBgylmeiV2k0qlYRJo6p15tWCwrgH3eCPgB2ZcfVgOU9rQRHhT
WiK1LcBCm6b8dbU81d/E1vspMUYKFagdpok9dWU9vRwjalsMn5PMCHSb9KJOzxqQc2ejB/b+pgpj
ge+e0wvVqEgJ0jaEw+EVUYrnxII22fzcEdz5luXuqNs7KUEw7yitS5YgwxgiSvF6jTX2HpWYCJob
XngTMQAjbzrjzLTsOqSABzOoozHuz79mb87u0aKvojhTlIFDduT2jtNr5XO76epLoeg/FLp+OqPe
lPDfuhmy2W3/PdI0jEsd2dtJ0ZFqEU3vSErySzCtf/v69ob+zo16QJh9vQ+hUq/n9UvBid3flsJt
VSL2/CMZuicOgbyelkByTcf4nCAxXfIvDFP8cnhGeDVwUGYTryVKSeqIoYwfEQilQxxxosz/4fEm
oEsTYQ8Fc3qhEngfqy3pk9hxOu7HzKDS2lmgeU4AkqTH/OysJNHjaOevaEK3aOv6ICAGPer/UglE
JOXHL12ztKaOqyhixoiu7eLz6XDfInJSxQt2EWvnSrbyOzmcbxlO9uERd/auao4Ep72mSMFc5AQ0
oqy0eWAfmZ9Bfv6gfxhjgx8NdNZqYoi13V7xLbgz3yf97g6LyZ2C+e/flbkpReXAaOgNDJaMm5Ph
SwaTlyJEcn3t5ys1BmMbVsUmbso9Cc6VbmTOp10TNtCMLs+UlKV5UQaxx2J1pRPV9PgU3W8vmmPl
/kGDlFCeNZQJz3Lf7AG9nEx0km35KNO+AOXcdPNcg7cEGI4eSK956xhL/3AFwtB2S4w0mc0lMMHi
p0tyt4LhW5+Y+pddRbmRq49wCsraXMhZ2ljnBeHjdsH0OBOV2DA9SBMmlkVuMreanVDSBKPSwCRX
Gh5oRWIKLNXHEjQ0uxtww1t8Fj8Wm30IYPQPVg7runHSXUqfJnvE+RsNd47fvzSH1yK1s8DtKZq2
eU0HUqM3f118oC9XW0vvJWDPBbeovAo1A1JypO987pAHr5uPMsNuhulON5uPFOiNm4tgPtcozwAY
+yiyyAzAAWpfz6bdgD4jxMGSP8RTcE2vrIrcEhLoXH4CZC1ZNxQ4PIMHxkJGtFVr+7zDSRlzrwtD
g7TJVU16XmPvSs9Sl3s8c8DlvYWGUY6K56bMbsdl2Ag6JV1HSi3KMwcmcnPHhb8V/1obFNbArALm
87oh9QuFKmzDCwZ1BLLnICYO0+2ysXvREr8o4u7H561eEKQgk6odspksRK/soiT1bo4kzeYruiTq
7Dyy4m0zxeYMjvQVIN437XnxHklflkSgMpqJapEvK91uTCOETMUS07n0IBzIDBFZGMSR8xms1MZ0
0SUfqWzVHyh0Wexlak66OtFlxW9uy4BMOcpnKBjQ7/cz4npFbTXFPY++kTLBgCjXvUMe1msgrL3i
AeHSjWlzD9pGhnEKZ/L2vbyySv5JcHy8hMSzNi/v422xn9Md3NPagqqxx0ZTFQtfq/0tFvd2M4IX
Q6t6dYgCBaB8go+Lh0r1oYdarXX6U3S0gFQ97ucZIwNz/XpALsFzfs+02y1RvZOcVzQDG0ywLrZv
e+0y0/huOUTgWqbRRk3jTUbM8GHV/8KEddAaGX5NoUsk66UvHRj/1JD0b8N4irwDwsb0JdXqnquf
y2x7KvJlSMVaxjZ0FMWO+GzCLhaQZ0clyWv3tbAqjG7DgVPpDQ8dX+WzqEkmRvaAHRsWwtTk6f4z
/IBPZmyxvV86VDsFoaWpyNIVqhO37liHM3MH9/NGpieFtiFwzlLd9mEwh6ncqo9Ppn8DShpJmoi0
b1DrpnPmeiR2o1bnNmFvXeKerhl68isxG7SAL/GChEsn+CdJFoW3FAaeunEWNuCwezX5FZdg3cEk
JfwSDRtVX6vegrhHE7Yiy0DX+Kx6W9gdbwpYV5iLi2UloemO2vowuop83rQuhA6ImWbefYnzbhTT
v09ujdyrjLBbbQ24EaHEScanGxaPyxCxC4P3ORE6KedX6t3JpdrEUFoyiK6lDtJYSJzqtZq6Nk+5
i52Xrt84uX04gKO57TLwE7gFtH1IMV9iBrY9E7LrR0qWXGMgK4zmy76XlRsh6iL4+Xs9JSiK1bFc
3+yQtaej2AuQsHjvFIySnWwBu/ZzeZFfMrm6UmdQZFIzCdgquGzPnRP1dhj2L4fn2tTq3Hc/6kbO
YSP2FMXGrQ6awBMvanI+pVjQvuVuRM+ddK+mRJq4Rm4AbCTNAX45yHVVtmneS9gMi2o9fpX0Lz5X
o673oMvBUsxxeLk6ZxyV78+xZbIb2UGcURuX1bOtquOdTLOkVAPnX5ksHPm1CasP88wG9DMv8SI8
iHuFtOih63DM2dSlenHiq3rWyK2uWgFN5qtkIPp56PizBZtaikSFQePWLjjPYRPUg/V88VzHocwC
XmNjLvrllhmqzPc1ZiJUyEWk3GhY3y/ra7zt8z2P7SEGK09ImTpKRND/FRgoSK/UK7Fu+h7SUH7z
g1ARTjpJKHtgAdRTUxiWrhpmsFOuOwBpi1OfqoDpj4JiQnJn+k4eo0+ZyCq16IbMxl4BnL9TorHU
NaezLxB6rrv6TIwhV/YXHKUj8XNrRKkQ+dBs9/hbjagZJpd8fyPak7Y91mOmIzZPoC6gJGIgRKgy
nKgbm0eBdR2rlEd/DLmAF/VpIPfqM40g2Wl1v+VbNRQtiIBodctAN07RThqFJS/e/jrY69Pm+7nV
Q2oedakFNv/jHagRgnzxX1k3nscFFhTGEO8P88PDRywtN0GPh3sAiR4yqKlEpr+18Lz8Lc2BUlhH
Gu2+/hfLIDmOa3ni08Msi5PvZ2QcHfyZ3p3uzXgE5eH+iPsHtBkUsCUA1eXxJsSaK9Tp7dYE/cT4
HGbtgtvU4rTF5CGh4wIV4Rdsp9j5LjTSHoMLBYmhyXZj9Zw1R4mdVK3x9Hx4aBngy/8M44QwRaJh
05xQobdv0atCTo+2Y+yqD3I7ixpf46DVADjLNTA/bIdBFDHrx8Kr19BbngPOu/9eIXR6vhGhMv+U
gBYfjugYU2RgXgJLNGMV1pgxGxnZo83OGLlKzRB22+bTov6lLm4hdU9maFt18aFECJtSN654bkX9
f/ZQ5UQoJk8qWyTcYR4hshGqnFQsZaqw25tcBXqBY8WMxACTNvAg9YxQsp4Y+1kSVaJ6YO9lAa5a
FRm5jMLE82ktHr5/v0PEU5A+bU5Pb90JhFup35mA25nVRO1MUoUXg9cN8nVFh6hcjd4q46o3B2tq
2vs84wIh4wMX2/U4BdNxHzSJ1RDpgzdGM9MUItPMftIPkDoLgoBwpbgeM3UxESkxeRFOQAqjIjGD
QrU67PeDI7ILa3BByQ6/scVlw+YlmiSfT7G9cj6i3U7viM9dzMlMt5M948ovoMx040mG7Pc031NE
dJHtviuW5IzNc39Uq+zw3oj8c7Aj2UTQ7GUFJUFrVdF00wlUWXajq8A7k6bofwtixmRH+F4PjSlB
w0+jh2iPDadNptILBbdWYc2rsKP8P/CMvaVx/uwX+vdIyY4jJAnb1RvAR8/pb43UHPZ7Tj0PrOdM
QxgDqn4GJewePGQVHYO34ScD83tu31xQX6Z8YESs+2HqC4kq2cqOap46GFuJkjcq5rISDZ72RzCx
3KFGniwyap9pBvUQdKt2TQSNMajJ0N7Z+N7a9njG627+IYMxa49npic0KO06NTh4s8NiBfllJ/G2
4qrjXj42/N079pXgRyfHt4CEu8dYgvmxHSuRA3n8NreNXikpVPC0hxF2tB1O2ifZkYVri6g3MiAH
FrF9ukdTcGPFsItVcMgxeNCkfRZZ+MPM8k/NYw501RbVS1MivsGwUb8qWUBq67AzR2sBgC0nkb7B
KfSgqWS1S2YWSgW9hYe4AZ3maRmrRztyepXD6t/EhgEeDD5cW3RPULLJLKZ7G4gN6+1kzSuQ4Mr1
NPM6v7iD6VIhA07Pb1PuUsQeZCgZeCNkLgNMqgBiiRqlY37TslHYwZsCqeP4iXbQzF6Q34rj3lZ3
/PUcfq/9OPEeK7uQetD3e7AqgIgXxYL5+bbBYnob6i02z4if1xrxwfX9sIj6xZb7cVZms8wcXuTb
DRJuDThLt/USRZvUyHpKsPW4q7YXkrx29l0tObZxx/OPmk/ZNWjqrI04iBIdtY1gIw5pSHnMHHuQ
c1lVnR6wR5sUQ5HyL1FjXtY/uh5tTlTTS/CEXZ3FkaNpshn7adS/nBbixr8EpUtldBDdpRpw2BCR
PMz+eY5F0FUlgav5/qnvst7LJse0Gw8eLnQ4wVYAj6DDeWO2mnOVPbmJProoKN/eUmEyF2jRkD1F
RL2HIME6ldwiCe7oZ43SUuSQNwvFTPbwJu1LtSyMboTdx/VAOTb5yk1vv6c3eiIlSWVMr93bH71Y
kzL4WMX15wWLUxoglyVB1i+9gELcCYzKcOZXPTAVdV+9zXqhOckzDbNfY2y8GpQb1+ElIctc8aTU
gJ3XJmdcv2C63UmyrY0bcNJARXktvWqDXnjhiEod4miRfzTa86XnndN6bvUBeM00LmGZC7xnPZgA
eMCpnd1A9jAwQ4eUH42yutQYe3Bqt+KLW72Dz8CpApb7oE7p3+g6zn9iZ+C4H5XxtIobCt3dAzAB
NiIkctrggpxHaefuCKR5yCJsr6nvin5QOjHUXLNyuyo/8kieUTXYchixCmWx8uaAG82la/sXLZt7
/JsxKFttUVwSa/2uZIY8zNFbNNiXK02iN6FDpvn4gcAcg7Mc3XDxAfXW9m16SFoSRa7yohhsmADq
gVKiMtOo+jgmQjWDtPcsdZ0j2h+M4PRz9uakEQ8dKIFVJi2kyvdWau+0KzEB/qkfhsi1Kr/qCSUY
/O+rjJ9NVI5AfIJpqrtu5z13I0M3FvYVradGoi6d5OTEFlOYwURdiNsCwHI6kbgnDw6gyJi9uwBq
3KG7FH3GPFWPcHuda2mi2rjjbBfhpNuXtmF0MlDXccp62wEPgrYftqRkDVuBsSrPSah/jza9pwpu
SdiZuQ26by2w3mizTcC/ExFiEAhYPHdCScJqA2Wk4NxLmv/B7k6giyFFquJSx+ITG2aayw2EBLCy
MD6lzqakp8jG4ZpSLO71LoCmtS8v471Y1H1dwKZ5d/dswtd10XhopJ6EWK5mHl7CD+KPUAJhpaRV
itNJ9wQdAgTXVMRpllR41N2dXpo6gxFOHCUMIjKxL5O4LPlNZoDe5PyyMcQBr+6d0QGlfdgbN9mE
JitO25yYw0B7d1JIMJZE7VPskW4v0kFiD0bLJUh+jwM6VLrsxlnBllVVs4kPb9YA6kmgbFOjl5X3
2XxO7byjreVFFI9IK3FJ+h4H/g5epjd2Ny1D4MIOME/I64hOpNqBqCFB3KPD4aM5W/jiDFiylzw5
KBW/IEk1neQogugHdMZlFllIizpzVMPp4Q99SMV91lDRFuLJPJ9C49WjE5YZgEDQixgRWzrzERrV
RLrOoyDmcJ5aNjc3ZoNIIbbsQ5bSkN9WDeeeU5uTh4ld7lqUc7soWzuSd+rzpl+swgl9N2OC2+Yn
iZDB6+1qT+vXBSfHxQJul9ezx9xQe43sDvTiuXomEGPXJmGypHDt/IFej+5ys9DysibTJv5SckQ2
p6BSJuHt5vVOwb6Cn3t9WJ4jtJI+6QQDS1f1NUMSYZEa57fm6WVlGYhL2n8RAxB8Xtdg3XhVg6UA
hN/MW3eKlb7LlSU+oARY0d/B3tNijpGfAk1elsN9TTkT6yQhHFLfLIJSbMF0Rr+IwYlXD0tHkR82
Ki/lW7jWXT2AAbeqE7DtwSl3U+ic/7+aMHAzGpIrnKCd0qM/Jd+3/1gN/kk4D4GtCw/rtZvBkzXM
mzI/D0ySi+xju4bKRv6C5ua+uRPLjPqokKL4+bNKM2NMhzIFdfniiJKcSgn+j2d5PEn15wkSsnmu
n8j3nRt8u8JLeH3eTmT0SdWUfNvkkXr3pFoaOis3M67XbyAOLds95yqHueeurl8xuYkqbWYMa2CF
6HbJmk30o4AcchjZy/UD/Er1+VBtORjVgt6ENxNqAtWFOY6Ao8tgfMYumOlvcHHC6lkEqZVvwWx6
8ZqzgPNLK5Hs9JpnLTyXSQBa69F75Ox07U/gXsBV0nJww342JNfLl0Yu+dHgDJEPC5X+QOIbkx5e
dEIEaV/JJK9+2se/yzZ5UcDibHXyk5gqG5VnTMQnF6HSUrT+9iqGmT5E7Tt/4wHcG5jgsAFv7dtS
FldFUaqfzJSfY1ZNbvk52uNe73lPcYxOgFt3NpPPtOPVLf62g3CbpYyb08FcU2t9zIg9wFa96M/M
MvEHq8Ph4oMfxXU/gnJxryoaciEtMyWq3HplQ9JE1WwRDHSkO7jJ7axq44orfHP5YnKPgs8GHJn0
EsxLshT5wfOyc/eqbU71e2UdDvAXuPyQImdFmQRwY6+EQzkrQ3fJ7xk79nbGQg+qJW7xjFpakK+/
66dC8j4D6Q07rkvbNov65KVyYs7pRiLG7yVJnQh8pa8Di8XHXDhq2IYWzJcqIkrSUBbMjhhRhIvM
8FvU51goFWmzhc40I8Vkh4vQKnTY2aIkEOOFe6QUBStK/R4ZwNCuYNpoUMCPDQgvcs+067F2yOs0
CdnFrdriHAVLhqnCF3woyxZkvwhAV+bkf4Bmn7LEyjokrr1MeLddrZzz62luBOrH99wK0FCl8gYn
DUoSFR/8jfXFqdfbZHkw+Wm+wYSN9wcoW1ojlSwxdPFoIG+ljS3xEmP/8ALlwOoXgKKJJ72lMDb/
QWzRmwPu4Tk/mY2x3z3r9fTwI9ZIxD7lJ4O8/wK25FEBnuMBvvChOJKB5eBfZADFI/H2CfNi/JDs
oxCJ7Sl1fp0S9H8Fx0dZmwA7Hlvs+MnG/AELFiB4SuuOwbebkk79g9PwNMj/4am3SpkxKuS88oe0
cgISGe9Hf9x6ghVcViiGd5loX3na8JFXNHnHVpuJaV6b5k+rZ0PJd6HA9HVk77B2prsJUhLt4VPJ
kKBC8Otlz+USPm+v8fipiadsZ5cXxDXWIZ3uDXlT2pwgzHJ6QZXnGlnsgbAXZrqpoQmLdHJundyq
8nX6XKY1T566etfbA8IZHgYPDbS7cGllkVlPC99f7/nSp8sh6v50DaIwFWiyp1kYo9OXlwGBGq3D
gLSbE+VQ/druOsoOAA8n2khzlcZggIvn2eKT5cDOq1jvmM19zpbYaBPeAw58G9RNyvrGD8r2vlTB
RbCpO3XLnt238+PrqpTxFO5rAUhNiE6yQEgxQ7Rgf94DYzbh/3XNxnc0/KAPqYjYzQNNCxgDcGb5
GKaLEOkm88jAUj0HQDLZJ7ZAZglt/3w2lo2fXLBeWdMJ1UXIXuzBEGaYPiYI3l1RrI5sdDKTDdfG
FsU0utk0HVJTRJIh5jQH0KU1Ml1cHLYKJAB3y9GcYVy0blyMIDThjixoZIvDXsA2lieuVECCWZZk
GsatzyeM59NOVWB4h0zh5nF46zS/YcHU9QSRB/ahkHptaiDDPEMiaJqUmKq9bGATeU+CIscwYquU
JsTvui6Pid6QGdWgw/IJ54F3Ds21zs05rkm0atKWF29rAy/fxg5Klv2/yHpsWfmALlIeDPQ/S0yN
1zt50n85K3b8aQFZ0tGxokSgSAFwbchQQ/O4ogjAMUIwO1uCksAeRWJuIbsy/FaRF2kFMxTdKqZ0
dgL/pgULiv9W6uc1QmsESD8MObu5RmS8OIOza9us1EzX1TRWJkrz9+vnzEBgg9GIUH1YzQG1zJY5
cfXM1F+3qE96vOq19EMwcIGIo247sKRItSKLFlsoCWndlKEaQVp3u6N5kqy7tHzVs1vycdKxCfbw
HDosyAuq1F+5JvOqw64KIP4T/LO8X0HA9RK+MR5UG64DFLxsUat37wDr3+1jGLBwJ5+43nq/VDqu
2XUn2kQs6nz+wdOTYiF5D9NjmjmEbZorKF2cXZx8GECbqZAjXV75yHKOn+HiMst2f0J+NyD+wI9b
HDx/eEqoICjPFShiCDDBx8MRBoXSH/Na5pl+9rq6AAeVVow6Hn2O48a9/LSgoWBfiyxAYwalAzrr
CGN5sgcP8XdEOPmVXPoiMfyUAsBbXOICNl6Mue21S6MhxJd7jkYvqkItanokJvGXkZS2Gk0yDovS
+VEFc9LG1ZuNE9RLMKklzHwDnNaxK90QvSss1l/xr6LiufTC4DbfCwU3qntHGu3BNw9frI7bgeE9
Mtf8W2eu8m9X0/nfHkVJyLXfpCql7ABIxzFG8KcdqRJGmfXyyduh9U/Pi5Xf+JiinuDnmOM9w30Y
wdvAphgGRI1XaiyLyK1mAIBMjQg9DF53WPGSPrLfR9xMOafjzwOwUSQpU3WumpWxmR2+PDy+LbSp
cOsMk0/xLB6jK9PB6FIpIeKyPudaZDkeQZt1/8jI5bdS5MC6pPyU2Ybi3DQx75ZU/s0a7NDeISo5
T6wOVbbGpBiVqAQmGxe7js/6jaNngJPgbsVj7gPxZ0jy2FXfjXFZ9qB5FyrncsR0iy4BtmYR7xWf
peTeijmknlCh0PWHAZHApSs8OQ/RyxjoCXndBIsKOyKu0C9h10K6zkHo92wpGlAPTHHJKA3t/We5
Eud1lbydaTSw9BzEyMJJFWKpEqUJo7dm0NCblj/RhpUekGLnYyY+O+3wGxpX9zM8gChQm1Wsjc2K
55qE4MwwDvRV92G0KpFO6f/xlYqRNvRBc7bLxbiMpkK2Cv4g32ZpbexoHkMColqgIcnaOZv9/SWb
yuaAZ3iTybwedE1qClwoHyQY/TfYgqNjflzfvpR6YmSmiJZw3kA7/GwFS4vsy5gOyXdPhnZIux7c
Y4j5hamVO8VkcV5/rYx6UKu0KsaK8JxzmRJjEOv6PqehNRJbAgCSVNdep+WNaVpWgb0OTvfgSe9M
bRQPh5L/D3gvgCj1xGprstbpshmPDTrqA814NVsujggRbgVUArwYcQvZeCe2421rKwa2ezl36ZL3
Vllm35ihSB0zzz3IuAdlY9B+JquP5i8/t5o0gL61DDQLZA50ycC9zBn9qSTnlb3LJKzmxkjcHIQz
Mu+3HAlnLam2KrKOY1CZPsIFT9jUXRSBDQyu3Jp6972OIocmn2nLLxOA7uKe4zQckCC0yuKJaCUW
TTh9ia/8n9C+Th3UWcLhv4hyOFi/PkdsFkzY59UPWDKi4qkOA+GwG/hBhpY5FFkNckPmWKpdMa0x
iTjkfpw3qe8O20au9X3UaKq+4eT0AOGZSWZuDzWSqoNOVTLPQntuh991K/4KkMobmcPzc5dhmm8q
w2t0YesiMmt07G0Zq0kzEoNaGomEcyUEh+PfEKFHNMFBicHlsoVZrDoh4FmhW1yxyXhRqXQ7fF+C
N7Mi0xlwrmOitwi7q6/BPNzP5iJqGt/+L9tZyjtA3FOy3sQXaobdiWqUuAazN2lmWGUNQbiI6Gb3
DxU/3UpV0OdmqsQqrk8twSuEPUN+T08cZtdi5QGGbpm8OtRY1W8kQKEtL+kSz4U1wvDwUMa0EV0p
Gq+epHqaWTeV0Ruaf7SwSym3z7Kn0XBgT2x+m/2YW7uIPHj8cc1OugIU5nfQBaIC39Ffatmi6NsN
yByQYNVpmOGV3uZ1BRnfDahnn1pVe6EOq9fJnJ7ogisjzlmyAWT+EmfrugO4ApIw+rIWamjbWwpi
QzjUlJk5E3aIF8pa+01cM1nfL2fyZIA4VgnPm1LxMyHuAEdUXaw1trBZ91/BikAOSTd8Yfod3NOG
qymzJzJD9oNmf1BhgJUamE2YJOcDgnBB7EG15AT2/k4Ju+NV6Bv0m36hwtsonKiG+VM5q3CRYZ1O
k3C+B6kOHF2XNCp0qFP0q8acQpwytrMh6yRF8cB7GskmlZDyZOlMg2ghyl/i2Fl6ldBcscLQsquf
C4iNaShofJ51+IxdOqj/84mo+4F68Tm8D3e+sn/leWeknMzErWU/WKJWHEgjjNHqd208M2hlMrsr
u2zOnmcYwU4RmYEoC9fMfFM4dPMuBpXUtVSN0dKul51S0Q3fNqEGRvWLAJZ510jjNhYsIHqlrw4a
YlU0bXByZDCU5jY2Ss3XQ1dUYChZaDc0DEZS/k4aukxA9LmkbDVuWJvmXXvgrvPSQR9+Y7QizAQD
0uPeyRVEVMnLDh0BzNgNDsu90cAW/amXJ4K8ESc4PpLq7Uo8E60Jh8mKAwVCuTDwo80r3h53PmIE
rHHkqWcJ6Zq4Y0NMAOJ7EQdUSuADb9QJhwuVfBpjpC6fWkc0QzaSfIDsLExG3ntyGfS3ofMVjuKT
H0pcoy7t2eS6htl5RUxD8p8ozqBPcFF4j2pp/uDX/hMZnPt2c8w3tzDDTvZWkSW8xfFJKS0RHqVF
Rk3KQccHv9ZhG/Lv8X8b7NrVTKwHjZGGYI1O1AZTAFmK8wN/B0b4GKxuLuMwWbn8LuhRtxk6clKL
vAeWjhl2WR4aK/wp+EvMrFoXIMtd54Jdf/9R9Kzy5ncv4L3egaj2KlAEU4wynhQIFX/haKKawvvY
eTTPDUm7GjtHsLwGiDJ0No6A+sUhbRsJJxnltFS+zvrtFrxsTXnBcY/g9yzTPWr6pXawuZvGxYlR
uKN/gZCM53vRWxNJ1JQS6Ui7Bl6om5GYRs5hOiGm12x5LxD+4qcW6f2ChNHwjMycOVnLAhL6MmP1
mmIHdFGAUkwA8tY1pG3cDRPfhTcXr4Tuw+u23RqfxrwLabeIBpT/xJGwllxK0qKyXcT2aMSTiV3P
vhsoWlIvvYjimbjxim67FotjVrCfsvimZyblLJ2Io7NZZSQyPsisb1cpdGoQXBx7liQmhbAxfefa
/44T68vuLShxulcL5w+vN+EQJ25kQGodj2xG2yxcXe4tzf3IwAnzjVJ1zr5SxgRdATkWSVzchu0u
5UzX+mqLrZCC5i7HdQgYZEd96lpz/2hL3T4uNa9m+uujQCi7UfnqXQqxG0ievTeBgC1EE9L812NN
ciVZk6m1uZbkm4U4aUOnc6TuVq/QVX8FqtHYOIVUlo3/Vmsps2mpy0q5zQVctOPU9w8YR+aQ+baT
WPAwt6jCbv3gnDgrBfsNJ6HLVllJ4/9CdawLrKlXhV4je1EfpHDbIsblcdBrybUk38WPWquZNfiV
RW/dzdZZnp4qSO69xvkel1ReX+h2K6ObsHT/yeDMAyzwen3AjljuPrmTNy80oZAL3/CdfJkH6hNH
zy3CETSjMhyrh2Dcln+DW0v3eeQomZx353yUC62EIAKzh8cZrL2dmgQbUdnJ6ZUOn6bPIKYlyele
7uEpWIQpqC3Hd6hMibPdLt5EVJo4JdWHtmo7DACCsEhkG3QoGLFIPLLw69MLOAaRCNZoCy9Phom/
a4tcuxtwQUXu/MEAxyUSaNwBRb2Ru4gTBQCrsP0rKkTtyxnqrQ+qY3wYToWH+50fWBFoC4gjGCeq
ZJiTKQgko7GFgUTByfjCNZmWXRcgfXeJDS6tXvkQmGgfXBHspljraC4hYmD58//GZiZzhOPtuX2Z
t3TGeokGhctynMsS2pRkJ0mdRiJWmOPIH4a2FtsiswZONeB+k2lhULGJYTKiXYYWdiHWcE4vNb1r
F0TQ/3ksZ5NjPIuSj1PPVndj+e3V6VcuIkcw/NNeCJUVtO+nbZyjeGUDO8Lfo1cPqp4rl3yIBI50
l75znIyN/8v6Hm0GYVnY2NH1SOxdXq2Vn9LSm9ldnq4dZIX0Eo6nN24C5XarjgtTjNEdefCyow0i
IVUkENNRPeodKWF49fEZR9NmoJHx+MWLPSQiFbsn+j+TaPIUnIenAQ184EllaUZjDHKIjEqlEQuc
jV+MfTyd3HN9Wj28JR2zEHx54b7+iH5J/aZipymD5nAhLWjSEMHBeCpLKLjRicRM8V/7cIJVpynn
v1jh5kSJEqm/aWDMOJl02d73qWq1rgYJJGQOpf1PwovW7eX05ANyCNihpUOlRfdLlQLw7Jl5QuTP
R4HFkmYykQqBbmPj9BUgb3HN9uC/PFaGVM1ukt6GPxWLCTxr7Pdox+HEDcqfYORnKeM+Ej4iGtx7
RVnH7B2B4Fv4tC3kTie/LyLhLn6mccOaT5//fLM/5qj7qWuAtxV+fgaXdmuZRS35ApGV+qNIGULy
nRoMRhAnFj+ZCmZnT2ZLiVbdG6Le0nU2vgZd4E9/CswyR7+CnUx1BP5MyptI9F9Qy0wnvfyXgeGQ
tWXZVVzt+G8M4vhmQU7DIK6KciZ2KNvOHBTvMxVN7Y4agZoxbrl2tcJtd/a6muUZwKCdLIfEQqou
Pew1vesZcMkT+uk80oemsGf7w/MpAbkDWofh8MaCox0zAJ9UEiDifLi1uOZ+l5pCKioAzZitCrvu
ab2HY2HrttYjyo/vCoE6Xrv2XsViRx2IQpY6f896ZyiXuNLbtpdv0OC40rTd6p3DdvQZ1Vbx2sMO
czkTuDjWb3QFzBaqNQ9zA4a9f7ER7VuOEKZNtxzWsHfdDbc3T8D2l2Z4SaYMGYfgb4S5eL0KVcar
UlBdn1Pbw+7ixjkKXG2mrDT7D6FXT8bdAEFjyOolrr/iJjutLUhgyzYsbrSqx2UdhfS4oj/IuIzs
9DaELvuZHWhPfuL94e0gXQorZiJlVQEIHXdxyiWfy//k+RLFDmpQCZDaSVF3LRhiPyFYWFdmndfw
X/JyJFsQ7CUYEcFnPVAZdYHmZqjEWgcwDGL8USvqcB2quGexGFFoDVdOy+O7cS08c7ZozcSDXfL+
UxNKRsDLLNgPGvoMizk52FjKPYrL5X1bo+MI5V9wWYe+lliHe96MsKu49z+GG1je3wUIizwl9Ius
cf3LP1FwpNAJTN9Th8r0Rhl7sVpj8v5dbQ5t1xUqXog+XO08fvgEwGnsLmZPZHmaN3bADDgV7au0
+JpCShXh+GQTY6X/cQRv//GZbsBVRb0aktxiCOg9DEaz+cyoJ4ddYgow0dPuB0pA5RSuBs1qXiUZ
NpHzsIqRM6yJ3+Y1HtBeDbub3Fe0enphBCyC541YcV4/qvo0bqoZ6GIp4yNhQGtAF/o29840mCp0
RBRqPx8aZrRvyApJ97NVIN3x5yWcFGLhfOvSHCO7ORe2qjfiI24HtyybXA747gLKuvywtwfeSMy+
dXbwG9pn7iDt8+alBAcuRiFXxta1hPzrq1GC4ERx9IYJc7o0DdS3F5GQ4Hw03T70vR4z8gAhB22D
zbCkQZypixbze22pc/41xjGD7PG149iyoOytzyErhWICtFIcE4iZS7h3HStUx0DL512pwNE8sCKC
UfYPsa0znQY7JeNd+M6JOtocuXuj85rvZ7uZcpJWZDkJaE52zRPoFESruqT8y19iwqR1Chyk/r9A
0+IgAilPsbI9uEPu8KFdqS0evFBNJG1L5b8gfNIbQ2ShDVK4l3yLPc1SS8x3HzAEcHII8qlHKpui
JxcFXzhfd5y4pa6ykjUuOq/C68QjaBT9cp0hTpEWUKTqVli3isajRnxeD3GDE+ecEXzU/u7o6UMo
CJxSWgV/daSIM34LwGZgAC96e1WL2p/vp547lIjIJlMzsuC1pNdxHA1EQJ4D/Ks39bU9gXGWnzuc
iGuJSR0p9gdvtiQnF3hGjZR3YkzIuPs00Q1BfiPwP2nSKnDUDagPWLkeVJkVUgX/O6xzA44uflYx
A31FWK/njm/AV6j9/wRhK+8vR/NuoO9PgJS5SJQzhrO6PWeBImY/jSNLi1RVJjcMK2qqUrjbslLd
BNrL7fLvrS+2jcEuIu5BtUMP5Lylb7YS5vPd/0WXmIZJnmWEwqJ7Fsgk6nTQV6eOtAljTG5eFUEb
RV4ogA+m4GQPZaThD6wIUlkJd6vbvEGAUF62J6lkpa1fzo/Xke+7RXrUgmXUB46AQT/yV/YbdLDD
8Qv5EI/XEVGMl3N61+VcJ5rMaD4Cz0tw7U/z6DdQBkGgx9j/+zaWBuRlxdRUYGpfE6FsIhoeH/co
VFMzvmTGtgo8v+wUTUqPzfkwg3QBh0uO+HG8ux85o7/dpoJPyljVkFBR8xcnCD2N9LK5RMsy/Ope
yXOdjbr+e4pnja1B04qun3wuWbeoHnDK4U2MfcnWBNtVtWMX/A+D+wn2XpnlIDkeTSdTjdk+v9mF
FAlwZDhKVcor1mvUEpvLoHx/1xFkGpr//kj/yW9abQdjbo7hm4ms2JLJ61mWl/h7CA/4TU6nmdP5
HikoSFNR/GC4rcW1ol8kqoBerp6CfJ/oCJBQnbeg8mZ0y+yQIYGeZDxx3/Y0bCsy1y7/Epy+EXBi
8cmVYueQosQ17CKV31RqC1/WeR/m0VBT7FbICSAIjoPcQGbN7t/I2Mm9VMwltbA0LMa6qHEzM2cb
08IojMokBMWrsSJwHcGR4yU/AbV0d2ABEguKxFED+Gwuw5t2Ba9DE7SWdTzxQj3rII6dAl8KNGMu
j49Dysqqy3clsmTWGeZ30FnqU3PBKwBmI2P/Iyarx+Gx+68YFfmOvHjitHdCM/OWbO8Ar6tk3RxH
mGcCYubpizp9p7BhFfSQpTHFqKJmNWlXW349s0FIAdeA3GkAr5aZWohLZk/0rEWSMYTqBS5cJW1U
P5kdGUixetBOb5oC0BdbhtuO6520eHYNYM/rcTIkYaSpL7XhcBDZuuWKzRMlxDQjsVoFjigDsqe0
x3bVIK6B0/9lHHzo6A2D+rslcVaMfjRsDYHrjZGGlTXzJCupk6dFO7vKuc85MK07jCNQoCr70DF0
iYxDREKsdHRF9AmDH15i4+jq2dFWawueVWRuyJPr7OdT5L/UOEC5MCv/MKmHzUuYMSD2o497mhIM
HLyQW28skAecYASSjswfzrNyxewsjq47rtzMcBOk8wTFPqeV2CAx72zgPpA2Is/k3Bc2JMCxRmZD
Ww3cmAeJ5vLjdS95bwZEXkPEtdKa1pGKLJAOmu8PszKP6HNJO2PA4b4GPCR/RC/9OvQovCRtZXTT
iGhXKI9X/+//f1+5KwtOvhdJlFRivy1uRfD0+b0MBRyKBcyDaqkSwAYDQReJs9ntkEMS2QJQRQhC
89DlPOshJovTxgi8XuCNkc7E8ryg6OyPan0dEQcuHgvSfDmNAKbwhlOVXZGvNCLYjkHb/DYW5CoA
RhwddrcFOpKA9wACvnR+Cn2lEBncAVKq++FnBT5SvCGMdvFbnvCRVT0VBQ3mzHkJ7KQByL1f+rId
aV9ztA/gP+42hkDrHyR66kYGTUcE9ahRhwBuZ/lB+jwNuf70C0akPfP3Qmx9dhLtMUlWpajGqB3T
NHKF+601cYu8QST8WZK0h5lTSe2Xm9Y8t0XntarCmGZVcV8v4FY4ry5TrYkMv/h9TuyjLd5qEdVd
XO93l+3TDiHvn9tZax5hLHdunjAC3sNSHc/XBpZ8E/PCBpHXvug+mpOczwspG+kBuXnsQ/tjhBAo
WHrYniUuztamgKwtSNdcCpu8XLShipdBKBvGvq7x2BJC6Gjp8sd//HgyifkjKEHgGPbvlmCVwpIf
KyM/eQSx9Dn6+KFJMGfs6F+fbKHf3K/hGQmGxZY7zUVzg8pllQ/6dTZpgTcEXV6dzc42pDggjclV
ooOcbqUcdkC6WORUqhqRPrULBtnk+RTfgDBkA32Z/VGU6EcQAfK1hNDj2SYs/jU4CrFz8v+xYAku
6RxwZ0u2wKCeKacIiT127p4ea179/vkprSNc6BrUl0cD2GOcbS72TAuEfuwSrrcn2kFWFrVSrOVP
3d7/86kuyFYnFtYX8m6D+ki2aCE08JOchWe2WuoFrEC9wkoKLQHjggxNq1zkuv9tilV8tna4GcZb
TB42A1UQMGXyN+50uDhQ2Rl/dz8wEQvnqEnC9DTkrOHULfy3PCtsTw0JGfI8SaByeGDPzL7vFvmL
M8xmTSBPNK/w10YFGrEbBkognNjkolgKPwLrD7ZRjB+zGLpZvF1peosCNOG3tMi32drdqpaaEBUy
gU8djDP3vvlwg5S2wre2WHObI/JhnK+xGbVy+QkwiyXbbI9Z56xfMZfLEWyALbdgZbPhGZ6sHKml
ch5rVU0u1q39gYUp0ciqlZz9pQQD1EoqzrelHsZD+AGFLAJiLhTGxmes5yV85a3578piKFf9p7jA
1n6xAecxUswbTht6EJAwKunxkTnEOovboOGB/pNIW60gEwlvpPDwDQt231iUtyC4th8/lZ60IMMl
IAUQ4IjuGyhY5P5iPQL63ZxdvsYqYhM8cW3+ycLHNSoWmGEQxBmHApPN28IxG2jY8Ri376wZ2rPt
PqNTLoghxVRqxk/ekf5UtRWO954Xm7in/HbMngMYAP9UaqssC6Ts5NNGXHpVYROSuxZSKqoZ1x0q
KEHH+yN38uGXfeW4IpHcdQvxquopKwisdXIvl9lSC+KGK7nv1bF50bGSZPGPkH87W5daqaqZkIb1
fkDGvnZeZTByvSJ2+prtMSmDcTRdnYL4E5zWtX+SdU3XXNAn1VNh9icNgk2COGrUDIHmaURwI4om
IDcAxBUq6y5PFk+SEUKXcZn8ttlh3QtMSFWGefttYV8nLoEUQ1KThCLgB719CmDoiC409O25QnMD
Kz3gou1kUzQFV4CITeHpy8uNzgkRARchAc/vJeo33G2IlmRPqh/C29SGW2HttIEcf053iV/nUAve
Xdg+IVL4oyRv2CJD0MWBydx6b8ijk+nfA+9PfEW+s7+WpL4yq4hv5CHEiPw5euYPLtJmZu8TgbeO
GE8SZNnsW/AX+F4oxTQehpk1WVDXcwl08YOdYdV2PhUsfr2iBZk4eZSfStn+btAfC4gVOeb7woat
WxW86fSmzjjyFnDc6HysCYC9hyX0Yv9/iO/II6lB7AJVNMukw5kQBT+39eBWbF/dYiZvN74uEWoJ
J4jonaxAx2BDuU8nVDI0juQeGLtcgypOk0w+U3d+lieqHFN7JJFzn8LcxJjraie/HlpBUI4NTs2S
D24PvxICRE118c/fXIbhTCNg7wTivBjdqzVHyNqBfJhCOpPE+96zkK2J0bKjx87Oo4Rt7DkzuUlV
w/3dXnNgQUj93Xy/wyhX0dCLQK5BIvMf3EUnNYmjFjU6y9SX48BMcGs1LYCzq2395Q4z0o1vpA5V
0FS+/HtiezfJ0+zx32Z5lvfxlxxpfgjM3kSrzGxnBgl8w6GeEhADczKm7NnkbCQBmHLmQ3tI0fJA
JmLcPJJXrRhcJ7/PwAigHaGXYUwIYQlzv5eyjqTXQrwx3QcrXhojVSOn4GPDgHKKsO2mwmtwdufq
ZPOlrVTigQehtOxrBzRxbOuhg7kD3mXP3wIoOBusaG9xEXW18stobUnCEJzXhNrm/A9CzPPjtC0N
E4OZ0B/dR7u8RxB2CEwXVPnLAVApH1pwBP5RrFZPIlD+eqpREPkZXkYZQJg2Y5euDFidnYaNQ+nd
5B+Z3YJhK7h4REONSzF0qWRMOJEReK3MDx5bDBgu790c1x4I7Qa01hwGDtwndcuIeWMrKBqtDkt7
XjHhVJYE+g/quS0rqn5oK+sNuwmkrXNGfcyiRPjh0xFTGKDt64TH3NtJdSXcJRR8+EtB6QsdYnuY
TlEfu+g3E/mAgTQUdzdkX0U0//fZKTX0W4/n5x5RDixxLWBiEvIJUBEjM0QXQURzHySyYsk22Y4s
mJPW1Wl5cGfUcuuqPUelEYIUiuz5ydVD4PgqR2BusiuTv7FSzswxrCtfJpfndUikLhMhCWJdOAn1
Pw1+zLeF+waJ5JqtqdNpIlsXj4aYEtFtqiMoI7xbz3DtoKUA5uJdoD5oZImFt+KT98cZyZTd6ZAK
9Z5qmUeQ/Ecxnil1ATcGGbGSrUA6jPwqvNwjhBCzZ/hc81Ba1SN4GTECmSg8eGHXsKKylR0qYBff
X/dfI/cgGOYVby+jDtvWgSqGMt+OUiJrOtcX1Cy5baJKdua2oVvAx63EbQn5StmAMLE6KIFQy78g
JnOoyRPwPED8zn6D8/R4FAo9vY2f0Ut8jsif4tgzigi9pHx2GxmFt8xNYEAgnP/gwdd/oU3Xs8nc
RAWCHBEn+U0ORbzCXUacIn+eXUQKqBnGvXBQWYnXyahkCJ5FM8/UZzIb7HFdYddDfCe1igj1WZS6
sl47nwYpsCt/kCktz7av/1l4fw6rle6uJJX1eFMuUJhfd8m9vU3GDP0Bj/j6gHljU0iSO+RZVBqh
DLg8UmCpdaAyuxM5g3OIQCgk3i5Wmo1kf9rBGcCFs0z8MQtQifNonnZfp+GyMK5duRjIVLsvh/ts
o5YhtG5kGgtlXBRPFsSvNECgBBdVokqBYe1aYBa/MVLznWXeq4R9clTuLzl84dk02VjGPKdTLt+C
h7njNvTVy/l2Uqloqv7X1dmyRpk2OZlXPxSpo+DXyof2M243LTJCpHvGOX6x2D23jn82sVVz5oqr
BtMHqSvu+2RqYkj1cwGPulatnUSInRf0WeM1kpodYxvFkajhiy15eTjBqaZ5iI8DyqOZ5JFP5sai
jNgZOYrmh1ZNXkkdHv3SF0VwvDBgq8/BGmbs0AJBfHijNZljEDdLkEXBE4nImlS9llNXRCnmubK3
5sjsswPbcfdTW5f4k+uWs3665Xu0cRhi0g038deqoxqaSEn+g29zrUapSRD6K9lYvbc2NS/ROcjt
0FjoBy+y1bw5PWUnrQHHL84QiAQXRhc/MZ/dnsuqB7AwGaO4Uck8C+sM3+5ZXSf7zFlytVglkwZ7
23Q4gQtpQACQXJZM0w3l0VxmUA44vxM/RxwSdMfjptM3iVXBlFflkUgqkxG8HXBEU9zyeK7TXcp2
AsYOT9cfaMHdsa/YfPXxzBTSVaC+UVsKhDrBiRzG2R/0sNREr4cYO8QEmR58XElgUzjPMux/UFVh
LzH0vmr3BMUiG1U2h++LHhiuV0Q4LquSbonVbNLIxrbhJ8qaNTXV/aIM+tN94yvo22wNsFQ3jSPo
zKOoSTrDMPYnn+DxrARaVVamiGX/O5CyWykipMErSaqdcPVF0JIpLJ5mVjyIINmZIa2tiummxtBj
BPUFDXCmMLRU9JlCVQ/jXUXI/hGETmV/pqNzfIPF+R3k61vO2mAOgLeJAQ7mUF7mwupGICbr2Xy1
tXyDKO7Y2dIf4Xrfk4fLn+jYBIb2OE5wFiyrFm1L8ZSdf3mO88PtoC3w6SDUKvzvkmWbXaNd2luy
WniaiiffXr6xNevU67/QSyL5EITdpk2IbFdV6AizYC4SaY2rz7TPXb2cOc6LOYa/Xp21eGt8JaxF
lNgox3bD8eAgAKgyYE61rrGBHhnuFB0Y1q0R/2AoE8/Sgw5R/fIXRMW1tB16EXTjiQceJzgDAEro
HxrRJeMTQAk/poYSnzhYfRDKu82BfAk91xs7uuKk3WueqoMvByen9cgq21sSQ1rfcytfRLIxFpHc
KTkl/QcdHoovnueSWVH24UgYlQr4kQJg1kEtVlVy3GMnH8wE6+hDwgIO7Whd/GfxSubKR0MFmSLX
ENixIO6QAMUYSOqH+XusMaUw3tmdSITyu7h5B8ZsX5+lrACtNqXiSLQCYb956qWblhkJkXKCWgz6
HrDNqGqOYgscOuLjR7wF6X5OWPvSYxmJil1aCB7tg9DXrwY7yvWDKMOkEjN8Wsqqy1qpf/ERv9lg
TSxm/ke8lcwh5y0rtA2H3S0h5XxWvwxcT9o47Rj+V/8cizVwrfGpqJYrrywhi0Ud4Gj5JIw2d61w
za6JnEs+7v6vq5ad54Y+OFDCO+YVp+yivaSozjn4rHr3evpYvEFxHvlY8I3dsxZKKef/jRP5HmK/
TmLzRzSXZBZQgcRlW/donr7NfrQJYZFK0G4WXGerV1g2LdfyZcsbfcu58ZNqPs3Yj5gDP1kke+Yq
Kv7p+1Z35sVsE0Fy3IHsN0ebJSyB4mSjZ26Gaz/VxI3PpXMBDyisBh4pLCnZnD1GV4XyoVrev9gS
1md3N2cMO6lya0HssRZojaGOINOyhG6lxSxcqxNUtbBREEoMsP16QMvoFb+iEYB0W9C8o/X2qTwX
e5JVsiKEx890D1e72oypxmmi3CSndMoqai6EfaZRe5wMuiOI8fgQeqvyNnSkMO0a/pYXKSCpXeA9
Sreaqw7bAaUEejwXkoHeQFvaUlMX7nSWfum5Uj1NKECmjGadq4+OZahY/RI7WxKAfPDSYoT6S2Xp
9stpnQPPJx/83dcs9b7wp4b4YA/Qn2FztE/K7IAuM0MgNuzWzXtXsl8NVeT6Zw59hmcbks5Jef+p
LFCK93ZLw49+sRgjE0v/tl1xvhjilf1SmNgoLkq6F4TnW4OxHqTNxwx6Dyg20OTILwe8UAqzeUGP
TQ85XnIf2Qaf+4B2iyGvcpyXxjNfhkZsBDUOdu+1JUGlFOAa7WALZPMiHFVNMS1GpO07xfg85k6g
1zu9QKn+nj5irZ/ONN/lr/N9wivwIc4QAPnSyOJ7A3+uwgGmbzT5DNcDBvLwEl23uW2OEl+7wOgo
XwzBEEDr7uSS/QQiswStHyqfXg/VDq+Y+FjzCNm++MWVnJfGwjvoWr36i4Q0dAA5I+kT0jXhy05K
2cVNqrFKx7xndAdDN77IRe2eXwd4h5Pzp3iKsIHpHtvvW/QkJM+EuYG6bd6vLZHb2fn47HL1GLS0
8MeMOD3p/fdmbyK16qkG1U3vIRRnEz4U06rSjMowkW5RN3JuWQcQxzH8CfUGsORCF1tUqV0LIY5A
H3ZNaOZlITHEtWEeD7ZAJAVmEjjV/AoLtXLJ7GgHxyhwzs3QEGCkkyZg8PJ6svirvMnaITW5iyzq
hqiNkTiSDtxNTnEfULdN5NWSWNMvA/GFVvnAtaNFio3dllY/hrhmd1RyySm93j3xQYH5Fc7WrAs4
ayesToWI9qlMwH8KzFSrCww+RNhBW7SClfNCeTI432iakb9SnHxiH+j5frsrGpND3/VEE2O9AFZ8
pb2ydXj0QBbQIKTgBAYaH3AMcILQLqMkF6N0P0YLTCeuglrFqdP5AfjGB8MMHHu257rWtSl1yPUi
f0DzmifJQg0/LWyGX5P4KwDjpeaGdonOT5g8i7F1EG/iDQyC4++Hg8JUDLOrrxN665Dh6xTLbCnf
UsxwLL2rT7JKenK9mPIfahkqRV6Ed+vcXL2taxRioAN/DUDha6lB6qZ9J48CUG69HsH8mgt4Ps5q
++xeTKK2Ggo0z7pjE3KoDogGk7LIpznooaMNlRNGZx2SApY9MGKyK9RRDJ861ZjB8GI5I/HPezmk
9tpFH5VedBRyTmCRNInun/4ARZ3mmOg7GBEzjteRjHWX6cLwsr91WpFQ9JCs7Wyc8NK0MxZGZoJc
s6vuyNeImoXFzOA8JnM9N0vCf24N2o/c1fvuQjWXW0RoHSeJ1OiDFC0tFucTFcXAqQXKdF0/OQyO
kiMEEigY9wmMi0flVrTCoU/j/RxeALT3HMqbuYJPht716R5ZPj5AS7rngABxtt5/29B4AnYIPUFK
5pY/1oSVsqgztjp3yN21D6sNp5V+7z+YtCkZOS+ZVllH5yEZOJW4ge/Uzq2nTHiPTzqTnjO9XWiU
mmHmAeLRgzM8AH5skocY/6ofgC4ep4CZ5te6jVhlLeQ39WPFUaPUN/zJYHYLEA1WvBCol/ZQ9nuu
8Hsv1kM5vXFgJBf8rZ7usM7XA8XHMz5CSg5N3/aKxRmWVVjbT463ul0qlcsZKAojxqOWyAjA07I1
bduMIWoJ8f9LbwWOz/du5i925n1WbLmOrt7+l41AwXRMTcPiqLiRec25LIUYvnjRN/ey0WusJPLQ
RwTAqEdmeajqKTGEJNzH3jWYIPiQ1yYCm1Qaz6gHG46YJdOXkju82HHiePG3WMS52DDheRxr1fZX
u11JHBO/LoQAIY/0U9WiHuqyiMdXCYXtt99ndQbUJfPGDXA0tp9pFsE2e2yN5P5hWfka+hHspSHz
dGzScyZ3ygBSxabQyfm86kU//+D9F0UJx4G4XZwYdLli5BNbyDurawK8vcjf2Tnnz3oy88kYRtar
g0xIdk7rQibB2oP/FOyclsq1AbhFV/U8Nr/HVpKb6azgF4gaBkILhkkem6zEKVSIJ0yyxRxhWLJ7
l1K/BiDFbLI1xHu2E3Z0Zi7uhMFQ0ZBz4zLjIwEK1nyCxyQ7CrcUTglQhIPQFMnyoujxS55wlwT/
lpB0Md67J+bs6v84adClDRgZT59gak93y5ugQlKqUUdw5P/CfuBrScKd+SONzktw3Updxy5IW06X
t06/7hRkMAEUHiIioCBowdxfHLiYZ+pzmK469HxhHhXJcQhmnEjSb9TR4hglK54WGrYtiOGiGntg
5Zk2It82a8ADSdEg5SqDqIoak53v8TOBJHveskUzz9vuaGZi+rPUnZaMSokaay/GWbWiI43ysvt/
vq0oeK8VnrsWfSrGPDy0UsbcvKC8YR1xVxGv6PPIeJKGHT2F1VdAPktQnjw4i4zSi+EXJ2xzWDba
DC5hPXMfQ5giz3Fz1l/nICi1Rpyff8FpWH2OuQ74mfUENtLaDpij4RodjAMum4kvafiZ+bWwo2aU
NuBVNyrQhD3q0MNFbBjHSe2PISJ9K+6SbWiS/TmNqV0yavl1XioA6DdUkAVvFboXIdXnbMZW/Eug
ugsethi/05Cqdt5tqtv6RGlCnZUU/lOw3WgNqTMc1ADnIxVWez0RVVhIvJ8NBLmg6Y8lQGMUYCIc
xRTf3KH83tqWWGqw4jssDm0TKN3LWOoDBmZzYS2RXlUdAduCGIT7XH0PP2nTZPb5GNV6CTc3Qvht
ZtQWxPYGQH316AWo60zZim17KYVSYliOVJu0HUKq5x9OQ7UHNuuAcymWbn8m5GzlNOG1aJQaUb7s
ULg86KIgsO5/P60BUZrbQY3a+5Poi1a3mQysE7R5FeaNqsJGYMTWXjkQT7b3VR2YdJ47YZ69ex1C
tFXx9Dw11COm/wO2c3uCx/E+lqKqUmgKpU8+n+yOCKPvtjrIjCG5r2VsYB+ZcMFyHChnJ2Aliant
S4rBNvole+vujbOOyz12FkeuByljyKaXUjEvc+41FXz/F35yVQtLo+x6pyOnIUwIE3WrG1qtX7zF
zc3Yms9ZRBBnxCqLGbZWL5kLXlbz1ajZPTKbhpH3tFg01TbiKpW38MBmKiSjDkRSh/fwvE8xPdgs
xLwRxbqhDTd2UkzlT0p3mc0c3NP6Cz6biRmhxNvYwhZrJIAXaAVWux9PiLjmPUIREi/D//ycHrt1
GBMmQoyM8Sr9UlPijUGO8ShafDl3Ww3F+WFYy0ePCo1bbzwH5d4o8ynKX3CBr+qsHAv6x0BB66IW
FlCMA3ruqCgcIF5nD/fZKKqmuhw7XrKvXNFPlQBVvEaqrC24SRTYwjrH1fxWCVW2XSBse+4Ceu07
al8b7mepNhUYw/Ki7ZVdjztV2ELxwWalkLH5WO1wCeg4K+ipHnv4k/5D3i+YW72LSgVXUo1qIKqn
DzwGaE3q+VrJDv5h2onXOcxvsza7gEqFRLVmFtdDoDP6v32PZEIY4ailw+jvbqAk8ZZRvL5tZi1s
WNvGHvlum9z/xlZasFVyPqUuLKET52LTKAHh6DtGiqlj9EvMYHrE5e5ownWtl9Z0FFAAhYsDn5Eo
YmwFFBM0rIiIEA7lnzh7gwUDBOD6OHEOVSKfojfuCfmmGxjvWB3TFQ5oo79GaDAE5uUB4Kk7aNEt
of5aeJAqezwW0TdTLwb9gHNPwaplgPjKxJdKwp8qzGJoSKSW0X99r8tZHG2IuPrRpQeYywtKisxr
jMlDZltqAVy7GJJL53laRa+OSE5z9XFW/hrRI3m8xnSL3nm2jYeP0xAreGjzciTpAj9okF7g06/x
KSaHzjTl6amVUKGiSU80qsLO4QnpWlalQsEK+N+5BiZbpJQhG23SjreZSq436WsOIo7lPXi9OptE
imBl3W+795q9McpOPPHRVwND5cJN9+4zWqf1QvY4GCASVr/T39PBZbNcqHcVJQJkBT+8ozgOP8WW
kQgCDFf6vKrks8V6E5SCd/nXJIhFKZjU5byQbKXNYyp1CEqs4hp1rtRGLE5LwG4oIfL5cimCfcAT
5xymukYsDxV8Stj28bD2ipERrd4wb60AwktfzosJsVcZKXQynWZ+Jsi3/cmTNgpEtW7bUyw00GC4
FA/lEbFgswNTVzu3oHx7x636gEdLdTN/lps2lB4yfLdpd+zWX+EcWp0YEnNaeZP3cj2nAXH9E1Bu
Haj4rGvjlYdMtcW44Ez7gvUYyJTH2aH8AZtvoQXC5TnprVMWHr6O35VdY6asVUJ8TasW4wRT90im
gGKApaxyhYL8ywcvuNeqQopP0xFgm+Ka4YKtOZcConTRVNBVV4zSyeKy1Kye1YxltiBdJmZ6El21
lgIdc+m928tMT3UkI6h5cVuGgtAxZrcwaN0EI5xb0wTb3H+Ip7T6BAxUn2pa/o8ArdF4bnDI39Al
VT9K6ewKzoSJdacoNwVcf+QBKme7t9pXV1WnxjrzpoUItef08w9naFfoEk96hzNgWDHyc9ag6+DA
kQb1kxlN2S+ljYauFAXxhD2H1YPo4R83hJX+i8OUXeqYEJyAbhKxAf5aZoSI5Q94E8cgNIWJCS5k
AdzI6kNnjjugDUuHAVIHhiZn98bw7R+/XxTYX3PZxZKONnAPdwMsEJ8t1Q+LSpz79oP3Yp321+YZ
xgNqfUudfmKhFGLv+2wegpol3G1AaHoDpdjllu++y85nY8hrLzSjYmkijAa4NC27vtazHi2+bJl9
dnAK9rOWzHRN0YtdNzc9bIjpJ/xlAxoF1kIzQjS25hr+1bUgP0Oj/wF79qyDxZI/q8DHdrTbrMiF
u5nlocusDUQPv62NGxJiwTmPY6h36/npanCXUuQvicpkejn/gk0cWVsnz5AkdSyUcra01lPFHB/U
GC28dVqJQ6/U0sIt5Le3+INlbadHMQb4C7idxNl1lJyTx9QWpjZErvP/d60rYZL3metP89u374BY
CPL3xRznioFXNFfwYZfYu/gU92Uxc4pRghQcdA0A1phIXUu8SEYu+oB+g1C6tLZd6G9rNiKtsUR1
Ze3h+bz+ljvXLNpG5IUqu8wAB/QCzvpHqK2suQ/37MKpwgDUCJCoxA9lCPasaBhW4OP28Rc/wl1X
Sj3pE4FYjI6MSrhGv4TT0BrD0oc3B36H05tVbTtfK1WBGtOHTVQOuxnrWuOmcSyjn2xrDYB52KLP
kUo3QHcgL4TscwYzhZkcQpZ2oZ4ZiwVzAL7m46s6nTse+ccQdbeWolphL2wcJyJC5DHFKG6Gfskb
PzBx6jEt6Z1v6ZALqQsPZr8iKCSUjLRK32LbeGVy2lX+9XIg2Ak3PHVG56sERp33nQWDyDGV16Nm
dgrs0IDVjkOWHHZD4d+xIXiV+Y/7Q2paeGav9Xui9KXyNkk8hpPejG674SmMPdxFHtJb39CJVTqW
ui4XpJIAJ8SHWBKwl1xEG7R5PrrIIvXdVmHN7A+cwXC/N0Tp03Do6f38lcRJdxWtqvzm6JPFsQxC
zkcGZkhSFHrvKxHjcixBVtLYflx8ZzMYGhvHTelCjnUMrSfGJUbvwsPD6U0Oi77QOMtvguNet4L/
t68v5As4w/DK3ciKvQO68FxnVLPGwCfCNUuyAC6qwhn/F3KOBvQYwmLkjEqHwvcsHuT+PDA9qHmA
gFIAk2gv9ebmyD0WCqY+J3Zgaj8ci/Tyib/+RVzA/asSnOzRMSC5OkVR8a3VLG4epIGHnYHJQ08v
Pt405qiNOPBfsd7KSuj7Q56/LRuJjEY5+Fl3FcccSQiBXeW+KACodwJ3NuA4AL/FnOOZtBoylNNY
Mm5KKp4ABhqXvVJxz0MZe3/F7o/GKQTV3qoPeyJRKKKdrpEBD9nWy6MRpUvoXW/sT25ke9gu7tC3
nIFD1oSyRLFQVxoU+ZU5s4QHHpK9mBS6Agb9OWvjKyA291XoaAf4P9ksz8k6Pgve1D6LY9Z75eao
rw21CTDUuSlMf3ExmnrUW0UxkgHSfFYdl3EIEi+9DeihqiWYrlyYmNCA/2A/iutl244eGo+CgehY
X/fNf0ghc9JbB6XKcs4kvP0HTOScy7a3vm6hlXGltdZkhGlbOpzxKJCKo3ajXfUWETrv0hQgZZKZ
mVf+cfof08eD7eIf9UsH6a3X2BZtWOewVM6TwbGQHa9bm27NUZw3ZcopgMgGiN2cwt6P0rZAv1l+
sA3DKBGzHnIkzmkN967prgqetNcx6JpBF+TZVwlxSgzYMROojhHQqcAimqqhfBq7s+fKk2yqH3Au
QR3OrebINULjiY4LyT8C/9GfA817iOOaL0lDAhdzmGPLe1ODoEr9SymnrPtDujMKeExYCttE/Ffe
1b+oZ1hYQJplvTdQ4h0k3wt55ie3XZsVtjLnQgZfze7wEJHXurQPx90imGa9UTA9oqQeri2e/kSl
9PDTbw3p6kPYQ8Ka9brM1tUEeAL2O2CShgmFZ7XnlsohHS7DX/PF0wi5YPTPuFQnJVMBasZJU3AM
2NOoBEWuP0OJfup+eQRwPEuHgi8pJPJ4RKLMP6v5hOVHGM45MYI4UNKT7AjC7SWAS+Ry08LoFXlg
ps67L+DZe7PHbYmq5NO6/WdwSxxpqNSsMaATwId019c8F++HbbjrchXwlbUr5Dq4Ark9IBcUNfd4
bahvya5YqjIH+46G4j10NXhtOKdV3HXuF20RY48TnTq+NXcYY8bKgeCs32TtLPs1d0lS/RvxRlRp
biapxQIRyYqBcAyHkgS34566F5QaS+5/DyIWMXgKjr5vEeRGs35T08s40txZKSec6wqdpuUAx491
5z6lzsGmh8gqesvnHvHcGNiFYOLauQN9JRddHRUa0HAj8sQ1/qNsE5kDn753i9PP4rYC/JSwZP8r
BN3slBKrzGEfZVENWXMAODjOPtFnE3J8BxPrqWnlkpI2Zh8Q6mxMhxVSOt0x+BStw0z2U69rKHYy
LXpMB7Kev3BiALA9UNPogHcryqR4VHhY8MIeEK6dBrObDHBuKln63YLCsji053RbF+I+G9UNnQ3W
OwjzQ84EzUEt8n3PAFW4WCTut6k6nHzbUfV/kCiCQXOz9+neUdt0HsuCvx3azx1i7vtREOOqrTUv
o/wBEJnC7pUwENe3sdw8z5Vc7WIsVb/ODCWnu3OLhQJs6xPoRZIdS+4FIeplRpbgT0ohtQlzVtgt
IMDctgxhOqiiB2sGbl2ancSuRVNHwL1GGXie0wpYkLq9zJJRW056mBIG/qxhIQ47e/Px7lUCOTTe
SW/XiWHnK/bgag/f4BIQPIJtT5k18oNxKoIkwNvtHV9q1LIcMpL6nPHAUNH5BYivb4b+Gm6shd2/
YoA+M1QswkiCgcA6Hw6nQxD+C8c1QwIB8Z34VKlAZDgszA0lgVDUsrmpqr5fAS1Jdkvav2Lp1Ufe
1u9RMIxuPPK7YwbCzPPPqahthzaLbaQfbZ6y4XKjgcEcw1WcfnNDhP5hirNVfUQ3JUCG8yoHryvt
6PXTIqKQMKZYUGArmOFYzO4xD6NKWyxCTv0gkgxNmxgsHTWlAhIZGJ6ZKsc3UXRiNjs+gmACQrkG
DR2y2m+EfWf219rGANictuTdc7+cVvo0jx45s8/RJShZiu9gMBBWdArLbqRwrs14xl+l1izxVq2J
K05k/tX5ltJiOJZ3y0l3O8muyLd3ZT8A0idZGomdiwSNjocTjO2g804YzMNBbc0Xa+N9DEVqAEoF
2I+YNGB0e3q7/I6MsYGgtRoujhP0NbUweNZwjyZgbfsuqHYf1RyosmR3Ck+tYz8j7P+4lFml5cqW
6JQBkRnqBeCvp+KvSurHin1+c87Mg8giyCb0MrakG4DGV4nsNuuGV1ua+Gy3KSDEKCC1OIRBilSI
sHvGr0HNmZZDL/GDNpQdQysr8CUjjwXUw4VOpXfJuTdRnUNAKDFx4ksEEY5NUvbjIACYtlLAtcsa
Q+ej4LYHfdjukQiGUHun7+jF1LbzVZfShe2cEqw4vgPJ8pNBqLOvAVSEgGmnR78rJhmpooYbzO5Y
6bpALmBDrb8jiNc41TBAs660Pc1rKNDgtAnz1IjZAx4FhgPRIomAvskgDEtAIzsC/x/CXCFFHYdt
pTV5T/ZGJ/VormwdVkqbegiQjKB8o4z0mN6vGnyoWWp+HIT3kV1+Je4xzcufH8sqiQ5LoM4nCosE
PtpMvZeWPgQVr/lSCtl78u4GgOAyTR1aBwfFia78vEqdcJd9xx9ZKyql008EuPMdcMsFevnrs/eZ
koOJgYFN+dv0gmb5zOMEeHKGLYC+jnfow5Q9CK18w8JUxzeuXMq86n40FwvoqZJIcFqOq0Czy+lH
6NJHGS/7no4myzo1muatZJdD/r3im56ykdTpE9kDhhQ5LAISYaIVj+AW9ehi+Drr229UQcUWRCx0
4s2Xl3EI+MO6Jx3sREVHNYtF75AccpclW81Bbj7QK8Ac7QWboMzhr01UpWA8DVNndITqoUTP3kwb
RwUq+nAdf3hMdmV9jJ/WJxAUhtpiJdFGoKzK7xBhYy39O6RzDDel4Z5IUFig4CjnRVa7GaIzYKr/
sGHcAoFvKNlxLWCipKF5En6e3/ac/vBTeYdsVHCcsiHryebcbehIDiyFa70z0MzN2heQuJC1r2Vv
lUC48vowzRqa0G2rWCRCW48G30zHEbDE5EDaUphXpX2vrN5okGcE/4nuqt+Xd1Tu1jsFbYELq0mp
0HE3hA+/B1fp87ZA8dgUuVimN+DWponaCCbh9UXyEf/bLSe4Ox7D7/iA/1NrLktWHQKwod+0KjDo
On3da1bL2HYbZwe4qANy6y3OqTckXOsJKpr3VvnX50SmKbzQnJ03/+wRHgEw6dVv2fwRV5hAM+Zp
+9+ME2i8asGK85ll93HyLS1CbfxfYoo2pjFft3Zh2+8eSV7AP34iecHjoYQfzGYC9TZC6rIMeBqa
UQF/zqzJUH0dBrDXS8SFOEDL/A/jwOjEWEjA5jZuXx4buX/Va7cLfVwm8IsQeQ+NDjnDI4kfRW3G
26qKuWkvPTx/F2O5rHTAh1FjVQTnPCajYNfEiXP1l+CPCLUZrGoZaALvtU8H3u3ljoDYcelPfTwk
VsdlCqUW2JVjPwGZNHP3GLZg5HtWSwY5PFBRkPR4VQkiYeUQOTxvqO9v4mhU3bccxrTkZa9LAOsi
AtDR9BH9DgfEBSoAZCyzgHQEcEg5tvqR5F3CyoA+0VQuAyGbpCn4Ln2GyMvrcz40LbeOjGFFNVwi
so/3EfAXqST2OA0XjEBMc/h7MQ0SLn6p5L+ZBHbOd68TNAjyrlBiNf+jB47yWk+5ytusAnXFyKFI
Z0NnQXgi2/xLKAUZDNhxnak7hZUvQHFMEg016v6bLhsQ2WhEB313FQN4lYoxhcOq2ARQXW+AR++f
P1lrH50kfkL6W0i6xKZpQ+sJ+qwLTTKZcf12u9+ELy1CfvZ1qYkjYxxi4MdW9bS9by/ZePv32UI+
RJ3XSuMvy30hOTGrrPCbNz+/bBcHgdA3odCHbxkJHmxjJzCejPSAd+ZgayAGona5TFTC6V07OagK
6GEe9bUiLaQfN0YgkO0w/Fgb5IMlhjttCoSKcW6hoiZgaaz7jnRFxpVzpQDDgX1HfXKHGlWy9uQe
/TFDiVXaxX8pk/MyY3Xx2FpaQ9cCmsgcj7zgkLxc+7SBsZQZyRo2aS9cW5sYKOzIAOqipOmoFUa4
X5yWE4kMYeFKqt1PzPcbOHqPw4/Gir9vMA6rREhxt8iok6ol4KLFTnCbpr8xbfj0aiBS/So0lqpF
dgEg5qFcLCO45vJN41o1rAGhkrBRfA/lU0eZNRoK257xXoZ6ZnkQbtthbReMsLwRLV3YPHe2IPbT
FmU+/uKrPEuajmcKyaNKEl57I55AWp3USxISEmgnQ8WML11q97bEqgOUHMXihUorQC41P4K+4vJR
J+f0CgwNSOVsHEuxWv4aHgrjxVVx5dB6Qqjpa9/ywCgSQM1qTt/6d3mYZaTnk69BPN9teKQ7sdH/
GNpkOEXrcFbapGt9kmXsaIzvJvJ04j7YNwk2r36G38Jd/yYRg3ANEUZZxRIm9VcG+5tP8kpQw1L0
FRy/bIaWE6nAuSY9RHI1DnWdIPR+TQ+NgWgSQpkILhhSPph9GjA0LCXzqwB3GUUx0gCNKqmlDyC7
JP59rXymaRGl/34P6bu2A2xMieEWc+A+f0q98faAYesQ/87XEd65mnJSlBlJercz0nnzOPMDrXv2
Q5n+KfK5jjhj5ZPwUiUNrrWWNl0cQKehiOzdI57jJV859W0V+Au/CcitBG/Tnwkl/KM2TUPcGD8h
zWjwpvbPbLCzH3+8MvlpBT6bFbITYlvUgkT3qLwJxrJadEkD0pdwESpBIgmnq9hr68eRmrgR+Oie
PtS0WkBFe+PL91boDT9NdeSsi375gvTlupW4r65E18fTLJ7/k9NskAfW+BEcYEotKOKEcFl+4MAY
xgWrkcGnoO2dviAUeHcZ+m/7kVN/Q1ZNTrJX+wUk3fHkak718ZSlmS1vpfBrs0RvnRIy54d/ngUM
ZC6n2OViPnFCZj0D2kKC67KPsOTfZx+O6dC9m35oy0K9zw3w5+Iz2n66zQzAVhiVHHeFwkJOoC13
5edSNSawqFlQxferyc2NYiGbOURMdUoM1h1KCA1GpVFIKRjAbRhEMyMK9tQqLehKNE2dOqGm6gwd
bwzAShmG7Dtx1dREzBk1e94Cwn3WBI0710x7hfqVWw1opwo+cc3TDiqWmwimqQxmgmSB6TaKkXlm
lVl4KWgLGVV4NusUyqLBdEPi5YyYl6kuhvjn5gXHiE92kkhzIuomA/5WY9vKQLDKvU88Gxhg1HfK
NzfptgAJFNDejqv7saD6R9xZ8n40HZcJdyvNVd8Ru4fSYpJSd1xHOiuiXzTUiW9mcEIiE+Kce/13
PQHSYMafwHIRxcVR9b5RkQNWzy7ISX1Xne3KDkIpJrvUHweibojnXmiMLGdaXDUetEO25G9v8l7n
euM4PnblSBdBmvfZxzMZypdbgKgTFeajWnF3pcm99PhXDEP5CogDD8tgmzAomJMizB3F27MgfdSK
PMWotWDke1VzUT+UB5MlYNETnY9nrsr9OgP+E08zELhnvkRf2eHF4TTrIUh5sIAgKG2aZ7oNbEpf
gQ5j36fulWOxwSAOjc6WG5Ay2GxlqakPr9mISbGQm6IiDf36G4JcU+QxPvHbzSOtKPvoeGDyO1g7
ZD2VU0JTmVP8NgzDuM3zYGmgOE2BVVPn0nyBN0Ncv7Rz6JAe+n4Wm0yw/kXr0wudMfeIkDiELYPR
OZ3tvpCoO9VbXWDbKG/JIaf1NlRn8+v0w4H3OTKiZrbs+fnN33TdSpVrqdiFZ/2oSleXy16Bmnkf
H7uxTR9GA2p6ovuYKgATPtJnpVYgy2GPAPZO7/4NpN9sx8vKKWfctGeVWOaKWw+BX5mg5XRG4u4o
luSy2AXYBw3ZGx4TYswwLmEt/VZERzTafVwvLTo1R/qm5UfwYpGjpTu4j8DQwkZqeQE6jw039WHo
d1gYm7gcXEdaERkBWov/sBPJ3pMt+b3QJH19JQh9GYvYDLNWdYsMZQ6QDe2ak+NmEYl0a9Bj93o+
g200825H06n9SJmT0/22grEUbYvJpjQQPFMVv4R56c81TuWlrVXbqyS/pwz0MNi+B5ATgxu5kf8X
atIpo3D1XltGBypPGlqiIO0wrKi/lq3nu9s4DrnrRDLi83aAb8ul3G2rRAv4iOTewK8GvrfVGfjU
g7cakK2SLgReI7MP36Ak1EDuW5dYBHbFrQhCNYKeVFP9IjuurZ104Napdwd4EqByYYsZIBY9srCo
r5KrKhXuR38wB1UvFdxtHYXnYDXz6TpYsiigdqBfMYfc1Xod4aOWWJAwvJgMjWnuwmCWipPxw545
6p8kJP7AmqwUo8kLt7lrkgz5cgBLoVE7B0I59rKfuU+aj/GIELftBxNitjSn0Smkjdp8ZqtwAkrP
rur6mQ2jMBrYLMnutBVlBN/y6Ec00HI92BzQSOO+JEpUZOc2pZ0zC4fczRFzZ+l4ofsQF22Sn+gm
iZyx2LyFSeQPKcYvSQJMcCbkUxYdh+qXZNXE4zRCVxNSSJUjv/nKAMGZOiPo2HlQgDRQgacL1DX6
EqzjED1PIuIJ0uLNRQPJaYjEET2qCUZPP5hJyzPccXMcalFJxz2UmK6BNzsmnROPK6g61NsNMQdg
PqkGHe6Zv12v1GLYMILXohl4ZnJjlu0RQHyC/2aZ/V80CJFGEPAgiMBGazrTlqpF/DyCCVwXTHV7
QJrVIEMnRfNK3Rpn+EVoNhOJ/RkYrC2ymeYeOkADE+jEjha/+vhKEdzfPVxmlcQQxwnzTpdi/rOx
M2e2MJkc+1BErVg8oj+WeOc/YfryJWZ+Zh0sK8QprTo9RqAJsOYVhA+WHpu/g1DNLEioexIPfRru
WLvOEE5b+zPvAO9CqHW0OXKMlhERmWBPCB5lljslxcHHETJHRSgL6D4sKnWrUe8w3PTpnAz5NXZv
At7GpShRTsD7rTOY2sL91CLtY5vac0SyJ2oGITinz3Rx/ULlWaQka01jfimz8o6GproXMBhs0Fp4
A75oXhiWMx3GYgs1oPmgis3zDOMlqLDf252HFpoBdqk+WWS6yYxVwObvJchJTz1k3D+hd++LZGwL
dAplCjlQBJLWj1js2YCcqU/MCtklFcMR7LH9tcT92mNCBFBewE8malI+dJUnattQyZiWyfmjErAu
C6zPu/jndQHNOX8pCUhTjOt14tz4SmmkKsIjBUS/FdwW/edY0XP5tFS/NlzBXDI32lJglnRPOnhQ
b1uVVJQhF3vdM2DJ4ZXgCLfrO4ZHR8/xh0+DV/Cq1hxA0smAVgKlL3D9ETT+uBjPdU6StjMvMAv3
uub8N4EjQNvaj75+ZaiO1Ax055q96Q9CiQyGI+1f0ufwOwjuCoZXpvc+atEKvCu3lR8KqE1ThLS+
41T/zKbC82SHq3Cod29zb17ZussNzF6UdbCKdtsQftiKompnT73O0p7VKwg1ZHy8LcEq3EreUHsf
P73iCce+YGNArJUD/h57nNAg8R69J2ViPzYvQjmZH4Kl59L1XKdiEgFcP2xnOwJ/d6HhqYsPmzWY
531ULl2MwcJOqhmY6HH0MkkoxtdO1Nvgj/b742/8qx4Q3/UPrHA91epcRlk08BFdLjdHx0hQyP+D
/8e35VpDeGI28gYnCAlgFkzkvTRo0r6l9nVDVUx4Mzek1TFq7tZh+eO77povsEEp0gcBurQvqlF9
5iXiOjThzByf+qL7wmNXvpRKTG7M/vFOBthV+bRlhHSLpIXGEWAPZZwU1qI30vGNqhBUcP7JICJV
4bTSvjBs28h1fLPSwpsFavQvepTWM0VvmbowgGUcqI2bd1oy+R3MGgHoi/hFUfZo6moEd/v3D9i0
a8EP83M2xcRldTtIFH9eU7EUKxXBeKDbvhHYLB9zu3pw1BUYbGstcFoZODyY/7WD0fQyzhDoUVTB
YCoqZmYR/QU+Up1yj6XTY1YfPjEgDedENud7nKv9AsGafika0aTupZSk0Z2cs+dZ+lVfwRtkwS3M
4hD7ENdAuEhUwvI7BgGLIOqLo/vq/2Yypuv/FwW9lK275X13ZayOxo0cmUw0P7GnpKdY3fuZ+SwL
qBfevXz4PcaqFqOyKr4SPnPyegyYoHzZxlHUe7WGNInnAKtr0DxP4JmQssWiIv71DE9tsrgrAWYS
v7o9iK8mCKdD61Tffs6MijQ2UovJj0NTUIl8/bFcc+olgQ3czMbqxi1BsjtEe9hS3QX69ukbho04
gvAzPjNpCvEQmIn97AdYBLQbb/6e2EgbOR4a7NkgsUUuqpHEpH3zPO6zuc2FLtaG18PsRDyA4tEa
xFnsK4ZUZoSWR9PwakYwSRIGFF3LotE+h2QNB/MJoDR7zSvtdTwf8uCtZuup8df9SnuVtxjAzgl8
B6nbGA8JRmfxRptNVBaUyY/hkUirmlRU37HI0K0X3nduZSRyXdyOk+aEX9wY5UxNmOE97/oi+QHf
oLcm1HrtMPKANJB8YRePM+gt6oQK9HHpQUfK6pDgCw4/yUBwIiiJilaD+wNyySGRD24JHKkTbtfC
ZGNhvHndDfwovIF5XHwfKCcgIVVn6QbfpIcvdglS65Bd2Ad2z5dg8m9zCd3fR45Jp6d9QIrJKDWL
l9h08G0wrTAwDvlUEZaeVkK6Pda9Z36BxgWq7sKZB5GYKVNBkddB1jT9C/gfmEUnwuOhBdWPwtQq
Y8vCjs5kEYegbtqaNlSIBQ38lB2I5dH02Ht9tcJAk5evBX/S3XMRkm9jThRJr1CTtPWL92BiNUiz
38JECppGWMgIKJzaqH2fJz1MHy7Ah1vvheduIeswlxLIpafwxLDjCrY3ckKLaiwH0zJnY91iZNZ9
2JbCe0a7nTHfEIMOMYnDTXrD24sGdiDYh7zr7IGPbn8jMoihPSLDMeHNdHx4KkRugue+UK1KWlKo
kFAkjYmsEMnvkYSS6IrWSvdrL/1zF/Dfas90GzHFtfBQZXJ7dJaJy6kb7YXcVDNBJHUBC+WKQzMB
OXXQJRDrf5o4NQCuXnDP24jOX/wHLM9G2e0p43iVcHJP4543jNwBDkOqykaHkPayudHu1h3C8UIZ
RStNiP30rQAhYbiCQzMk+FwGbZSLK+DUj4liS1Wc9RAE4k4/wGxUn65VSN+HRF4VKpC0OMmMgy1K
SzZwvQVO5c2cjVLa+jPUkgTSeUDhFNynxdLQSWv9dfF29G/VQ00/BOG9MB2fCKwwRsIxSnuhJ9Pv
MLaVuCn6VxuvbAWJB6gl57UfFnX7euS6HrX6as+sc1cXGDI2xlKP50mHxIGV0fBmP9393DPLiWPr
4BejmU6yGWtIX3B8mzwnzxatoUK8x7dyJiMJBXs9yVomjZUyPn5hG2V3ABNhy9YiCwQNlIRi3y4f
9Spi+4boQvHoR4W6jzXaV5UJR8JJ2whVfl/Bwy9tZEtuPgTRp+huvMTaXvTB975mWavrt5K0vu1p
35l9XmyuRtVjH56uA7MSOoVVvVEvvIIXsMXpjXtYviTHaCqw5I6s1m/Y1HCIjPK8r7XUZzWM2tWm
RrLDSWc+ffBXmz3hdnZHTW2PHRvgmQarl6hQ0GMnFTlQVro1e/ZC44mbchbyb5degMdxN4FPRs8V
AeD5IxIjsTCUGRmPscveXabyyyB8LupQdTUzN8T1P7eQaJllORVLqQHskYEZM6/k0CKvJeCOEYia
PE1MJEcqbBxkR5TxSbDwNIzX7LfMk0eQ8uqGp447jIaJWYMoM0xpPANyMPVXvd7a3n09rBArW8vx
YtN+Jk7Z+/qM/TFlBRjeFzEpFrXk8D7m/pngPxb6Dlhe08QU3g2kImYZuqIra0jMqy05mcne0z2w
MQEwXAMDHMdilG/OZeniI/soLT5szmdATPLF/1S4w9X4USL2CbryZfNqh9pu8NqqRs3e+qxDkCk5
w448+dOc8fjxFrwgT2J/cA7rOd0LY4FR7nIPV+/N6qxH8lrjGDOLTjWbr0K3nfLMAEzQADmaPi5x
DalJ3/wKNIi2zhlWY4GWhircIVytc+uJvlcEQ1+KjkO53YTfK9AzIhuBQxbwsWIYLns6LsjEAu11
kXyuHz5TMzr2U8bju5NokoWiIAzmjKLwU4/aJ4vw8LP24P54PykhCVdtPr70aEnwgLEucFbxQ9oJ
HZEPUbeN/Gf8qli/soh1p4qz1Bwwl9Yq9Em7jv/9LCc1NUrqwFtVBQUK3UBcniGV388TY2VjUBpM
2JpI5yOOd5ru7XsGaJNOufdmAP69C+SHKZo1gBRL4V49g8M4uPMwEgmjyuPfHVtRYErDGjkZh7ES
R2T0JE33qqrMPonRPliwWavJXz1nsgp3V4CJYe9o6AP8SNY0A0AWUJbTDrwks51+QiqefH5X7Jic
2PF7GpaWoAULe3Cucge4u+3bD90xMk2GXMgGvI8682Nn4lOAhObaA/WtC7xqHJQKayFeTghfLu9x
AItwQXx3m01mGmVF6DKcLpVO3n9weihxEAQZJrcVSq55bS56VcqUiLI0jpO0zmUwVJnbM46b1nHK
/kn0tgDKdVM8B+xk3ENWvltOFJ44UvDAtaskesUo9GG/iegzxOvrIA9FZM9eV48qs5hCP2uVd+yK
zosvf84TL/Urhpio5Jp4lKO+q1r9yV70SFAu3e8nnWKFZZN6SnUePs/SSeLiSHQ+XjTSPliazGcO
n0HzKxJoIjqn1BrM4SLFbaDB/TDFuD66Ko51zkkPRg2hNwI4EFhTQacCjkZAXha+rfSuMXLXooBt
V7Ote+lJD8ctDUIP4EvX5voH/mPA8Rk9wNnxVuCJM1Bo0XqFdEdWO+E7qzM4UJTvbStyr6mFqpdr
5eIaA0WQ2BAQVnIN59O1y7ZSqSZUg3pi3U78LHKotfGyEy7qBeHfTg0FRIej06vsVn505nQpwQzk
hoV/nAXZDwTHuqy45q8pXZLpWqwyY7FIY3S3bKvDIJVr5nzHAxa1ReDIuu1VxtwRb8tk0+8tFGXe
gtaR7u/pXERzF19BvK20pf14ZcYn5ZPl9JnmQU/Em5jMG0FUPKT2WZRQ2csN67+OMfGKDcxGz8ur
NSLHcTgKo2idSP7T4Iesj1faLqohlOBkW+riDoqbcQXWVioj0NnfHh9Z7zGjAKEs358iumgkkUB1
V9ZLCw6ZBfLbafVZziYgNqS0sg8XFnCQJhPJ12jpHHZtzHBU/PvZe+xQ22+uwLTQx/pcXanrFHIb
FPcmhct8fzZQ3ALADpXtCio74PYFE792j/Itcqmug1HEMOmXfMj4cCOJkRHswDnaDvEOP7Ld4ODR
ezBfbQXZ5elbuQjO3np31OvAmwlQ4LC0aLhyGwLmssHo6h9eccHyC0joFeBsyj48rQ3E0QVblHu7
n8T2gQGyeVAKrKXXX14DNzSWdN3EsEFDj+j7Wwgfahg/5BzdR3wEPWsM2Y/mY1zEAPv52k69vcSM
6GIQ1PJOgeMByeGGnGXgWceZW034umNVZKGd7ViyZ5HnA8o5C3VQ7PqknBO+FfX//hBa/TADIfLe
X10tVzpgWp613bXLv08MhkWP0V+vD6o6yD92BhngGQBN3E6Vobfzk1/CNVgmpAGTk/cJLSngwgcJ
qjwnHu6oxn4ZFw7is99d9U+4d+YFCaHBEBKLTiLtD5ujdAz6sPKymyMY17uh96pybnA8iYmlxlSB
E9FoD+3hOJ6vXX1hQBU8hoXheeAC5fRyd3xTwObUgWXuf0Ukvc6LXFj4BVvBNtQRU5ImtPINUIOZ
xvr4zPABDVv2CFW4RSvwKXYEEDeKSW4eB2uSS1YQTYEyM9450U02322kyII7BhEGHp349xf+CILE
K8bNaKyN5hjPDCV4hVBw/J+Qpj/Jmknko3MypFfarK/u/9vwLjFS3HLa47l7yx4aZ7xuR4PeDyRT
4B+q8FAUoCSRHIaD+viXnU+GnwgdFQRpYQrq0f6ZuB5otWZ224HRBFdFJKRakoZIzm7+diBbafYG
Lichc251pRmRCozLXwAhmNAFvvkt4t2QtArHzoCa9Eva7dza9CXiDix9W9v0mbtNpfZ29qpRB4th
URmAROLsJEflR/u67MBbET5Rx9BpGjd7ORwwVGXEhBarpAKv/PTcI1jktJ4nWrmmRRWfZ86QPiCH
+quGArqCGOLYftu+hx9bmKL5p8o/Rm0sKMxkyBFRJgoM0SFRgFS9Gt1e7lejYJoLvlSOKH+dmEwY
CPSuy5tE7HLX0q87VjVpwbsHfEiah77T48/nIPXO6V5yQ/7e0nAXuocnMPuX0FA4n+SWcZJsJq9r
IFaHTryys2od3XPLiyWtpeHSDx+wZVXGVj3zjXu6KFeiqTaLYLnFEvbNicWE3/XyyTRiaA/vaeOL
oNipl6TT5SbFYr4XKS6GDdnqtsy4TFqnbfm4boX1WAnPb9lz0f3zqq+pITKSM1abYpQzNFwRDmdl
3edfpgt15MR5hfQthSpKSWYkE9MsTRwAxt7IJmVMuWzr6q+1M88bW3BU5EPaGtG/s2ULu8osBFyK
/fUaBMZY3P4mNAkPuFyJtz6SsGlDi+Zz3LsdI0Ykur2BeJx6wZg8t8Q/6EqY9qvkOAewlg1Cgth3
Ice5YJq036SVonIVRj++BAd26MWUOSj+oS+fcfBlpKkY2hvOdktyr4jTVf+91u3rQLHygU+2IZgH
w26jvlGvX2OmpPpk9p1gjz0EtUlB6qwSTu7DW4CjiVoePuDbDNWUHBNeb8qtfDRCf4yKwpDSyYAj
LAhd0yslp6P2BMHv2fshEqaGKzkhq21UYSsrwrM3Ls1BhnDCeexGO+uclGP19gbWC9snPgK1O85B
6VD23O8pVFzOyhDxwkamK6fTb4IGotr2Uvw6f3L4PNG424AvRsgg2peoFUizs7pLP+vuWIrHUNis
bijIJAzg26op6WjbA2oHhYXIj/XbSRepe9Wlz7LmsSTh/fTwyWRG39OO1xlr0YNvp0EfvX+TEPCR
q3UF9H8ZKYdfCwmoW9iA6Dupml9CyrecydTT34LGO+qbOp6hcefEo1ER0pHDkOl7PM9usqjtfawE
T7EuVufx6VHzad3DcbRYP9xXux6XRxa1ysMy7J6KOe6Tb3BdsRc+M13N1GgWP+uGJJMiwZdMWkGR
nk1rh1JMUxW+Yh+dOTrK6zMGZxbuq8dr9qHAmix+1yzZYMX26PJe+B9Ek4OWihNSPEOCnfyIu53+
r6CQcR3qQ077a+pBhqk/ImYoVd/WLXgO7deaXR5sy9ft36jSxYb+AVwgv7wmXoCeFbNuncBOClK5
zxHtka2dTOxrYN5p8mfWMIloYOGsWOjaJVjKms4gu8oejvU2OC3Zu7l6eyyUeCJ8TbX3Lix2AoJo
V72SsZ8W/M1PZR0zXr6CWSbodDps6v+4TdqcwURaYg/gQE452bW2HueaNxUoUufDroaiAfwra1+O
8mBcub3WBJTWl8wvvSsQioaEeg68Ow+dDFQ3nvXtSExQGJPMeDlvsgQpOcf8ZkUvAFfhj0cGos8V
9dJRl54YGRrJvqUDFpg1MC2jRKaEgMKqEvWyMM4d6PnN+F/BeE58t1VH0B30lYYSpkU/mQzZtdVQ
lrAicB/Paxb8ljl+0AsYN77hAyvwBfkqofqjX1JTiu5IPq2wu/YpvbVL36mNcs6tz9A0to+XA4RW
3egePYz/JKFXfcTURUvgFDGbFXIieDTHqLTkcvIbTUwsUuYAoPM/T4Y4uZ2ekYTaDlOcE4sf8qA2
rVpADVOa8ujY1Lkk/1u8JcFrx7ONbY7d3u+wb8yx/SW3KD/+Hg/i84cL1f2rHrqCVFxrjW+/Z+z9
iHHatxwBUzyp5i3s3eGhegpewpXwmC8dxNkBfOnmR9jHMF0ZgWwFLdu8wyqcC8VGkE2M6y+qVAug
wOUV2uqFJtKCt8PfT76l+q2j3C3GX1d2z15jGscyztiM2C18u/qdOzU52S77LazE3uSTNaS5pyQQ
1fCe9WHl5340dyGn60JzYE4wg4xHFIXvD+jt3pn8+wlZ4KkG1v7AQqVhFirjyGLzNVUaCAorwVty
5nd1xNQY4chN+xFesMeuaDESYD+JYsBziJQ/eUmAfMO8YUN76M80u4OpRnN9D8DoB26+JOhT+OCL
0Izh/5EnLvNsKdjapii07C96EFs+yAQaRuB/EguwRj6AW5hX90KUgAwVGSOGGdInGc+iFiJwDtE5
voD1DbyzR4uFcjAQCpmnca8TYkoSV/OaqqUv7fjocK14BoAZKCfJ3SSXiaJObKqKCI7J7HSIRiPt
FpP19ZENiXeFjGLrsshWbmKGbk7ISaAmoN6dkU29BviW27qAhZheUmTymA21Yu1EL9DfLxzi+l6U
wW26mHBTvayo68Ug4HTws2RKf04DxSDbGIsFcySEeDeA9F5nSDPsawKCvam5zkdnk8qpvIeQLpzU
wXcvVEj6XZdMkQOEhMPKJ5Z3kggiHBdYS+PNDN/Y2fH7r/G7EePEgYbjgLJ3dpTgHl8ZOUy9axxD
VNBSu+i4Tbj2YsuN6qzG7hi5OtHz522vLNbXgfn9u03lYUcX/4q7kYRBiSf8xG9dUAlmkDic2WHK
yFo99rhc9mfA1w3YHmyI/N8RltrgVX8GA7o9NIGMzZb8ddrva/cZOZFGW9AwNb3XbmP15R8q3JTc
YLrPtScM0Fi3yK4kOL/PF7K6R3AMt1RtdOgjeBRYf6Oyzue2ofgEr766H177Kx9Y8qttBbjhMUft
HEgdmH7mjecWa0cVkOLaQjbejgkluQnLQAkyUKLgf4XcMNcdfK+rnQkTq+8iDu4fpcHRlNG9D565
ehnQvmuA7PKwbV12RvBKsNVGeDLWRK0mZ0UP/+05XUUEk8gTjCwSTOl7qfv/GC9UhLw7z63Rjxe9
6YKNBK2W4TX5eZFkGtAEGRYLRB+UDxvQ2gyN4V+Q/LNKv2Azcn90e43/A6KTMxnOkUv/PbJPebUT
1NYlU2G3ngIROOrpcmPEiGqUUZzTuOT5CHdY1BhFsxX0d+b2/6qZ3KtXQ1OMoRU4tJkzXF2PqzNy
89ouXStyoaGzeHtombqCuoKbEReLwtKwJ7gpk9Rri0VFC855MWOX9h3La1dEPlM7nGs3rtfDrXUE
K0I0BypNxe7y7PXZaBLWC7Ds1NDklhPlnT5JWX3rWCOeVGwrP1PqZqIEIz0/ZgTxa9mKGVbjI+0h
pvdsFc+3hGCBC+Jk7tS2+f4lCgjpQhJqy4mwQ1YPhd3u/mRAdHQDkof2b7FHXMP7iU+BtKY1aJ3v
eSMul0e87VDxRC3oR+MyArHvdPz2WsgzVFhYLfhjQQhVkV5TzXA877svXuzWnPz2GCYqZ9SWWeav
NEw3A2UquCer7cvUW/BeA8RrJ8MwCGyS+tL5xHYNfaIEEObaJkqigoOVtMtipMFIqbU80JV2FZBH
FXeERDw4zHNata8idCWEzBi2E63qBrtqBq5Ouhf0u/PH9RN6fzvpfcRMYtdENYek2c/5fE1PY7sS
DKa8vJ45+1b3j/0ocQHn6uArBeOSCw4eQM2jkfNB6HdWUNsrT9LQFjZQ8fHVALyMVVc+3u3ctymi
yogQ22fHRFZqnWzRtG87Qeem0OFjcvOHm4pXC4CXxtKeZej0Pn/vKn2rNV0Fx1fQC6VeoLhQ8pJ1
kODgqdLS2NloUWBri7pu8O64inAGihSHrPHPZC49JukzvvTg8BeMetI+BqWJ3ZcaIVpgk7sHOZa4
1ZjwzsL+inlXqwY0UScJUsg0PyenAK4qGrgQIVcAi3eHXOQJiJCC1IR1m+22ZMeNxOvGfAQ8B5vS
g5GSsHq8ISICOm6oO0iT0F2HtqIpHTnly9QGQfiVXN5/+Z275e2vUmtK8BYbK9DXYp2iW8g2/AFC
6ypokBID7V7b7FbYTSCsH50rp5EL+krPmJYBJ+OqPk6JbS8kVN3MeQ37HnhNxWmVmwM4gA1BXtfe
jQOPqDeH0suEH+6fOKgGeDMjsZtk0WBKa3GIUyxPEPiYDCjxk830cjvpV2Gpre3cjvGasQoVRZv+
p7NWoOb5ivhNHIY10KUoz9v0obqu36e6aLSnWX4oiHyaiKf38tSrie6FQAMSZnma41dcGh7b+8An
zGUufb6X17LWYZ0jPLCBZIsqhf85Yl2YVTkyVeEfEEGeHSC9Jhda7ffk76cd1IRfwRSb21BLA/o7
eFmFQNovltdb5M5be7tyldXK9t3Jv7OxFE2Dj3hzOxGzjokKGhnZTVm/lI5N5W7p0/oVBzgrxsem
QHKLIJvbLwKXs4kqjHWUW3Nvh/aVCW4R5Wc4kKdbaTE9ickktSUZOs1FtCfriH9Ih/H8tYttILRK
H4KfPRNQggBAh7fCQbgMhITILMG9qw2lZiY9rfey3zN+H5g7nmANX5bFahFahAlSc1dHM3Yi+V2T
KASDaNJZXtVBC+lu5FOfnOsStLhnPjIZww5qgsIcpIBMqatdVyWI9MCGO9Cv5+w3eLUVpYZH2Lya
rKh3PETHOrtKhk0ofCjv5nCHukVRvaTXipp2iFD42ZGvaG1lju8CZ0JjTqmAdFatHLrS++ouQ5ou
wLPWkmvrZ0df2DGvegCf/vbbAGGfG/oEXx3gnR+SS8w7NKlrbk8fl1px1bpmT9067aqpLQ6s4OZH
a7UTg70fIxFtGhwrazzcKMT9mSkG2sB6KzCrCQ0He5m7ZgRrna4EcjkKWDcW4/BHq7VmYqK5Baoq
Snfhh95o4H43aIqEUJcNTbnymTZk+d7EetCs5NV2FI7Kuz9Awi/JfqHMe/n/bD1XhaFLYoikcvto
oQVozL1Ecpkqgw8kS+RIAzzlv/A7C4HG+uY/Y/PHJS2LaOMOMDBP0EFCcyEzZW3PdjCQ7RuvRxEe
HEpv4lIZmKPjEmAFcFmRoGUNz9S/UKJOcI2pgleAfh4Z3Uh9eS1AzOP1JYz70W5TkSyXasdVgXH4
9TF5sb9lA0dnAx4Xc9QHrxkec0n2hGoaxGa4mmRzOGtX7aG7/R6VnvWWpGCJhMEDQ82C6VirT+SU
UbQLmn4Msju5hVEJEaE1GHCcn1yviVBgqOa4GJwF0G+Y/FdqAt8PqCwFlx+uIK5itO6Fb4DPMKTw
79k3upopTs7yE8dVJu49oJT5XLmBOdvBd/eFX6iyT8a3Fsw83D0AAugpUXenol/RpGTJxg7C9xJo
ZlzkfvFoQ6g8CWXCUpeLusI+3y3ZzhQ6kfwakrvwjdIf8PIco3p/ro9GtV6uEX17NEwN9Wv14MWZ
mrnwcs2K9/ifKQHdSCczIArEdXDepwI65U9ebAgNXHOvMh2vBo9t01E0ogb5bt/UiOERXYE77N1w
JUnCUpc5GPwaMTWqrfNcCpZaxR1PojfqcAnDNZYvqrxRLtFt6o8fBEO7IdKecbX5ZQkn5cQXxK4l
1vvwvMVR+MLJOb9ph3DMhlWZwFtDyebAEjnh7BIwRLseBTryKmGFB/lfV4aE+A3VHFwLZSxbRf3f
wU4UJ9lsubu5uWnPsxg1xUgeoDZoUMpI3BeE7MzBTdtPZ2Q1QlePIZGKrRB+BAsuiTVfB7tTGW0H
2xstU8ZUs67UPWwy+sBZfGO7tx5lXu9OdF6qRhKOdSfdH1jbUESOAYGlZEfOgHpDBsqH/z8pcH3t
WoiSX6s/13erbeVjvpsQULyWL150emPGG2UuKlmqXmZqN42zI5lO2h1xgpHeFUPr9flPseY3UyHc
ba9Xiqwlz0FoRDltzBIeoxGvOJGRmCiaEVjMDVppPrIiB/HuAs31ToHxwjmsWdzymh9KdoMAsUSw
npQsFS9nBhe+62ZiuxKtp7QGi96sgCOn1La1MG0MVpgEJG6W0Gfxtn/vDmBvj53rJr+pyMNnb8ip
npguuRsnfGLao7FGzB0Tf46Q4majVwyyEfj6krySIq6bWdh8stBdod/eAqYR9X6kfnuW5CkFGrH8
iZ6oO9lpZIY0ujCffK88F5VDcJyem15JttJ5XsmAmK5Bt12CTufNevCLD1QzkvFwrUSvJ4HkoMhl
1fkRTx4xl2CvHXJik1Vpd0yccEboU66ZJvRrukQGfZsE1fIEErZkr4udAAVV+YA3NA1zKg0xOPIj
VDxDmcnBJHXOUcVTJSC17mQj6yQdaOmM3ZC68Fw5brUretZoJRAR9O1VObS5pMla+N9nWb7WVOVm
Zhd3YWgV0YZDEbigdDr7WInFcK/IUBgpQtC0BSqkOkMOf9Rm6JeAX18GOlWG8B3XIIpxXpzg4PYV
X2otx7JkKbIoEBYdD2KrgXjm/+AWQCLag/QdvYxu33Pn3pSWoNslztxDkEOxzjR09UJ3lQjKFD1K
YduNT836/C0EI+tytu2lHxEIlw3M0N3GAgK4yJonUZI3apfXlAyfw4QkY8YhGizEnUVirIhh8IDn
P17DeoIrDjPRDr+QeSqPewySY2ce2iI1MP4/7twZQXmGEbHeKw/CJWqOMuQnkbvVgOaKejYsa1O2
OmOPP06cadFZVRqSdQc1wu/Pvjn1LAIRQE4yhv8LeXBBrzXUCkk6Mruwkwe0GOZ/izm+yLhGMmS8
lSmvRMwlCCfqDWBVApWsV0x6L4rFLN06uKN4ycL6debT/hDL2aHlslgXB8WFfAlCeh7zyLWyyM7w
Sb0GgSfaMzj8TA4Di1luhFPkGAd9XdBBJBxSmfta1HMew7M/48CAwxjxdwIymh1puKheF56bX9NG
8z88wycRkgQShgsI4xoLYjTNCgqnSfIQ6ti2ZYTeuixsrEYFvCsExkNg4x9dBcDW2xdfnv17IVDZ
Zei0hp5Le9FrvExgbcGmbpn0Q8Vum2jdyRpPpEMtk1G6BSnFOrQybb4h5/WNllNv9Rd6WMAj5E3j
K5ribIOnQOvX0G2gLBgHY9g7H51nEDRFChdvkkgC98Rt+6N3sRPy4qtb1Jgb+QK+x9hloq+x9QZn
d4AKkRLCCz/7wyqDHHlsgc8oTKgoki3UfVqTzuHiU17Z7SevjlvVmjRrDpzT92Z+Wcxn6A5cUb61
B90OPBqGG8BWKCtXWXTwqBHiwHFOuq8IUBD+sPG3p8TsiynmWOnj+vL8QI6RShhD1ydbMjVRHPnv
X3bEcMbs3kIc9YSVZk/sYwsZpBZ7l3ogvLWs3YkWFIgy0TOb1yEmf17Ggx6prkDf1DYeMDQk22vj
mC69l2+RbCVXrhYeVAlYHWfXvx/kbZfpIz7cu7q/xzSVRdfB0498I31P8XY09pfnMD08kbx/f8Zr
XS5nEjtRO8cw2s8CQSS0S3rCQ+47fVXF4xswM+VUFPzJitk7CC6qszIk+jCbsYnmyV/+71h/IJ3r
VcXpETTtJJIBYRsbsOzeaU88Wv5ofxn5XvlED2882yJEMdFn18MMv/JlN5KA9zlDCPadbEtdEFZs
lzSUkl7BRfFThp1wPyPGgqqwgUUtETgvRkU3824oRoZc6/MmLPHyB0gorD/tRoGHctD5JfaEIc0H
lZlQQl5m23o++TOxvTdpPFemFydfY8KckRhWhcm0j7Sl9XzMp2g0IWXlNMDveOkO6f5Y/NISSsSE
zCtgQafxEUDfnZsrBoB55gLhqommwsJJQclYXYq+DWOSL8u4+3b+9jvVeQ12GuezTp6ow/pegBx2
tU2lD7jQJKzxX+yrmW2snsALRFYFcQyQYCh6/+cf4rLTXw07ccGOPmwE+AuVO0vERXf/IknFHeOq
HzHXpSPK014qJoLJrhcIu1qzXyBXCr3558KDWezwkWQePPn/afRsGz7I9BXbMdqjcS/SStXPtttu
6qDfA8kxPo++q1hKkcRk8uHvtsEQu9OB1n8Aw/Mp7Kv9L8q+7ul64mjZKmj7nTi4uFLn/o7XgnJD
OePxFHtEvlYfFrr2VBvLO9ALGZDW3pOxoIi9Ok4CsEkDOLFI1v+6OPquyzCXxOH+JUwhNjYC4rRv
UHoKUn4PnHrKngiMoqmK078a0U+bZYKWiPCjFrF2WjO37PDO2tQDX9vF0V5EqRGesBVJVnaANezz
DG2MHfZntpAkJfTRjNClsDT2aOTNafIqGEgIRBOTU5DSVq9urZZh9ij4FWhTmath4cI95dW1YRij
pY52TcP9/TGeOBXu2Cx5rmRwiVkGgqOFNzCNTcUT5RJeFDkzgWQvL8lRynr2b6zKmtYzTqgFyCvW
Xqrl4u2M3A0HXYCkzAe4dghJ+tVjmYOPUDB673lZV/mCFdnD59JiK4HW9N4ATcc3PRQAQ5+QFngp
NEPR39nJ3rXye45V3ZvQfS6LE44LHUGUYeJq0tOMWKT6WZ0Bif5Wm6YC7qA2deMBV+Z1oUKtSG76
3/eLCbR5n/B7tnRTtiaKIze5hF4Mbvg3hTRwxo2Lh/EedbuQY9ItbgqhkQD3NggAoJNXB3Nc9dJ1
hHwpLMjEVx7XjmpOz6hwZjFbYIUJiZTIQnfNKgM3DvdpYgi78WW7A29+r4wqWLqnd46/VzWbfI+H
6wBUYWWOvokuu+4nkbJ9c37qbdy7a4HiqJFRrsyDbBwmVBK1DHJl9vaaPTdsV63Ef5DQ2MS8G3t6
yd2GOEWg22nHef/GjQ+hkMHPAIMq3Cz0duqUiaVyb44CfIfqaquCvwDl3FcI1KTgnNXlpM/Ec5Ka
A6uUSJDFPeKjZAlWwjXMgly4aUNCrg4o4FC/It24ZRMsqZY3FTEOuQjTMh1Ryq4sPlq7UgDUH0Ns
nrFdu+F7bo3dMZerkX1lVnQ1SDXU5rlcgqFmJ01BFacDcEpyHuuN2bhzqDe7F868SThzj55J9K4q
azAmtwmAEOhSJeV7mlk8UJYXV1Vyc8SZwVGgHekSy86uvYxBLK6XcFIM0if9+YFQU6UwJxlA5Nu7
KfGT+fIdEznt/WmKmaXhngKIG4qD1rGH3TV+4toiwMcJLYuweuNCQQ0XqvGF0MpRWToiOorilR95
o+QA87SEO00c2uwtIQ++nyHAN5v5U5jygLsBGjm7LMRFWEfh6euYGjvRKfSQcWlJryfP+H4qEKQT
Tr3T4ZclnPInanlONmFFuTs16n5SmkNmfAB2peNQO3xU4KMF6iemj3sawRSgygAwpBno+fbkRtpq
7S1VCWRANBvfbxqbZ3JMhth25wr8Fz8yHdLzXd1A4lbgofMOO6MKDc5s4QX6xmHhCKoUtwnYDf/4
d4vCOQuMLLr1iKrXAql6+z87brnI071sE5Be/VwZxaJ4EkG/nPpok2btxLDrnZZ73q81YnxlB4uQ
+lT4ViAD046UHcOtE/zphBO4GSLyn8jiEGEj+vjrBTxxsCByc/0FEOvDQWbFY+6Q56Q1LXVWLHL+
DtcmuEFoVOKUsw/h13CzHxHG3JE/fuTSoR0gKneTshkGl7GbRNi++bCsF4T7vgTdOEMkcZTgFrUg
p/k4ieT33yGGZOEO6HFWf1sOI00xOz6XwAQAJ8dHy9WIKN0sTdsbFyDOAr5zZKmRrKZBDjnRiC/I
c/jw3sN8gDp8xDY+UsVRlK2qZJVVzb+Ge0olYQzMn1zLp3R53/E3WquAeIKippmCMB3xXhfBoWQo
NFS/MdAmZ6KRs1Y98H8APmgHGjTIn0nUWkI3yt6QQ+1H3itIGI1VkiOuV7WY3/1dJT1iomk5FK5x
8rUnfKQQPj4KVW+0U3ow0SJE82ySwbWsVN08C+J0nmRPmoC4IyKQUvI9CLU3FPtCwR0cUOUrXmJH
9jeKqYehax+xX4E+0bgHYw7V/roRuZoXAbx7xAMP9z2jKMRvn+ek7qPNj9bCECraz+LJVeAZ+D2h
brvY70m2E08+NvLxFP4z0II0iy1LYwyVvhOr03ZS/K+P4EAmDHj5yVLFyJdrFQxXodCL3M7AbAVk
X6apcAyBUuP1Xd6rYUIzEKWVCE8tTjZ0UqWErmvyK286a0xNWSirLp+w88wBc1q3JRKTXsXBLucc
JQCdkqxTAXSlLfl/aLqkTQuvUVAJP5wLPo4RPu6HywIw/UKuQOWObV+Pxxuh/u7raby8MjiHopYv
n+EdQkRKMvJiuIgwdr/th1/xSjon6hnHU5qvVVEHuI428hrCIwJzcGDPduHgc4sNGsFbrtla3t0R
mD/X+tqXuvu7WrwUk6u5/+zkerpMoHhX8HUw3qPrKJKrceRqXv/dt44srLYR/K/J/CJoewrystFw
SFuwLkyLkMLKxBDg14vqoi85FHMkfA6m0kfBzavUXeePVRM/wEMyqJUC2GecgeBlaGyXjAqWnr1s
vsM3aD6Nc2GtDCv2QXqZCqEPXAMtiK07vstY5BSXW1O+PSPFahCgBuE/E/OaLWTWFRT22NzQMXRy
xyB5oQUCkDcPALjYqnPDas7AXrwypt+07Vq/ijJTjJmu4rE+QEbZ5YxzPL0vSA7s8ZAl/rfyAxM7
XWiS0iYnh//0ykIb2Foa7lSWYTe1SW6/qsz8yNbcAcWnGTxwwHLPt6HGOJdPWusR2qYyMRKz1XFE
y489kEZrOv/gY01T/bHOCbc4RK5t4nzHK8ymwXt8B1NB5CPBIFgY/uzgLZtNq8uEkNTzaR8NGPbU
fIBPIHQKQY715/tkauNveUxU2lWOh6ok24Mh4zg4jAtWT2f2/RjfPBg8v4ZjuueYzMJUatjdJYUa
+n+UUQrgnIT6QJR1OnY/IouNAKydiQdJvtN2kdmk4SEWJeVc/2goNhjpWa820qi3jExateEYVO/p
2CBM5RT+imll2Xdo0wHur8xrcxLFmbVgPBdSpO2qZvBvT+4tmoPc5hLyUKNDKDRKknT5ODU4Kdo1
a0UJG53jKoPSy/tkuHtWrkPehHk8jG3LdB7FdHcmZIB9pONvfJdMJBJIDKZ/tTWXDBK/cMihr9HH
OX5NUxpM9RoxtKvgrEgxeHfcvOiLjRFtjkII+If3TlRzaXIKcJEZ2hXnFdTXyqSh8GAZmvDCbz7I
6Ed+Mz6wDRJlArvu1XPFEYt/+O8wacnsZDlqbsGE3bGkzbMbmeBSMgEpdodNWChx44zh4OQWktok
S1tzJGMbEGtexLDFLLffRRlNwHsQVqcxPTsS7qJRHvmJBtU9CBBGrpAC/oqrXeyHdWATRudw1MWQ
bZs2FNRTXvn9s7BL3jf4UHpS0gDJnUzb5V4l94rHomMviED4CclbIW5YqEoAbWNc9r8mGBsf6rLk
gRlXQR5aCpti6UsBJFJ6YAlMksB5q7+2iqzLem1PwZTecQjOoC8mN4jzN2QO392Ts1nXp38QKAxX
OIy+Kv+/2hEziiMhefDaKGQ7Q74pXOMqjBn2B01o2H496dZo+eKULzkKVIyELNLEuQFhes+zu+gM
tKZj3yEikqXYeZo57ASFMCUJd9S1W7ZpKIgnBuCw6uesWYZ2FhAky0jLavFaGPjsIaF2vBaqxZy4
4xQ3OOIDlke8Ne8KM2zURJTn4NgunN9bE7EP2SXR+kgAukKLdyztdw9JCuyAujX4Bz0aiHJRoOKI
wf+1REL4Il07gcqP7zqeBEIP8gX0HZc2X8ex4qgZqe1UeLp/EaaF0XMaKJxPB2NXAjEJXsAvALCU
CmZ5JHky7YumyraWFKPi9Vdt/sH+13htBPWDqBsML7bJqlfUqDvCSdsIEsp8CBMznQ3HrE0QQ/uA
36Jfzc+K7ch26dxDJnFVxmRc5rRWFWxagmsNHlaauI3yvDELssse95A7CGbMEjPqcwoWJ94IM2Sw
8l7st/HjX7aqoKnIWJFmO5VpscNB2eh5aShkjY1aZKBrE2uYfEknpZGFIjLsxaqzLQccQypWzhJ+
PSVoyouDYaSkRLNMiLU0NfsYkXwxuMl94VRrLtoHjgMB/3A7u6iuhM4RFrdUDHr2lS4lInm9RrdM
myBTJO6XeejFy8qRS/1cMaiQqBGAOSqmxrZlZcLjIlYSbUoWki0g53zEz1cZLf3Anquvof57oiPu
Rbdqvlo+HapXwKtvUGd2fbOqTNhT4G2Dqgme+v6pcoKTciwORK2LQ/geaNMBEbRnoIRVvDGFQTcY
nslJXZB2WZlH7AtWhnJ4dJcCNX/eGTZUf2mjKUcvN0RPDOf+vsVS8A06KkrgeOZ/TqbN1jkDEPJP
JykMPpyRi9b909DRR8lgtFSBEBaBAB7dHxn0AUkGWq4bTXBLzSNVcG2FSs3gJnNP9PK/c1nEQGOw
uuIb2jtScd8EdMkqIR0myN8dlZjO6BiHFz7FmsmDfNgs5Lz/H4HP/u5brWKA9537/6/7mziP+WCA
le1I9DCgwmS2RySqRJduRGj0yEGgtC3Teq3wPVd4Q+bC1fvPEGU7Wa4+83ucfzHXWi75+pa5IyWQ
CzOuRJisYwMhYJ/qdpDbBM85rcK5fpMneDgmWDsRkTdVwCw/ZSlD6x3kUnXRwpKUC7y5Nt6fkKay
w/fAoosLeakaKdWv2aJHj8GwDNkl2xJbiQu5MuYKdPBwLm67NpkPoFW90YfWEomMZaymCCb8VYaj
CbEwEGa2diU9JNzIStkSvPbJBzsiOeNoD82yTlyXaWBhKVumG5iEdr2GvxBYLlOqMXP33551gQEX
sE1OuRZ2Oa+6th/SDiCnPS7Rag8yrGRbwAXNdcjQPQZ6U5AsXENORqFuhAYflEaRp2NUp0qVbdo6
IjIPcUZ0EdigeFbBfYhbs1dHkHiPi0e7dIn3tXaiZ0ub6c8ekQjQpP8g4EOKZN2gBaCfe7voXdhA
8I9GuIMsqifx+gpaWDHPKezQgzsWRcYdl2/0qfSD0mGmS05bAINq34KKc4Ui46sNoP7Jjx8Y+BFa
IASeU43STHOT8F0QDU4f+w9+bcumrJQRHiYG7DQomgl9vBVE2J6ZFYEF23Us/WAYzBwFO+FPDCVo
0p+cadyQmkB5rbvARxJ/8a2Bwhri/X0E5IdxxOKtjJwBQCzn7Q/2ajWbjE1Cr5wG9kM8XuQgfb1G
BVIKgQnpw+fSilRpKTb5BbHUK76nLKXAQlrpAOarxxVdGZ6R5RAcE5PgYfGQfCREzqCSI08YcHNk
//nEKmBu43yrAN3zahKXeH7GuXQPcVSYM/89t3h42aHBgORbdHkNbpTblQVSyYQt7eFOyG7vecuV
ovEbzju+PC2G6xypo3wcxex4Z5fRaTam7+7eevqYVFZK+mLjZ5zJ0deTJhlqphlE2urmu4HiLh0/
DWQehwrFidGqdh0krxiNw01xgdKVfw7Ga6zfn48oKvQPZe0fg0Y2K6rxtxfbA96YSGYnqeHIFhnU
3LFq/YiXgIh0ZyGIRb+KpvFubnf6nZ4jC7sfuE5jdeWgfuGZUKKTOtq290K0WAG2PsvKCQPVw3vy
FSINg/oYoaymLdzt477rVpIRafkgagg0Wz9BbawfusMq/nkUm5a24XdPs09bAjeSgyWkyIxzOt+k
SwUNP3rfKeVvZlJFNcEWKnrQhwpSUWmtbKLw9CietTxKpkdanXE9sdnkT4OjIK8nmCnS14Hx3XLZ
bEU3PVLI+4KJU5marXLjPei6R5NN/Klyb3TkLadX4C/dq8t25QUiS/Q+Uci5yJzWCFK6BriPTC2T
+a31Ydr1Op8ZY5BbP0olXwkbMJeBhrIVHwzKxLUrIORLFjY++UKBJ9DSwrrQl/YzH2HL14/ffOxH
3mSA+XKl/ufjHWPSkxLfpMmDPCA1GBBxyG2uccMHfylKjpDrPWpW2RlL/ZJhXCd0f4pWwm/rhXiq
Ckx/bARB9x2t0FYoI98KxKvbsIr694RMn3KZQG4NOhi/A7QpHJxtcdGwbM0ykXn4CkIiFWreoH2h
OS6jOHm7xEU7OFT08keyB1egy+jQ5oRAUr9Z9GiMtPQsb1MnZMFde2WMctsa3Uts1W4X89NaYyRU
DS7Hy1iW7OXE1H4MQvsyTGNI0cl82gONNpQQseEruQD+/wbu2GX/QZajLJudvDYTEa1PoahPjf9e
Kvamw5TJn/B1sIizNUYPCqkhDknKjxycyaRg0Ck2pP1nH9BGfOzovZsJEz6ZaKEbgQnh0CWeuB2H
4Yn/yCOpUQUauWgk2VNDxpR7neBSm5faB8+u9apkYQuDwVJmeT7jFxRsjBH2kOdwxovUPtJLyiLY
/Bb7t8cFBjFH5jnNKVTv6GcKR/Q8/7UB9kA+0I+EAWUKc0Fmwl6jE1rebAO7rrGYPtQWDxAcMDJY
Oi6Read+nViubZ8QChQioUZgKGQl5NY3zCa8/jDQenrc0skN/A06ZkuJcAjFyjCJE6suFeKPtSuz
ZZMr/mkgtO9x3d+VtYSPjQW37H6ISYPcWJ4uUBDsA9WhaeJQmhxREKfhemH89it1S7eZo9zR4MZH
Q1D6DEZyEAwud3J/2P38m1Hm8tO0fEwWmMqk6f496AJ1O1E67R6nqBrzBrsx8mYSCavM4CQ8TZk9
VUcxM/6/8N654arzuLGv5CqFcTtOUx1DDsPMFHPva+FbTgIa+E7xFHrE3PDAJuONlqRqs2i85N/s
CgDZYKRZkT/wyoyJ2gurugjQGA2vvsOGdgDq6CB9Cj/2d1TLz9GZJ+dslzMUfhtsQY5tYsZeg2u7
fGkf4URnzmVF+cDACtkTW00mFfI2QggTNt1jrO70ceb5LPEFIz64snExouPeC26VqB53elzKXoDr
7gP2mY4X+fHq6BMBAsYoY2msPfDqygPLRlxscDejuTwuj+lRCZ+ppYajE0UCLS9K59s7oySbWLv5
AQiJnXULlqlptC1K+h3HtPZk8bYEt/5RSwNKzq1MKvIiPhdBPwZ6Io1uC4wuENjUanDR1nD8KXNu
3OybOaxMsQdZ9fc/Rc1tlyjhtddlHKZd8NhyIuWLNSjsURANQjwgH2HHDcdOSll6liDR2sz5aBXF
Hth10TwH8f/Mv91v7p3z2SPFem0viQmg4F8ZI3f4aXKz53MziLvjkVb6tOQOdFPm4OChB2hadEl1
q6xgQhDpFtx0CUEKCBkHx3zYuLmQbFbssspEFwdg8D37Vp2DqtG1aPVFEixEzbA2/AShO02asUkW
1Jg70xC8hXoRbl/ki1E+m5lS3DE+0LUgC51XlmYeLsEF8dz/QX4EjcjtVeJLbqrYVpeXyUS4CV0g
KvjxJ75tShw17I8+lxKxTlCf8tMqWmFI4FXgNg2XP0upDGXu+hZVnNBNNUsnZJeJQIegEfxnqxu1
Hr2nweNGXJiIpy6I76Y3xCv2gMbsWEJ5LWA2iGPuaH6HFsp5Le8m4HGzDB1uyz6180+4T+oFU6Z8
U/kWyLgmy6XXJw4Upo76/epEHczGm4wrny7QjrbvfagRZlsNfNeGZlS9PAylAb/QTwt9O+G5KKjE
CDnmqt72KFgV8v/mxBgGAmwgUAAQRw1XWcKkM27kkFRrDVCsjU+zGadEOTPLJrkTXRojwts4iSHL
zMjnpxBzRAvWTKabuIf3oPlRobVrI8rCDOFN2HKQ/XmLsYMW7EETzdQj52VCHFtIqkKflpZxG6gR
/mjasfMZDqCJMEn8MEvCvoTOwF2dCPbjXI6kkT0XdFpZJbOZSLhn8U+i20cvaOB07Z1FhAh3Mybo
pTbMWscmckH5pC3j3mRLRxfTuX5udqyBKhyiJOHZRsBFHa+6HVMR/1qy8L5Ru68hsVwdcLpN2RIK
t/UDzHoarKc910+yV87xAbiX9ti2t7XOp1fBfenUJ+x9oMcIpqgbZDVbT2mwAJ+JucNY2kWYapCU
dHkd1w3c4lFN6X/Z65ljwA0FO5ya8Prj0W/HeNxpJX8/aHB0E/jmcSAGMatUr2egXRCqZ6M9xZVQ
fXOpQUT02BTMuYd4qvlWIIsOIFJGhxOiEzEpxG/yPS75ZvCk9FN46ucqSk4rUy0RDJuiUXG7AEEG
DYM6SltuxbSeicTvBQFFEjb9OHzY7eThAzTGw4zjQcvk3mMmCk8jkr6FXqE1zMSKuC9NGaLEmqTT
L4IcjLwIKGtu0i3BCzYXD4gwGWhZFXsAy6XedGk2P0n8vR2FNrUTntvJTGk6C7d1RvHjZta1XuGQ
GK9TUT4PsQHCHQsrhbqRIUgf8z9+nWQZktR1uqcW+pDRUGoW74DR9X2Jwi6m6oeztjktBngYt2y0
Eexev87NMdONxNeLsnKeYcsYKNqMTZuXJhAVVdyZxQiCryQ+Ru5Sp4+tbk6LvzQX/wX1S7U8H0OQ
riA6hWDakrBGiCw88uYTC9iW4YhPrJkqfYrxZe/UiLrzQa7PAXah1qS6nx3RXj1puAdci/fEbYo5
nerwZe/kWLUJfuCle73Ku5g8mXMHc4Hk44jnX99bv6ZAkPvxSlTEHdvb+pAEqiCdPtJDMcJuUO/4
OZ8P0cR6wPsxZTtB/WJkP5zt5ocfekBggbVUD8PmAJjKEVnWomvfCZhut1JJQ6rVIJVapqBKgt2n
FcRw0bjoGAYgRjFaF5uH77xd3tvH4W6XJXPQUlks1pfWtJMJEx7nmccFdUttuN0UKY1sUl32zJ0R
RjOSucr5k62jO8xGBbLu9X+Vuc6OdaP33Y0M5Mm9DmG6+Yql9Q7ueSXdnS3Qx+IY62ebyZI4+SuC
2byMiJ4Hwspj2bFuBiqeW+SxZgXkhNZsZQ2ZpCjomKcGj7riXNxf34qXxV3bEmisNyWqGZGJp95h
hF4UlcuvkKS45uEH7O/0qDX9QHnis2nsGSD8qpVU+E6TMvwKIKXLsCx9iZLGVfr3+zxhxIMZv03T
i93FmJgbNDJ9OnAeC8o6Ua951xXUpG7G8ML3mbekZ8NC+jfZWav2PUq4Ofay9c5sSOea0Numu8TV
3pD+2S4QMwBZGRRVd9MygfuqhBScFFa3ra1BSsiWicaniS502WfFvqhDG5xkOmJjAuT1GVehP36H
KfaG09QRvCfCQ4Z7uYhcx3yhs3DBwvuzRVn0SuQiT5n3rdah1KjKCgXFbk62L5gnnIycETx+ARDd
D+l39NIoD06f2KWM5fE+kOKjwQM/gtInpFJNgBm6XVkHpIrFAuYL7TFFtJE326QyLqyXr/v2eTyA
WCAuWHQ5VTu4KZ0WTKUUwBCWLQDzxNOvSkDUHFE6EUu/FwApstEam8GjtECRltgB/OxNZmhXAlZY
RFjUnL1Q765SLooAQugqLlSybqrAj/0fgbapsJEVwRn18r82eiWLAYjWkXFJWBP2gv9k5DRuWjof
bSB9Q7yyi+z43eggUhm8P7QY5EcbAGLEQeCji6/g4PADFTAHybhG2PK+pnqlMa9F60nO59UGK9sR
MlsWicxdg2oBv6o3yefHtEnR46CcZ/6SM3+u697MS7+Cx10fbFRpanFasdd68URnCVM2QSeHwsKZ
QkUa+Y/czEjp/15rLX4c0lioc/a/10EjaI0pB7WeKZ8FAHZzCiDPu42VqUqCoz8JoBPA+f4Wepb/
YF9IMS60XwMI/c/AXnm0QtnagFoY5VKIcUoNaamd/WLNu4jNrl/hzzOHuZd+dbVJe/gv4C5xrrBE
mzY3ziQDXGr7qFCkQe+FMmCpFdBzOSbGl5Ci2u6uSDxoM46MX8qTO8PdUGGoZVAuSLtjA9Ahimfc
qwPt3PX5pxwKUSYB0Ro5/yIa4O4hkWBkzuhyyJiN5BZLFfQkTdNmZxwUHef/EvdAt7zKpentddjQ
6CYDTxkpTeUx7iJLgsHSCQyw7CDvnnww09/eDxudLPYYjd6nMCnbu2F+7PVJoOUwQzH7k+uiAq+r
u2+giaiF/tIWsV+4Zgz6/P1U/+zYG2hqeqceqUwVe6U5F3mhHIISotctR26eWDPH+AbWBrLvohhI
85gtKXMW9VtkrMhpWSE3SgO/GHlui8E2Vi2ii0GX/k69jWGZZU612kmRMeTRm6puaqdxYCz9x1vs
BRmDqKbm9bruTqtB6cV4nc39N/YwMlizsjJtjjIpYH2U6Y6JB7OtaHyFDqvOp97QwWIH+dz5piXw
fPVEe/FP/JHmn+YMeXYvT5Kx/NraoO/G8sI8y4SFzzsfqzLu2k9xL4cikZC4GQFVfJYxqpBU08ml
lgq13PhvWaKskmMB2EsvNORrSyyqMyGnwFYrGVJcg+k4YDHuG6ceQsXvxxAHKl1xKT9xpsJ7FynU
AlN+ktV71O68pGxpLKQv4b45brGJcv2ZWmJ4LR5b4V6DLuyKay3jHR7sisXJ3c1XfP5oPRIgJmS7
fJBTe/LK2O6x2xHoGN6PPHyC/ooU5zE9YbLEOn5SgKQE8RG4dpotRO4CSVuSm/kNX2kkmabm0MkW
braBfuqWBu3ZC0pTb42/islubPaMEnSmD41n+pOv07CKkBdxhGXgPDcRwxKD7C1rKGWs4ngZcKPH
ztHC9lanRu0PFcchgzKzUsI0WvG923avk0YcRCFBTjdIKgc6ps++OMDTl4c2js4FZwlcqvSmp+bN
dLjffgEjQC9UBzP3kjIB+QccF8/3K18/SwnLIcqqAvm0d4OqyNzY5HN05pnXKXqhJ9TkLo370U+j
aO3DBr8ZS/UTbLpR1s7DpMfRHU67RxqWMaNtyJA25+utYVxRHMPmjF8bJJmkQSLS4f1y6qffWNPx
4ySwekZeC5khxxum46PdIT8Q/Jnq8pylwP7Uh7uUU1MIPI9AtXiU5IiOKiFZZcxmmDyBfcZegELX
/ECidzatUx/R/Wfe/0fge+dqB+Qm5hMg8yJVlZv6fiaFUi2Jzxv29y++ZDx59WIgLP10Y6FdO2mQ
e+sYBzE6KuLC8yTJEMb49dpuGAftckhsQZx8GXP2w3WNHfQvg9tGGNFE8nxqAD1LRTdEBK6TGg1Y
M0PUuDLoryy7LVLx03QUZGg3TD8lYOvqrPdeR67E1CbgbIrg96QAnh+JGNmrkOgi/rRMxiNTcLjt
3kKKA/trnuJvz1IPs+QzPgg2hCZW5oKXArRv9s8mpFmvLCtJ+EiAmE+9RqsnXW2MZrGtnYPfKcwO
iOV8tWIpDKzEVS545Q2lpQ+HRM2R5J6Yxj2CIf6b9WKpDmdEVxZTDFDwMCLe2a3B0XdfC04YgsFx
ZgkxQPOqpDx5qm+eDakjrZtTvgLwKc61XTNmCA5fl7w4kp9XRvlmDxiWOjP3r6pdXSplwd1D6r+k
Lxna8JOCVZWTJFLEsZJTI4jV1s0i3ISj3nkx+32cI3yKU6G7aUL92jXcD6c6CAFADuMv/x2olzAg
/5Hco+vQm7v/Xj1Au1lSBIWg3My3lH5qFwnCXCysncStahgP/rckZ97cyH9dOjSmJDHIbglw0eIM
2Z3yKZ8cHF3XJW8ioLJ1Hs8hIxjpcPu4TPTRxxWeTtYt3vH/Mtvh3kwVNp8oOESJt59xaSlEBS1T
m9IIderXi8ltrr9jUUFYHB4DJFjfQg3YhPyyVgnmw38/0hdcy8b/98SAzdiSs+1ctN31Ois+vsK4
sg65lh8ztejwRtvnOc3o9tuhVWF/PGhAIN1aCSdFz8K21FjXFW9Hu3NihlDiHT3aYfgs+BWJEkeO
LmX6KkAyVAqGZVLl+IeC9ZJUsX6eH1ZZy94zV00SxT0UVaX1rAsdk/RPUcxTVF7T86/D0EHC30Zo
C5ragJVG9/eMtmpGtOAaow/kSe4/6zb9Axp7ui1xG+IWKPkkEze9WVCSL+DyYTwnUu1VvkMsiFBz
27cXVChcIFNOwUXE88sI6e0trhk/xgum7GSs2t+eRMk1oUPIC80OcpbRNryKlGhp2cmGN7xan5/D
mGRL138bzDeXdyoLP1iGsqGB9qSvWS/Y/ouW0NGEpF9Yrqp9z7gEH5yW2i3JfFJLS9/fa9S6lqGP
t/RUpddva1TZDVnMSkvWrf9tJDIJhEkKZtaACcWq0mncs32fr8x7Y4aedxK3qEyjs0SJbKVHfajV
AlVyLcGgOXavwmTNnMCuerXX6GywlF6oET6CuK5NER/jxNbi5Qps+b4EscR9u1jYs8cQU/GCdP4a
9YkUIXlCm0DVLwirFbMuh2BSpGLPQI0sSsiwlkh0xjOFXM8bnhBgUySzWeYCuauyGvgKq3Hgkn0W
t7wvAglRd1SfSqglSl1T9gFG2np7QVnJdtFQGo+Qg0NTkyJaTPXb1lXdF0oWp2U1OIVFhkLqD10X
b3L3rtd7NuPwfv0KLvIRoMy8McVQVFuqQP4y3U+5Iu+D1oNez0N3YxxAfYGrx9wGVaJbK80+kBbR
4rns9kM3mrrZK4h0iU83xWYd4eWqtP565iy2zgATD7c6mhitZw3AdCpFtl+ezr04W4Mb6Uo+7NZL
R7IP7ChZ340v8Rfud7vkHR8OvwgPwo1E15qumsJ/yk3uKoRQUxVCcv7jmdiiSWq2RQs3jz/jclKC
S8mvDEppfCknZmusZdHakuERbpdhhawQeYimtmoRXges0ynMemtQVOOnuWvl5OlLBezc57YqbiUF
Bhv6tfcSO/xHTHkQ0LbdOKN4j1DXPcVdW4nrOC+bcgITmvZIALEWu9K1/RjkA99IaAcTQkKAf56L
4XmIHkS/2IWmQ/DtpkjtWAADSMsuVeq9BZrPfsAcxUvAKc7nxkOuqcsRSXrDeLaYOsTuWTpI3zq2
NWZso6ddpDMmB4Rx2874vT7HESGMG5G3NevLX536ZReKsmz9wMuYZ4XLw8a/U00qjCFxT3J1PbXj
Bnop4Jakof61TRmtaCcgTpLhvrULFBgKj3Urb6+cz4s93XBxTVWicdxfko1PWN6KNa4Luj1tue6s
P8ulRs1fpTDQ/JA/Rr/vRsQEyqVXdD/WCjf6P+tZGbc9p1K3PUro9nsdYjQ9B+yfd7mOz+mTLgo2
ZxN/X9VP+c36tuK5fxiNwikKYmXaNC25wIgHfzRMaWtle1B5mExJa+N31FWrCWRhNPCkf7boWC//
QdxqHcM0iqNezPVDUUNkgtAOtwfKcylFYbP7qGkrll1Qz5baQPEkGwhoRMesGfWL0eFVGmB0htI9
Jm/gWZhJc9mpvM4oHNNeYhUAp7IlLqXfGzfMnOMtsrsOXs1geEYGMNRqbSIvPeFhNbPHBtzGAAE6
wMqvfGFEDAy4VjNr/hFuwzY/51FtEWbnJ6CvLoOeW+7Gt4GWkXPh4f8FIzZVWopW8teXNVXZ/Bm6
tZ0rjqvLIwUuqQkceWbPP2u7P/2YWmLq3zYhbkDtVfqawuo6WgGbUed0ahKJcLIZc6na7OG8/rWo
bUleO+gA5KoimYJxbsoGpX6TQA/oJ55uv1WPjVwxxpUFOoFKhYsf8FeCSLzR+R3Vd8KjWf17t3uy
4kKfSFnj/H3l2tslOsZEbcpnctkof1o8/of2ZEScpqEVntEUsRLbR3i7OyF4QEHain2AHanAgRcl
/Jdjt+ejYC4mFJmMSEqdPao5sd7LpQFTKXosFRDPYRw3Fl4bpXwX/fn9OJCBFx3VcZYH3m7gn9/+
QDger9v+jvQrZMRQJFYYZzF/gHkP5V7bEjCYk1NU4hi42YoV+Am59WC85bUl4oU4l8jkicJK97D6
zU+6NIezyLTLoI1+5OLIcbSXbRO+gskv46umYpuNNA5fFSDj8UG+Q/xkBtp0NScUvYr5ihQYZffy
RKdQRe9S8Wl14PS3BNQP1Yi4SbbduGZ+vNtNKpbRU/6rHteoQBYGXYoJfvsuCGsgPqx1emrldwRo
JVbpPHyNn4z/8c4WluazVQ8Unf0jKrfdHXYNEFlmaJ7mgalu88F0Xyt5Ge6yF7A5Pm+va8cVty2A
AeXnc0wSODFr572NtwOxlmodOeljKNdEnXGZ8AcITf2X8Cw5LElquqoJwVWXZ9/TeYXESfc9I5mH
P3+6blb19WNLZ2eT2eweXQ/bye+XLNYRCd8lz2SAIQvDePdOXnwnvpIlJD2J4WxZPEfHbmtCWyqh
MX0VPQ7YAfBUhCK5Fd78vcQ=
`pragma protect end_protected
