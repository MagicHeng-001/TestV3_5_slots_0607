// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
gru55x3r60eM3JqyyeW6nQzXXd78GZTMjMNF58BimkcWUAfyC7o4kPMTAQbfqUcpb+djEExmnqdg
UnoDg5RqgzNCzy8RiuwFfIkvsKwTi3Dt8HXztzO4NmBWuUb3ykcmaeXxJF/IOurxDvpt9BC8Ov0o
x4zlj5be5RpLjyjlaD0XEqgGhEm5tl3ZSt5fchcu/AD/kXczKTOKNn9Tz6BKrRi0/Wa70okC9vzS
bWpZv9GOY+6ge1DYt/ZDY4W8rIJFbcfmHeXuNtlQx3FLb0KajpXODysw1PQWgHNjFzf3cWe4atpg
fX7Gly3DKY1wDlT4WAr/RY4JecXWmamLysJLZw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 90592)
yTlqf0aixyS5WtOhEAEzDJ9jbExbEk/3EA0H6+Um3y/Urjsw4wFX2nfhpDyzpZ4ETSnyKLRpDCDA
Eac/PGlwlnFKZ1bcZo8EyNCcgNrd+iuLcsdVlJmwO9AztRfgeYwq2mnp8MqItYrcr9MAnrwLCFs2
m6p4Y1N5zmGfdhtMKpvz4Vk3HSDybA5zQUl07kQd3J5kCZyc/747GFP5p5qgya3n1h2WNkdUHeHQ
4gu0SbVwlAqcZFEhIyjFUwM3YPpUP1InJaLHEZQSA7fHIiZM5qkN2nkVIPLO7/7BL9i6NQrFNT47
dI25HdnwUNh1Jp6Yuct/Qo2KHDFONBMUvx7l8MHvHg84UMGgQusbMB/XjMdkisqKfBOpgn72Blm7
FBTQ4OXhICQHT4Yz7/9OdGhMU6CSa3H3M5TSum2uuM3YMKxtSZDowRZkdCtuVLLdAbjTJ/P+gacx
o2BacPKeA6t9x3EK1ySZ94s7OzpMLr/ICWvx8Jq+g7JT9cLzfmLvoPnhAExd3NtBy6BSCWD8cZVm
THGcgRdgay0ub69R2LsQH6eemcZkXbf18wmv2xmDW6Truod5B9NQFH5XG8Xmr3R+DIDDgZ/Bo+A/
a44mtWIZpax2OEztzT0I24FBzHRMCBDwWE362UJ+Odec44bZ9PEWvLuaEECEt+l7SpePamzT+eH/
DB7qvKFqUMdF1JLKpa63gFcMqBBAgM0nfw0iHyLCZtMBEzNzgeTnNcU04Re+eFmPNpZv/kiIqYou
De0rErzEn0h5u0s8L2nQ5dDNk/M5NPApUKk1Rq6k1rtIFXYXys5wpJ3Xb2EYiPcwR2xWc9rjcLaA
rP4bzyoqVXlQxdIFNn2CdrF6Y412OuOnNmOk8/PXUMGa0rfRlolZQ/2ERYPPLAd65I/vmUkknkNK
lRtMGLn4R7c9aVDiuGHKoCnH07Yvwj0up/b1pKGVgKOg7GSS+z95vlNgsWyLXlFoIFsOTcjaL2fP
JSacgclIfpf38rB7T3heGDuejDKNO2e5r2Nc4YmKSKdyzCwHrUWbhYF6REf5ip2fBmuBXoJjgdUG
053ZMjOkLtrIfrfDbk4EYjyvc//GDJ6hQY37x1VDCnnmdTJXmeBAiEHtYKiF8W4WmMEXJ7jJGI0J
ai72QUgT8/GOBiOR3zA0AFpGbZwbeEkFon0OQbie1lB5LJq7bw3LJ0coTjfhjlpkKpS+0x8pzbKh
d/dcmd/Nhpib9ZBTq1LaRtmZLIv6BEK1mVZhpSUMTG++FsPn50qDh129bvGZmZsgygidIfG2wsDP
SPjA9abjM3HWSiHNqRc8o7O8KGexUEjNeRX/vKP2eUb58H7TAaNFnNzCyBfaEZv/pdvQuY4PyzHl
PyO72bdcCK+PPE4QY1AuJb54hNybvpVZnBkacj00PgLg3AZ5M2HEgppBE64eTRP0r+X09Sn82VAL
UwNINGK9PVsWh+sO5FZ7xuYFs8u4uSD/OnDXMJisbLuW3LQGln6+ItqTLp7yJhnPNCo5UbHDpTcW
PESQE0cXceTf1DocsDZ+1GL7APfjcCziDnnxLQ0sX4sQvUTtaazGrLeZenu+ddCthgYSbI35nqyN
/fgYZ/eoWEkbDC9CRc1S2CuocGU3y/MPfH03rwL461QKfI1T3qt0umk0ldnZ157kjl7K9CcBT4mS
izpLy2QcFducxITL3wqwpbxZNDpBJ7ZwZaDXDULo7PGWUO4czoI6YT7DG4jRSgPgfyDsEYP9Wpys
h+V23C3sS0nTDUNGmqnMxrgkW4aCngNdziucW/6rlBk5rrccRp2cNTeU5cU+42pYzrV6Yul9JFqt
DDUZjnkwHjFpKC5bEsVQgI2Ui4cYiVRE+kDrGsge5yQ/mje6ck8sR+xbWtpP5rdgnhHtu9I/pyLQ
ntL7lUwYWbM6FM4vFPPQD1TdExlCWy58ht4DHT8phor1ykHbcxwsbNU21xKHJ+UAoFXW3N70vmpx
jM+us5TsC6VRv99TuFnRAkzBrgf38lwyIo28/AMycFPKHon/rZ7gxgYzwZnLwE256cYHAGsSUhxU
Q+NAfbPQAPPvnBegHav38oKYKUNN18Df03YKkZCZAvG4yNcZZJiGWlMywd+QRXo1QYrKV47LTnSh
LMF9GGXH63iqSVGsl5VNOmgmKzhvQvYzvL+8YbP4NUS9eW0XHm2Pxvs/E14sTWhFkpbGz94C9cgX
32wmiD4yTaN7/QPUx2Yik6xx0Kyt/et0Gehi3g3v5LpnDnp5FgxWYiN0ejvf0jey1iYvKuXqDij1
LJjfsqmJgXH40cXyeMnmWULWwvwzpAshUEfBX8UGgUGbck0zFqURsjnZi0QLLwUy72yJnmCzL2t4
UAFUAHZaaLI5Kklib6EaYbDb9U/YpAo9Ot8NGTKsLymrWStUS6i7yA6sWLJR7fgJUv+OLTKyWqtk
NVLrHS++bMTwVZvSIp+061fls9P9V+E6RztQ9s7Y0NdqqkE0e7xp5dG1t5VsRJXo3Ycyk7TG7GBx
/xG0Vfsq9am7EulS6OzKVvA3hNlb3C8WDNQWOr8XzuwpjXXiU5otiGa42Y2adkTZXmQfbpWqTxQ6
NFjmszNeTLkpYydU6VgQhllN57GnyobrZSQVzfLmxwovXnFzJSiT28DcMqezevxeSTmQ3bmFrogJ
2745J8n30EbbcDWnma7pX5rklImVKrxuE8GVwUHnzjHa22jai7Cxh2G+DPWDExgq8xowWUUz2b6G
dDdfP1Mz4c05sdcmdb3ODWvJY0Z1DidjFV97pptD8emL67CfU947qw1ukHcog9XCMoRalh4Rbzv4
DnB/1aF/rgknOqeGASha2YZft+0XgBy1YtlHis/IBV8RmII46vfURkdZbgdHQv7CIRBP1AcSpFxY
RnDiA7/cEWdIxG5DL13jv2V8pOurAIM086YkBs1OfjSisVVkXPvDHTbIoid0rHbsM3Llzwzc4dPu
2cBu6L1laivcB5FsvoHi7ayq7mBP4x8HUjdTVtA6rphfnKwwVumL1qIpNYpNw1Np2t0NqZO2T+ck
hw33NuduIxI7UnuAAzZrp3ZvyuNv1y8IG+xolvZulN0x7ajZD5WJm1A3TVvl0W6f5PEyuhUbrXDf
hzLtAD8DKyiitlPNT4LbJVlxpoatHqezCaqHM5vOZM59eSvZq0aAbcCAM4jorAnofIz4pioZAFnf
/Fa9gkBnS/V8WrU2FhEw5HHftvmJp4kYxWWa+RlEbTvP9c/HjDN4AKJ8HR48YnujqnDCH2UcvLQN
YlLe5ZmhgCp+0nSVHSpmf61wGKbnzRCIUQfAD5naC0yh6REmQzqt1rCXHBWi2JX8wjzcN5sTelEa
w20kJsc/ss3VOP0MGJQanQ8olZBNe1D1/LgHCLaCdXxZp0hPBLeRKPFkcCFCN6M+g9og+nFK6nFX
vWIZ05+ZV1VdCWM1vlu3lD1m/UrLeH4/RE4gR4cRdt6sIqC+4kfQz9OA/VOhLmvKY1d5Zl3ov6CG
xcxl7g8n/GoIp7lbJ2u1IPbs8jdhI9KbspHTdSc4j5XjkOXSAQLVb7a5g4XYfOfeh36kuW3UVxvK
7qx//ou8WgNkm8M/4h5j2m4dXiztEkTV8Maknszpi01+N7SIX/0OTw3G3MRBcAj1ht9AikTatAd9
slPxsjd8rZB+pxmdyzZ6cPSJAdMuED2FQbmce7aBqhvqTR4y5Xpb3fObRw9/giFbU4QkWieOf8jt
IYh/Mhd8Qe6X8FweUjqAP+aW8rWwiprHYJfRnp+e65nIgraDqOce0RVLVNYYsPSq9GVb/l3kgo8+
1xaFrnQ0el6y+xZnp4Z4/4QUDNR68d++d04QizMfC6pVGuiPlsZdKrBdd96ooKhlMkBSOpQNpYVp
VKM4qsVNflJSm2fXPDc0VnB2jtV1jH+TqRHzT9hipTD5ABeMh1UGGXKIiHulnZuHk3qe/WKT8yoS
zRpMsDEC4yiXXTfJUgB8vSiN5SN35E9/VWJsfbNhuVIJg9+M3mE2S+SR7++J0NyuvcngwDAnxyaa
jCb+WZ9GC6QGNL54WDMnlxH0Lwpy7wzR8GgOOl/JwVeQGAOIGSReIX87xQotI3+DkGnFX83UqejD
a5y4w2HJ0VU1N5PNrYtEVZ8ZsM1/fjQSGx/iiQxmUIle//0+Zt1ko12p9AfMji4dmQu/GqJqfOmz
2iPmN09K3Zb1G2muriFeKPBsBQaE0VftaJbETSdYt3q/8ajMyxlpXa6fZu8dRkJHyETGAi/t1QsK
uqsbDEGzYy5UCIjdFv0rjuicT2UNnM5De/CSjI1g51o8Z8QeD8FKn2M3hGGUWLRT4WfuwjKI/o4J
UPO8+b6kB+kj2CRpLkQO7KYykumT9x9pGRV6mA+zwM0rwtMj490eIVGE4XJQiJwqUQnA8rkuabpw
DvvRUOmuc+sWkXVDInuLFFOeZ6esrLPnTZjdQKAQLZjtnLoM3VKEBia+o5FhbSGv/y6oSdut6FBf
CCRm8o7chHRSKqhUmHeGI4mCS0i0NDZhzfO6ZuCWy24aV9bKFQUDxwaUTW9LVOQ8s0nTwdCekP6C
VoBVoEuCXkyIn1YhStL9BM6ZI7EnI+xvl0G7HidNt1GRswgC8UC5XUlwn8HRS80723Q8EWO2+9+2
UQPIqWoLpwr6MXAQliqrXwjC12aYTmN7WjaFePjjNgkJ7gClovI2G508mlCmHxpvrxmTmBM3794M
2nxipqPr26nigFnF1IS4CkMExpUXE7HQyi+xhLiUSalHjfsz/03SaqauHlLnn5VCy+RVG31KQ+ge
1RoAHcmAOBGJf8e0pNtZyZoOivvkCVDSMixxC7dofqUd28YPjZ5nD4mXnImoOZw+k/nZeCO25hS+
5FOvSZ5/R0QdD5UUlw0maJPWMqYWm8we+HRHgk2MJbbezKSgK09wlFeEYNoE6x+TcHqyxTi7rUqM
ldI7LNudGKzi414/y0/NZqJCAf1gkYW723XfiUdFsrOJwihdZrp09BlZCZU3Vwcv3jeOVvSyVXXN
pmPhumwJ7VrLiqn9DHWlp43gQ7vU5NtQSNzgxiqBaWXTan7SiE1omVAI3hPoXP09Yt+2fk0Cjpbc
Mr80KUZamHOsizPTOXtmw6Tilecx390jeBDBxiuCXBLlKd+9Nmn2Xnorm2GWeYYqbZvHr7KOnGcQ
i85HXwCQzJ7Cxte9ktCy80JLvtqvQcXIRVu917/kxHoUKVPrHxXW6RtUtSdH26S5/T83zCt7BJRA
OgGT7/5B6OnjTwH8pu3UeOoPooAa1fqwZ9S9bYJna0gL85SCTJSn4YPiOsOmEpOZ9NFodOiIOfpw
RmpROEppt5gshrzhGiYtLZwfeXJn21cplBaYL6+/47ZVgIAxK4GCJaNAV9kRwamxXKt278QkhtfL
THfkgQOFUrQP2MiYx/YVjve+Ht6eOoyjylwdyHWWnUhR5pDjyMXPgvhRtsUWUW1L+fNvAcH29ynC
LpJeMtUXOASvzOVfxhL+qp9xaWbEEhEAe8/KLUpl6gpvinnkzhgN47Eqb5xhG7RLdNLv6hXWA9jb
i9jyGWkXzjFFKarWrNoyzB30RM/ZsRp9aTFpIHwTX7DNR2oYxB4wozOGtZSmVAkqMQZqvC/tiQA7
RvtvbISVldVIhuU22XWsAju3OY9rlStJyGvDJH6JkNSlX86CfwmGV6WRwYKSE3nfJ2fqscqeCPoY
kmeM1Y0ty1I5WWzLYAxrV5HJkOnFrqpaRE6daRqZGh4knCHNYJKTMEW3xnf3W25y0/wUw0j93ZJX
SkLvaRz/vbHFUHEr1o+mzmoM1TWkWSqapV0mRHR1QY9d3a8n/jydU82JSt1o+uFAlvKeWysjDEZi
tOE7GyxfCSkHR427TTRbpD/enqsn6Mw1omrWPhRuImxOWxdZCLHwuf+1z9kpmMPGxpHqlJWHzXgf
TQJOcLoJH4FP7hI6wFtwRBXS7q9jUecfqmNBuvJPfgC1sQOvBae5mDxdTGf2HAwniXZo8Mz573FP
pRZWQCeZteca2fUNlGkYZ4Kqrd+34QivSr/tNOxohtmT2nnL93/AL7rTMAjw+OwV0YRzrnQWxku4
QipvOEHY9Eg848AklDAJNQOG0KA0H2EQti3oQ7xBNT9JfIqTgvru9s7LGXgPD4iUGcLF5nXTR8Rq
pNNYlTJn19czCLJ1RdW56hNkdFaNY2JMejyn8GPlZI6aMkKPxVgXTPxEqPYdDHaR4AV3O0fb2xuX
OGB5Qtbm73exGEi+C0G039AVE+6zL2MC3hsRu3zCQMjRdF51df26zz8lBLm+XeTeHXg8JQh1WrUh
hs6W+GgW0aqoxbuEq7yYDWE0+fg522ik6Yq5SfFeAnTKJcNeSf7aqX85+bnYZ5inNbysmaiwndbC
7ZNhFncUEQX/nCY2dxwJRcCJEzAgDS3B8ezfRRI7cCGys1/MMzXjmVBnEoVRhjeTSekpTFreokQX
cJhozg86u9d7QQ26GA29LI10XOmYG6gjLn59k82AVL+IXOZzAL7LfzPfmjaOedS7yzYOlOBKBjn2
V+lMmyZ1EdKu2Kl0X85fdQL2bUqq5lFrlfPazTg0Yyg3EQoy/N5+D/mbqSjirP9HtG0eWgNN00Gf
98ghhS3EwHEaVLt4/WD7kpu4b7G0wIp03MeEsB+/FpIw/GnnZuC+KLt2cScpIziQp3s5GTNjJw3i
ns0WOl18wAnypOI4DaJ+/gE+pM+Y0YRNTTLPkR91huUzj13HYt6xWgKo6PBY55ZvDp7AhTvuK8Ss
zqBqtpGif3XxraRUepiNQjp7ivMQykCXXl4UZhm8B52zisEhMViGdZ9JcqgwiTVkAnGGVkGCrxk6
Hw69mIPHC87Pl+Mmj9o2uqKmd7B8ssujerlaiMXEP6Pkn8xiayN6Tb0Hn9AMQElXdp4PpDkXTEp9
jdmY3i2Vl5z6ei5Z1HzjPg3jrUJASugjhD+XebhXasnhY7Vt6NgrTaW8Vidn1pvAgX3DWoH55Olq
wIffloNTfjiw5oOFqlf4nc8hPAFgbyiro9zlrE7foGg/91ggukqxcx3K4f6OPXffqocu3SqRoW09
6D9BSPoJkK36DJjG2MvhLPaUqFCjnFvrqd/FzNiwnHeNvzxcm3wEcQugd7Hwso6rchM1OSGX6lrr
rLdsR9khvH4d3uaggidJHhc355bdpYPK9eeNv4GFjFVwTVGKr+Cobd4MubE7ByINzqm2Xa7dWcPY
8w94XqKJkt5CxKS0IMWh8Wg0feA1fmD5gtn2MPoIrKAje8Jkyflcp68f2+XAB186dC0dCqU5Chtp
u6z1Mwq/NS4W0qHNbbDUX7vN5sLRmSvd0Vg84a7F/ztZ0JzwRfGexmdkYGXBnp7JS7nNNJ7qHC9m
JNyWkxQREUPCVHkVKv6MD31lh+dL3NDxhBj8ppyg5NVFhprnSeoa3Hta9NqKgSUOxWlXY6POQgUh
2htsPda2X5ZEy+3I2fVyscm7qtr4rzDA5ee61JsJjkidWVEN6XnQXgiXZM9Yij7nMNc+ri3s1lOu
RzEoXypHMsjsIurDNHCPJv79N0yBH7jA5MQ0M+l0QqWeVLixnZQ6UErluK/HuiUvuvTe2K3Befsf
PbYq22CLYFgDtln/dXCMhMPb4FVetdcryuhqkgKl6h1Ca5iPAndg1drNZmRh9ueRwx2Ailkzzs6z
KdQH0Vedfqpu67bv4c8ow9+lnxqt0iR8MfaeBvwYrqrmuylulBqrhAsBdqGwSPP0q+w+9gB7NFvq
gD47nSxhsWF7iQ8Zdcj11GbAmN5nx/HRh2pgQHJM/UWzb9vRn3SdLwX35dmf9jEadqP/Yp2sLY5s
JvyjNZYH5mGzWA+7sWqZzD7ZaWb2Nh1T2tJxyOry6X8LpnykBFLisQauMdUut5mJnx8GhnW6LoUo
q4gOFSyBQHWI9pWseRQeaKF3YVzuaTc18fnp8Pmopymj8BER04Xg0UCQSlyw/p0ofPdkbzDAu8/+
FRjaw1Xbsd5sRX+bVltyc7t5U8K831hmK5O2Ty5CNTor7+KEUlu1lB5lBZvWekp7LbqXeUxBnqRP
ZcaI5e6EZbBOgKAO7a2vxp5D61uigZDyfX/yqiHY9+SelwlVqUy8Fj+AIUMzSfOSBFKrR3HjIXrG
9bjWtq5/KeX4MsSEJWXM8BjVn7KPgYAb8enDl74FZcYNpDc9hevX543EHxuPNsc6ycAqQ11xgNLB
j+98hzt6fRkf1oVs4Izb60EupwSLuhPMTPV+BHDPeGZK3oACSYgvkgDh4JYMUs3frDm20CJbhm3k
Vs2m7BKRjRxxNGypoJb7TnqDlg3EGzuRGC/aIjRScx3392+AM9RHrhJoV7inTcg4hgxaL/d9Bd6I
X0npH3kAOZHTpwBXSDhkmiCE94ml7ZpSXaUBEhZ9IBVu9k6EygSk5EH6UhIHbKVUAWCXyToxhwj4
myLw097LzlO6cheFziI5wSPOH1TRq0l5GT3F+x00JEMLLpHrcrdYaHpNjnGdQot55p+3hHgBuV4U
kIx4Hp4xL1aAnwQ4SZYeB9eX/J0PHZtlFulbn+04IN5vc2DEcBZkE7r9LISuOLBHz78PNl+QGlBE
U5d0T4jY0aYWPR0IBPW+VFcA9DlBc24e1JnuW3lPiYnStqb9QWtUNn0i2GIy4YuytyVbYu0HmuZ9
T7LWFTfrC9zLY1KVlcjthxrgoq+LHLCBmKY7VP+nVbV3jC1HGyUuZg9gyXEPRdAr5GJxnK/YBRvN
DMohNcifl/T/sw0/U6f9WmbcOaaQMD3lRxTZYWD1akQIlN9UPKWtu1dsR6fIm7x8SvahWTE1EHq/
SUqNxCUgnfZ1xE1PHrfvEnsOC/GspjGeZ0n3fLfl24wLovjUPl0EF/+c3sjVA2U5imQ/bzmyryUB
mvSp/Uyv6bv1YYmjP3b0QKe1zQeB2WmWp/6K3Ge7p0hDwmpJw3ird7fEUK6beQJKQ2CLU3Gal7DP
yK/25h+biWIhs+1Ia4yo2cNnTSlghuPGfimSwuiTf16RxxFEd8r5Ar2U+h5QXC7vydoHUZVTTimy
eOrMvM2Yc7Ei1MIz5C+TDz7HQ98I9YGod2uyjI6xCJ1PF8GAMaDW18tSEl+uQ5GNSmSM58A3ibwS
UegCZiSi49pbrJodKefiBVWLrBKvKPPHFE95Ox4htHZH2kP+A+TYGt8X5ay3eo/tw9UjawFIlluD
tQeMI1fl/e/7okB0+2mKP0uhwjmg+lE3WZ9VCVe1ESIUx29FU8lv6RcP2UnCP+0ESbWTV90Xh12F
n28RiPJMqBERAd5jNfl9ua5EgPH35AK7XtCQFhlbLvUPJG4qoCSWcvLhA7OWdro8U9nWO4PaziO+
3oVOpfUDtENztm5GSx3raIl5+FqfFO54RI+YDHbz1Pm8T9VuI9TH6GvUl0Vc4DPfWxpQrloUm3IJ
MRGHE3MhB1hc1+ZWhonG77pBvRNSwuca3jRvZ8VFsknkn7j2+MiAmloGXbAWSpJWAlLDvXwa6ZfQ
GjtO8S0GsBNy2ZrJuig0Pjvo6+eJNWfEi+m0mYyX+nMFBWLH7dCiM4vsCFnWOAcTyb1HGckvJu9A
N58dQkdtr43FJNMLEpf1OIplK8I7UcM9F0exzo32YzVYE4RCPc42XTKvhWZmdmhOiEiZMgaaX2Ae
FgdjzBHELRiIMbj4LgQ7XrEFrJe98fs8WT0Avn9Vj2BSRIpRz/JnYHCDS6P/iPnvjZvip0QcKSEK
S0x3MDWuEwPtByv4XtBeyEYL54C5DxKhyB4c7os8yFNCu9tMtnALoAV9tjSaskEDivurlQkHDXZ4
+HHe7F+O01+79feM9CrcaGLIo992Ft6KqB67cB9xtgwSY/+oG1649oFB9ZnUH/PqGXoEDV2LRl+e
SLlgeVeJOcrDkNPGy5GgkMAdzBJptL9gNCvaLkLBv+vJN55lLOJpfgaL2YJPba74YMBNHyKGPzc1
iknMk/ZDjeFS1szgxuIrniGQ5AqbKjaEEdPWOKMzDu6n7tP7HNa9O6hUqw7Lw+SjTxz+Fta7aM42
cEUAz9RATOdA13gupMOsCiAG08m0tStLeiyLTjisl+lUtHXXDn7z2PfH0ag45hVuo1+qI+dpiLVn
KsCn+qHF+t39BnBBnD6h2cvNqYt7q2x7PBL8XPPkgcBKU6io/w+gZvJMesR2Jt8hjjOQ74EEjwzU
2ODCnHxmvtOFwdovmV0LqGylpq1l9JwGBJusXhRFqLYz6II3+jvxjiEk8XSV7W/dDm/lict+IesJ
5YDQz+psIOB+hEZTPdNRy+6pcsgBuItLVX2slX2X1iIRPf8BB4c+1iTG3pdrprqFRD1gAae0d+pj
j/ErwCgK2UcqI6lXWMBXS7I/lDPFxJR7i1TlcIbE5kTlZ3nUASx9mFWKunWp9Ny4uImZaKmwKCPF
/KZfCNmD10eZTALAk/Z/So6iazVpnoKtrdMzFnOKTD2SH+kx8U756NOZ6PfXQcrD3o99dYF24rRx
QVf0OzJ7euo94F/27wI1ybpDZVpR1O0++KOhOgFME3ovo8rH024cW2NX466ycQKjqu8R5imF0bwD
GTLUfrHW1ZIa8y5IkY6pecLF+7KN719Wz0IPMI4UkPMUthqSZpjJfspMAwnUBYiW4j6P0U8YzPG5
yRcmPfKyLNjymAg8KlF3bvKeJGsgDZDdxA/ge+im3HnfKC014RAwEfirO++qtCXwpXTMkDvl8I1K
kVlzxP1VGEpXGIas8JtIN0DAngWxvVlU10ww2oISzj1yBTA2hJfJjyLVV/llKlVZPhCqSqwdRjuK
Z5W6NoaT2NfPpzA0iXybGiHRR+rlrrNy7A3t5Z9V419PHrz0WbmJ1Sda5XfodMfBuADqKKLx3vw1
WE/O1NTcQd1NrVSYtna8FMpIDiHUVI+Ouk4Jb+LDlw5z8BSUbt6P4EYvwtPcgirTCDY0MxJs6R9V
A6NtHZONkpKSqRtroa8YgAVKvoj/C3VLjCYz3kWOqIQJoiDnnxr9EgbjSEhM89USAHfSQZJKKeag
ejnlqURjzDrX76qsTtcYQXy3zyxFu1azaLb74DWIYNhLyrLjKaXRQcBqMCxK5IrLg6Ejh2ha2oos
Eew1xk8PLwc/Aa0yuAhOkhCxdcwetRv7nOY7d2FaeOLGoWxghcTGunAgWNMCXpHsA1/A6wPqIv8D
25J0w5KxJbm0SlBUtwILBC1yCi1Z6EHiqdKZf4kD455dHRNp1NKkxb0tYblZSgPl5IMgQYHX2Iht
LtdDyiobdtBYt+P0GD0eaZdc4ItyEzGTNZOpNTTQPVBrr2rmW17WYJ5Cdw/ZSQ5jURaq6U2tCn2f
T0YMExJV6YrU9JjdjHFqrLMf26JybeRkkZ0xzSQ66+j2UPIEUCi/PYyhtO17QXXI9FsiFBt1XV5M
qbbwKL2PafaMT2Y/MOLn9XBQTcA3+x+RmdjteSCqSEaV0wCsrNi0wt/9Icz6cCPUkR4uhr4Aovrp
MGYOnscBHprc5fG1U9M5WoE9I6Owf6dAugVC2xCrRChGfaPf8IsaysbJUAbEOgu1uWouRhMS6dw3
SWa+M2DS4O+fOjZg4v1jT4YfY30qevTjdbg7uZQOu4EDXzEiIgLggY74uCAYomO9++3rtrNjQdv/
A80lKJlGhodmVsrsv3cdZTvSNByl/QopoV6bi1JPIXePfC3iM+Py/fslV60R7tv7G5ktV2+89eRU
H4aWWL1DKKSajx+hH4x4Jx072Exc2XSPSDQJnoejvl4Uxwo56DOwc+Cz1opNn+jxljzwkjSB6okp
GlT+bgxrFEv/dxJyRtdvcVzm0lSF8INWTys6OzAmwUzsS/jBugGFvEBtTYhKdNztzVe3m/eCUk3m
oJWqi5/l4juY6hxP1D18NLGvz38EEhONwZjuKoeNUcxo+BV6mkFl64NEvDhIMPaIc9geAyQaebyZ
XrGkzFNzLX0H4Ohj0y9tJOUEShzEw1W51tGnsImwVYX50hO29kK1T0TnzkJrSTYsseZJJ0/PoMOR
6pyMSRpikS2DPAlizdNRqTd8LnLmN/VJDbv/+DcH9nx3eCyAshrbw43tcT/KvOj3dgtUBJNVYLPK
VGNTmSQLRRT1movwc5gd6qCeKmPOqn03aQHt/6yXCPPI/qjGiiCg7cnNDr++JaGdGpfrsmxcglWQ
SnMGCyLAro6Z1ItAt/TUoj1EeTl4+vVqHwhqHxLX/5Huzoo2xCwbAK/58Ssbef3d1u8J0ttBO1N1
toGQVgGr9bdb+hwBA5b2mmxCYhKim3mwaomPSHxX0zcDfG/A7J73FAwIgMDiKdWHQnfINwvNrxEp
xxO7Zb/A/VYlSGD7wMAbOBiBaieoUqckh1zu/Z2QD3s7v+xxJU00Sm4b/HRJ3DvmJonD7fcJIELy
3vDqeU+kVQiYTjd/M80pVOFo0VF7D/9sAgMAqTmmTAvjI7xZuVRMm44oXSNQwN95w+a8vLLPZhvv
/mf16lzrirH1D5Re5ZB496cZRhS3zmnKuZD24QDqzdkcY+wk/0CwmmHNU4yJiax2zL989OLiaGSe
klOFcgpoZbswMtviqI7hp9Lvr7n/w1BvW7G+Po2osf7+tyyLH9GgEol794BtUVlDzpvhj4FPWL/I
4xy0tJLUp0PzzVLGoDFgZB7p570OQDOrk/MLuLXsmCc1rx2vYVBf+l81G4JETTyL80HG6Fz4hHyU
EmIXxE2k/IQki+Nkgp3bWnOlk6vVxfTV8lBEgv6KKTpPTj3lTNGq6Dv+jf0LShNVtuW5BMor0r5i
zd6WH5kmYL4PCT8BL96tdUA9KJF6jkohwWUGP+BFpU5pklPE9V7gx00X0YeFVcv6ovCIpYaL3pkN
LiCHt6/vYX9hjDUvUpofS1zHrTVJC6LzALomintpsBVwUeSg5f1efC55W/UVtiKpdG9hCee3EdZs
2Jrqxk9XirLeO7HPkRB+Gugs2sQGc2wzdB7PcMhtBmMnTCwRbY9VOz0BBRnh9quBg2wnmGwQthuN
oKc0uAO8s9BcH++71NzqIge+u/d6o4ra+4DdPRywsUhKhhYpSvg84kEQ1lEPV47v1JchuAA1lZh5
pvh2wvIy+x+mlcIqrAVCvc92kSpS6Rt8yzVM1gp5dRZUvE3an0vlFY2XE5QShYNX5FALV8gMcF9Y
r88N/X4UYYzgZIGAmBAZNPimYvXXkUA4AI2Ei72eFJEVVlkK2BPlSdtieIXIJyHFR9HasfvDl9Qi
fXo8pmA/Om6RVKIjydKLH+L/KhWC4LkRVhhfYRDJJULTu1A1yJrmo/z5vs3ydcIBM9P9s3dlunKK
snMVp77a1wO9iWQxnwMJF/2WsLqH6jxCFNblonNEaURYQ7A6OEovQNZEuGDoYBk6w9RZP7xTmruw
S8mr9Db6zloChJQ/Y5jSHaStiTeBdVf9e6PhjfiCHXa6dGGFvLRiyVRjkUfoyI/5O9JUh6YKBeU6
9XHLHJkoRZ6n5K9OHTGzbEPZVtSrHCwrBiUHX9eaNq8HE0gnCGt1FtbU0cqEGGBjrrK0JAx/k2bW
0IEkiVPQ4e2a9oT21ohdYDcYuxWwglUe5A5kSuY+G000WWaH2SxlXYtlQRsm+28vXT9uz0EzW/MJ
Kw8ME9EOkVNxR6cPalI09/s7X1nHI+XuTZDSjhh9dR2y3EBoHciZxs5+EwoId1Lp6EBgkgocuY/a
iN0ae4FajL5DMDnJEVAM1l9w6IG72cehbqjx8x8bA5SvkY7v5SKQTaFazol6sdrZTMYt+t2kDdiV
IaK4VTCteUjSKtMvov82HYWO+W8ulqpvAWhddmCS8atkO3BUKqdpt5MauLzw3RUVPEH2wgrQOBCq
vyKocEMmTnnoBkJjU2K5f7428lSuj8uFzxbU7u/DPTSAOLRGeEHcZSLJ1/Ns4RnJuY8iIrq0wMcr
tZBjSqjsFesOPdG8D2atD6VpzIA+9T/HjOVLHXiLyv3/ZJkkjVwaP47jgw7trAxeU3KRIw2AB9ad
XeGtbfU3rvQiE+uCkhduaT7gcMNslUfqdTqelv4/J4ha6k0s4XKIg+S/9L+m+iCvwfs3AnXzPfh8
I2BHnJ6Jk1Uxm+u616RWIi6bEMIdACc9xjgQeDsq9qVgZ2qgVy1brdE5i5HBJX2xHG/It3n2WSFe
onZPnSEooRKSt+lB3DlnvQktJGEFZ2t9wVvCkHv4M4XEtrHuKU/f3hqLt9lZr/nf3LoJDUHx4zFX
h6aGdbuM9u1bl31xwpkhuZQGC4NSKOmPwBL7MJy1exNTnUVVMoD0cJSKuEINzXJ219wNg+6tRNM+
uWPxEX2ifuOoWS5v55WVaFzDn/5NUsmQwBcX7EGPmrBsR6jirpq9O25oegAbcbb/ekv+rMeTDeYU
ELFaIDM57g+UfCy9ZvPdRehoN8dbleca/S3xUl7wF95vqHalNEUn2jRQODrqg4DNYemexCKcmUsN
s+qtp9wmUQdB2vIX/HZMEbh55Vvg7OIMJSVai9DYneF0aK+5jTPjrlLBYhAJDMZQGu7EcxZt8z+f
2Kq2JjDSG23p7UYmjY/syu+bwCSgYAZ2u5rXe0M7hDnpUm9j4D+FUGTwT1GDE3w2ybJYFPTGgR3B
PdD33xX60I8hFHyXGXPvD7KcFmLPGL2R5hBE1aFLnZ4vbTSe+52qhjNThcMwFTkS0PlVJdudbWfL
OVEcZ2wU/f7zfuh4AjJ21mwp9CusAiSjxuoUZKwlbXa350gyFofAVYqZhHD5oxzXQNc2IxFbiyLN
WcqUwYYT+GCLzXYCc4Ohfo4kDZ4eC1JSD5tHRyCMurIR+Y6HQGNuUz2Q7pu5l1vxbPM1sw/mdcgb
br7HqVNIZk63CjeZQgnws3CBxkbss4XcgfL4SHQLOALsZ8QkD/KpJr66HpsPVNkGRieNUXHs49zK
vFl5pU5N9XOiNnv89BNhValSc00WX9rpZKHVF9nRvAyA8S28tpiaSS1fX6hhC1m73ZSizM+maSHA
eqKnUjrs9j8J+VnrbFextfBf6XD0Ne2oEkZP+xILUOetnV2yXB2vZwpHpxAGyfSDs8jTyRVmdWKb
lXeVI7ctdTcPGcswTMvlfewNukZ2RPZMWTXEbRNXMNXsQqaLSU3HY5h6KqWTllqiP2Kz/MN5IsNP
lGPx9PUIjOt/GJBn0OsGjqyI53Nax1O6lNKw8wjN/V177wtHXcL0kNE4b4Q1KCJSgxXfWybru4Nq
tSviF1Af4e2Y0dffyGtS3SmI5y+Fmje5QkeuEaO+uXmMewkMeysltf/ziNzx0Fp+EIrU92ZKq1A9
AW6VUqfBz9ks6ohoQA4xBrx28YfpG2pjKDBd0OGRggmW0Im8QaVkllGu5SYblbY4uTNMWahZ4UPq
mOfzZ5Q45ISxlf5U/7AZe8ko88++2wld4E/Ib+Iq/TkAr6hgr5EZstVEbviMXtpWmmLt5eY1Lc32
/alR5ItklQC066ux6mDei4LZvbWN+cCqmc1QDGPlIj0/SCwTUKMAcfRccIhbOuG3QFI/MVBQh0FD
QcqdpCvKdo0WQ7h7zpySPTp3BCkucUx3iWXVqaXzyrE6sBHjM6o78mXCTC49fMg/tMLyQEHe9k6F
cHDWc2XPJXP2P/IARduO4wrmW6bFPiQNnnmgV7vX/DvXT5YrXGjS9brvtB44AKXtRDdG1fAnKjd1
qodzLwJ2ghQ7SHTNCpgN+07yLd0FdDQ9hhB7G2xgQePPC1PnY7rnzJTvtkbZeop9s+HUAobRo7sD
0D0LVbq9kZRbTcOUoYKjaraO+uxqceVGfOpJ14rAOJKO69cUEfbUa2sRnIM4oOKsv3OD66KyGob/
N80JEwHQ6qk2jLCzKB2Fp/I9fDsCRLdLhodTNJjedfeFtLm2UzboXBXuQG9JK4dYcJw8Y4GJQy2M
H7/uZAxbhHDJpOnol6s0srshOIz4Hq8NEDhBJ6ZFqpOitWWmnPByZNGCgbHV89x9+sVjqlP/wJKu
MdZMZOfjqJ/uoPf8URocDbuFHtxYNAZT5oyKS0UXZMRPu7q6hDnwCKWKCyAmZMf92GTDL1NT6GH7
aqNdNwHyer65zOo7Rb2celF0sZ6I2vKXPfnzC1WDkefytt0Hq1814XHwj0sAXIw+82I8pPsVyrUf
MGd7HyvpWA3l28SKWTdbIHJiFcAZCmRyonp4URfLGbX0ATQUe7zHMXmkF7vhJ1+7Fff0zePqtHj8
f2cfVd443VOow8At42EYbTtmnsxi2PNV9RzCu9JewIKawc7YZ5T4wq4v2aYWuIrEAWnKr1Iqc22Q
EaW9T0zLFX2fEorxdi35hhijPrVuNj7v/yvsQ6fkBgGZFs5fZrNKDHv5EJ4OAcJOp6dkXOKcn989
poM9zvPam+cbZS47R06nAPbasXWjv1KU7baWiLfwWiQLieRuGX6ievMpHpfcRNqVaTTKnF8BwGd5
cBWbHLCgc1OnNK8d/f2LyfJuOrRYQhcky00hPrRASgdgNZ0lLAoLU0fynF/zlJVL6SvrnDmyPsPD
RCBRW9eSzKwRLeYEz7qKFcNz1x4KnZgtpKlNRJuSh91A58cwE9q3f2P9JHgLhRUPgSIUats797nL
7fu3AOSjiy2pxSyyd2DMO7Q1SYH0rFKE2qN25d/h5/6JBsOZHnQ7gvX9g6z52Vb2/QFR/sMSE0dd
kPqtupvDGtWL9OOnBfxLvthJzxauzRMJCsHgPmKoE9JyNG0w9Hq+bvJ+j6CyHluOhZ3B2oEJmLxX
krbTuCJUOpk6+zqKW5oC71lP4khcSxVLAYUahvuB5C0+MyJMqfomvCcj0uhUlQjZlgwWWoQOkiNh
rsuAn6zzxOXQ35HVcSaUraIhD5NlkH1a2Af3aXycbYtAMxQPVcOiY+YebIKPi8qzgeNQn7fEpIU0
EkXg0yJ4LsaBG3QdcCdW1zA6uqnwOWnZu7zEUUAQOQ9gH/IYOwz29R4QtT648cAOx6LX++aApPWg
gJ6rPL3Q8/XP1KI+iAzphIwjN0A9z/C+7FL36NGzapeN/MaYxz61h+1PT60Ls3FjWIHK8mqB9NNh
P2hx7lIC+PfqeEirfsNgmVS0ky8cgaarYDxfK1VVniF85XqhVIXgWZfBI6bYRfmNyeIH6ufD/IJ1
APHg2oRCwNP2jrHsNgErcVvrEm+JZgIChHTvSgDzGPWGVk792RH0fhJT6obRLFZOE2gk4RtpOJHZ
LVeyaAn7aLHJpZqRr0sOqRy8qZPkgFXdmCXAcwBJl9KEFYI9ltQ3gtZqtAMjRBjqrvk8l7X+LaSI
91KLpuosa8YW403G2uyoHhFcz3JPtoObqGTvDWpngPS59c0i6V7NTwsyBQXVe4EP4DyrM4Sg9iwD
XSGeVMA6WlWK/sPtKEnXIa5aL+NwOx+QJhg2X/ghOJNlwEexAi/LGdUHkLzPf97v1eYjqq6agIhN
bIi+ojcBSAvVnWropC8NYO/cfsge4dcXrnRUitUhEExRzZXytd25ddxDWLGggAMiY3+0o0d2X5IS
GpBp3xVny4yBRjX3IUyCpr+HUPM/QfW92dki4eyJEo+5hWt9bOPEvIaETV4UhU0XjnKjgv/fZ1Ui
x5BiTyOQHvEfAybzrhiF1ETmR0a39bINAGL96+qnnt3NbW0gHzIqMdrmjNWP+llTXaQx0405gjWh
Yy0/yezp+Mnf2WicELmwUumo6orbmUmCG+ipwZxKW5IwhUEOHddc3dCURGvXt4xNjHT6e4wVmVzV
eteOXUe0Y8hV74ZxtHrIB5TtWwQh2R818m1V/dlIBHgNh08P5+HOAcXR7lJnHuKRfkJHgdeoWxP6
1zlt6LlU6O5ql0ynaxdHmEMjf7EsS49cC+omIpFxX/CPQaWbeLIJqbTr/xkPMTUV9rDvhKDHROcr
YP74RSU1fjxN+MJ4LKRUxEjxei4v19Ov9S3BYaugOQ3Bn9rGMlp5rzer5TIBb8RWs178CVJ80/Gk
jd9h14NzP7UbWnNmGDti9ZR/ma+i+B/GlcCFahXdRGPihORoNxnKkAC4Atn2GOcVGg2kbOwuV2S0
GpxKbd0Be8eTCpy/mjGu95gaROKhRuzRI5WNnDeLfjHwmGoZNvjVieWr6yAPCqNSR9kPN0ZO8sUS
t7MbZwkd+IMmYnJp5g9uG6M4Kat2uTgSu3+O8TJXbFVydTlb7iFeMLxdHB7Uy0//dKBidLhTtJVf
jR+CxeAzCytAL/d0Pzddo0BOYG+5xjk0nzzZMa4HQwODCjnzwZIrpVpwhASj5xRK1Z7m2+3Cath7
BayZ2F7naWsgxt6FQNmn0rj4iBsFUoIAVmhkvEmOi61UtDphAVZRlMeCoA3+kzcEK1rdVujIMuXh
SQzujgyEWN8WgkMPCvrUh76juugl9xB17o1VJoRtkeJi6SmQFZ0O9YOMGwM03T2vs17+8pFo6uvZ
WUGdakZtvW5en2UX8Eb3OPBizJWK7eeMKn9DGHIRHrZ9G/2qg2ZAB5DBnUIJbWupjDCj1qXOv4m6
m4m/kt/I9AsT33rBFrr4VwQdQGfNzAUN70Xb5fLkaQI+FGke8Qnnu001lQzZ3AJ/IXaAK3HUi9ya
Fwz7RDcxabXw+Oe0+rP1wAlbym2nPDWo3LxhlQG9C3/YLJFhv4MlbvITrhgFTgTC3LRehq0Bo9bN
CDeDiW8AZqCKTeI2l5hoELfN5ZzSpVTsuYOstVpJY3U6Vr+kOxe2+WiitQEnjNk3YuFeqrAHidHA
8rra87Q/yahsMfJ2Uxyab/ua6GXo8q2Vviyd/CtAybWpiga5Ah+7nKBn0fq7OLCs124k0k0anGnT
8rj/nqQMXZaTjWqxZBy2SzhmIV/qb1l5yrSTtz5wnRfKwmky302ArVs7+GWZYZQ2tJ0IVJLIO/09
lkLkrr3+Xck7Qv4P8RKwPgqcq7Jd1MJxc4wtzR1i7dt+wLMUoa6OzOhZ312CQknK9Bn9SGLpCLKi
dDdVq8V6+mzeBjWShxXYu72JrJo0b3BBFaI0UzcqObgIaO9iq7H4KvYUOOaWnfFbvwOxAAcCTBcH
fQa2T/c5BxxB6swlHYAhFrWxgeFBWfwItkBY9h8F6V+ssF5PL4CYfjbCT5/Thrw/w50elxUn/YEg
IsfyxbWEo2oAsTSP4gzFGoW7o6zfGfN2LsBgrvyQcJOc8vdizosk95Qt4i+nbBeANOAtPeL41lcm
QiGrraUbslgtpjRK6XBmL3y187fRE3jLP7+CQKEjaYIQkQym+AyZZGG/Bce9ryBIHP1CY1oIg8mo
16FlSJfh8g8Fi/1OGzTicoeDdM4JaEFDvzHu4/pnqDB7BihN0DlFVU8qfLHDuq+v/t91VIp8oyTH
dp+goOUO6rR5d8GnOcmaNZP0FK6n8JdjhDvFXxBubkNZNn6oB3EFlC+hTW7aXsvO0w0Vp7h92dWL
SKbSbM6e3zmytPnNrhDcL2BtJUoG59+VVe+j3x6Wg4RghB5xA0/s1TUvlq4SVG4EQHPSco3aBM6g
Fl5LllXT3MNks2Q0KoUhC8ik1MQYO4MAbTIyivmsYI/8EZPRAfVK2KLGcn6Jfpb4k8WcIm24Lf/y
nCAS3mlKJaV1oOI2qdGtxop58ZimQRjymROQn2QS9ENQ24E9D4IYTbw03tdm52TH8DwrfK+j1osY
bZyqGts+PUXaUWLs6pc3OEOG2+DtwAr6T4sVNRExI6/RQD8bGi0GrX7hJCbg4DbtRGxaqT/AVPsM
AYzPK+sbRauP++SWwzCWoSsx3yftm/UV2josbo7FcFJ0tUtoXjkklDvvkwLnGQ2Fi91wGZcjj8p0
OFL2mvYrXNGe2NOKoskXXC88+QeDhU0JtHen2eAd4642QC5Oj364re+QtioszNA1Oc/0rRmIkSBe
jFv7FHIlgX2PnG9gpDJHMbbvwsJp/MDgYE2Gh7lIKDe00Rf3o5l95Hg7cZeQafWR4tzvNU534LrN
Zwmt9o51AbrFQJuHgzknUWdithgh/HkdjHDLhBtvBI7blaT6W5wNaP324Lg2Hz08RGrhGzwFx7yp
tflrMT0DODrr859v6VsvFuoQSTPX5uDN9WOybZmMKHn/1J/B1lHY5lZxoCEKiXYE9UeYV1fLlLkU
ftPwaNL6XOy/Wkxotip+Jq6JAIwMN9m4do/v0gMMm5hkTOixKTnmYBNYPmnVwDH3HgU3JFp7wh/X
4MXRwCZitVjefT1p8FsnbVSxZjhxMQE1vgrBz8hVw7UxOEnJrktTBTzQfUPg9Nv/a0NqMUQM5v94
mO6p0vkmq6gyaZiPSCYckgHptXqivncTfc3X4W5FMMNBpRXVCe/curGUOndDftXU5TnnhVlp6TQ2
5obMLhyEZ1dRVlCELx/MMDnES0NcDu8//ibtctsc8r053lWtYpmnbaAwXyTaiWp4vFo8D0UAPjjh
AGVAW4JHrTLbw5mlrgdxf6LraTJLoZ2HoKDKUITJ7ZExfd1dkp+Ia1N/dTLr/F00pngw62NdeXcZ
TqtvAL71u/rnuDX4UgQq7z0B/dN3GuyzjfAQsko3GrGAYtBgEc2iMu63splCev19jOxXnyTjRymm
//33dKaQg69bTBxO1Ee0fRRs4dCJJDkO4Y2Bx3nmaajYF3PZt30xDJ4EsvJarlrtNWZuZxEuBMYk
mFWB1z82Ru+BF0qUTwBs3gHUT0rJv7yUsQpAywLFQrXEM0pOkfOcWzAim7frValqauADJ4zsh/gw
x1r3JKTtv96P7TFKADEA2kCdzv4PyZExjxhl8xyfG1I0QVsQ6uJk3nk89z/xSOpWFyjXr0icDMe4
bHEl+r3gPLMQyblWrwvMg4JVCFsR5B/9/lP5mHbtWxG5P7JU/12pwdwyczlMn1o3y+vTUxzP1yaN
LgWuwC1jkCFAi551FNC/JcbxUuJASP2fOk1ryb9G1HuKwKtTDXl+2MUnVQ3Zd7ziHwAs4r+p4UYp
rZbhG3zn/xO91dQo9JqcFQ5iG0OMQ4hDpXGUycYPQbeLQQa6+/x6Fe/QP2XY/F+hAqNQ7xl8mQMA
kzFo/qyfspxwQr6xHP4aBFoL3yfIbF2tLj0d0/sYakAX1hnOQYPOgoZ9cZfQAmu7Npbu4fMlgOCp
jvfvsOXn/KxR9/kzTBjswqTG0Tk5GYQ1ndRFoCb4BvqLxFvYayD2as7Ce/XsiKDTiNuiIpipWrYj
cmfsm7kUmFPD+9bKSZ8EYBD3idubz9sd6/7E37y3a7VIhAgMOxql9YffzeKzTCPw7NVGUGbIDylc
y02oKW4Fa9mApXRioa20x71XY92x+Sc7zeIzbBK00UgUWdCtigclH699LrrrlRUHxVwvcMEwB0Yr
JK/zl0SobCN8n/fwAgdC2dga2SaPH6IsTCByiwNSnAm2iKxtweGMWz15ZE9sDa8bw5TjMnSqyQs8
jnZUd1c7Yj2gzQaqSPwiL36pVMNEWMoz/aPEohY9c8z1b3qHrLbbkv66Qe76ODDk029bzJvyTBSo
ryBIkwzecw57zhF23wULZyI3vXAcqbMkmWwSNxxFDhASNg4GpHsEV++ulFdIKneoMW9RTaJjD+td
n+Ehph8eeR1FQPlzgEwOg6YW7gRJVJJP7Aw2uxUJNE23YtCGh5KF6seq2odU8CBY/0YBW4DiU5a7
Ga7K1FSY1Q6CGabDrcKk33MfK6UfZh/6no4U4htzpJOaY3VRCaB3Jy4NxCslMjtIXdLQwHJl4EWo
h4/KgvlZWVfwj4rJRanGdd1MbpjUZeSmp17n6dsQr4aptQMKkKgKgW9PsTM8b+KwhmUGZE29VqcD
09LIgIkpAaBaGFE85+5IAvqA7KEzha0V9yXcucbw4ZH3aM8rFe8cLB2eM8CEEYA3BSVyn/nxo6Ip
QdLYwP7fdUuyQjxt7VlL0dOq2bqna4G9jlOjWA7SF7HPEkxYdEIF4nKu4KA1MRc5jFx9tJKTjj2B
kHelKkYMd/5cdUcrnQIifVXLOEYAk0IsJAIZEtwq4RM4jNFPJRwzMsAcdiGZk6Q+ehO97eDwejMg
Ss0TWbz8Usz1/M6IFuCv0ntYB/aexK9B4m33wg9EntLWwFi7N5g687aBaAbwW0PI2LvbGju0hBrl
ISnv5JX5Sm526SWnVMbxuxRgNZz2U6WNSkQSOh96wgayHsrcYlqyzgmA4DmKd0vspTEYxbKF/64u
kevK2g56GpZzVW1hlLsmgcKZ1Lx31NG91DMs1CDSViteSHG+9P/ulVWG7XY6MFpd1NpgjjiBAOjV
kmdtvvAMU85AOcXN/Ytjgq39e6oR+onCqnfVCqvotk65UyeiKZYhYqWe9CTJLkS3T85E5C4cFc/F
Pga4vrvj8ccDpza6PlLY4yRPnBRqKKBat6w7xkkO4thGhIPs1DNHxTp9Q84OQlnpm/7AAWBQM/nP
Maoql/NsHJwvCm8//xpBSqV/3uCRLkgS1mGyTHn97oJufuU8ICjZ+rdoNHRcg6DCS21+VhfqPYCL
BEkceRMprhWHmNOkcJpJEE/lIK3i2AUKGkFBKyPFkdJILzZNX3OXUIvVNJCxAuOfw+EhfVa744uA
FqYYYhvtLlZXoLbUxNU20it3AVTuU3ipDvzFq11s88DEDFtvip6T1CePQ4jUOdQPuAus2giolYya
+N1zducF3osTRHDi9BZCe5dFLlAX9aY8W2Qhl8wr/TPoeYw7kYVUFnB+tnAg+cj6VSEo2e9f4u5g
CFxl4gtj1IFN0c5Si5mW0NFjpsJRBSl+4f56kfVt5z0WjpEDD4cl2yERWcGX0QWfjL+X9H4XSjTU
qIlGgrptrTSBkgQa79AgOtRqXpF4msJuRQ5ZBj1suxwffa8rm3uWjgN8WuVMU/CZUTkrQRJtsKxK
c4IG5rMXC1wnpehdQlWDMfKMfpAdDkGqOkhG1hWgx7vUtjcPwA4Cyjzn0GWd6oyMmHEqvSTbN9Rl
Tj18dSdbgwFtW9lmiZdM0/fv1iUfB6FZusxrnnB5/R3nVpn29asKJXbZ3FFepO8ovmc/AnffOXhF
KzqYmFscOOpQt/ZazyCgdIBf9JnaC0uN8TtWS5TU68JVrda7tUv4iOACHeQul8fYtO09kR88Oc9l
vw/w4oPzvcNRp5zFCoY4R9JAIPawSP6d8D420XxNBkU+JM8QiwIdtc0vcvwp6jDJ62C+FbYDEcKi
XGipaEIWCoE0fC5LHotanVZ7dI9hmz51HH+Mcl0XHPlQEt2KwftnIKf2fZwZQpUdF5DX2MHVOGtY
f9e7xv06Jz8uxFCeZZlRcLvOn+sg1jwKZnBVbgesEIgh5l9g8NXXr0cQ12ejVhU1YQPCxMEiijwn
IUc+8/YH64eKP4NOIq3mhlWMRkCC8E0F8G86qKqyVRS3ygHnX1aI+Z/nm0FIgV3nHgSTb4xxemp7
u3NK5oLF38vj3ykrCdridaTNfstSI6FIfM9u4SJ1gHvW0suFrNvmeT6F/ZM1cp8SSVSOFLrQGyfD
WQtIWmbhUm6IR77d5pHPUAmO4e4XLN5hvW/eDpG9m/aXdzUWNxAmr6yuYPzNaVdrGUiI3cHsW1OR
zmJMxts0sk+tyDtz9gAOVY9enZ0TJ8LEW+WQyAHjZ3Hmi88yDGVqb5GNrqJRiLaA2mcSKe58QMLq
KkGOyTpiZIz6TcvUc2ukkbJJPygnnVxgxGbXKSOYNoeKMCF7sh6oGvnUVr7btTmTWmLjsHnwOQX1
Lb32vBzifvbxcV0TApo4blSN/7PzU8JHiei6z+/2Byf3oil4ybhPoPd+Ns3dpkKF6WjOBXB0T/5b
Y8bCc9wvU0olrq5F5B0IYqXyEVOPSGsbrE+qE7V0+ByLmBMAIJGcAAeEvFZF5fTG+gP0WMFb1goJ
A+xMJTOXiBVW5j8/fP/061t9Vd6WwnMRkDoB2Ubnc7hrP+gYX1MiYpkLn4mcrqj/ozfq59Is0vWY
PRCz6vNiDwaYTd8XxS1bwId4zFWPELeqtmlvYdO9/lOvUHJyQP5kQhjoBh/zQuzYLX6WT6TK+Xou
1NYR74hBpSY7okP6aiLrtin3kLBVYkj1ApwHiLuC8I0U0OwjRFSxwglxK9fi2Cw18W0AQKCULDg4
xSA11dwWzx+lxUNMb77xcoIx3t2c19zyPpBr8eMcWXNSUipGGjOv9q3mvk6ibBoJVKM6JQqIyVlj
6jnqlXzd7QphvCZ9A85Rb68WxrgUt7ZD+DMWGxuHnOgXL74dVkDPKa9ZNYJpfC0ym+xBDGK7FJBb
GjR/nAQ+0bxmuZj0gKtT2xhwt3AtBepI0Pd+o11GAhhPZUujOvsU3okccGb7cmCx85RtqeWIM0ya
ipZK2VF25ESC2iDlg6V+jl7cJClQ6A1/iRmYqFkHnlLzlJSkaoZYIn5lwEGiZkxz0nabjXK8c8Pw
sa3XxRUvYhq9saMZB/w8qvrcPtp/daZu0EucmL2UiOoJbmFQmKnrcBKMiHUmZaxob+YZnlgAJHLD
Ho6hO47Kphk24ZS+JvzB41qYlTgtvgjPLwMD73cGBCDB7cXNH55u4Kjoqjp9aCwj7oud103Y5ULo
IannHtVcpuJtzW5dXwnUlMVTTOfov1Y6OGAczp1irLNKMwmAYfryzJk7goyidbu3JQMh+bm9tQLc
Sn5GOYgU7PtC4FQ2PmQ5jQldkIeOHq4PMLrIkcrM13fQjDpJIXD2tPR8AOfkWdF1LuvdOOPyCI4k
4ELl1Uyo8dFAPU+TNx9RVzDFfau1A5KAqEUM3wLFe9p/Kwyr+1aY5pzRcYskED+3au8u6vDkT9CT
7RSfZ21NNoIKB/yRckFSWjiopnNzarQyR75/YaGyqJMlYHQJAfQAUEmnvbl7jmLbC4hWMK2F8P/x
F7qxAfE/QU7IX8DL/vVLJ7W+WPMOeUU2VfjwFG5z+/oTYQ+D/WXFD5ZnSmniuvA7qHFaRyGGG12s
Z2skCRao3JOgGUVLmZtNAM2KXHC7rH0blC2gnUYWImBEuNrgEX8FdJ7MdiTg1t5ZNCT30JB+m7Ne
0pjPWe74MIuIycKoRu0MDNv9TKO52HFYQBSk5LrNMtdQh6+ojREte4Wme82Ry+kwM6R6KDBuwt1U
l5ehaEMST4rbS4gKEKKSmi2NcDFrEj/GJ29YRfVYrDOU+DcJNBeiScz8RR1S5N5XhoerI/dcuI/S
8djtVVF40qH9DCrMqM6SdJG5soLhIsuEbrZ/cW4pqGhUgz9Gh/TlxBPUb2DrDraklDRjc6o9pdRT
hKOXurT5FarCt+9rCXQhm/gBF4t0yM03uHNu5dwGhtgGA0Lznw/7SyQfDAQ2TWL4PgJ1Rj1nDbBB
aiStxJQFbHTbg1BDcGsiWUKx7aSuhbaxWERKxTDY2Tb5IfFa2U0qXrapjM3d7wsFrfg7kTRp0xVb
Kt4iVDKvP3D/6b90zhSXsGfvTSXEJ0OqgAxdcrahCJuDtPGvPD8e9BeNkhm8Lo8/jekhtkmKhPbf
nVfiCb2pJcm2Kgepsj0NBIuFkRcTMy0Jsw0EFvWuTv7I95bMltIDH/Hr14T0F1Gs+NVr3v3eHLDZ
W870YaJVC/4GNI2o3Fj7M46Yh+6LlVYcX4teOO8O0mJnqmujAAvkyydVrMff/fIjC5lzcgF31ynH
LbOfA2Fp/y+jHXycQntFgfeY4AE+Bz4UgkNvEst4xPHKfYh4vgtmP+GABLGtisQUkiAif90FpL92
bnJ3wZfYypslSuZWJpmWMznt6siakP8Nr4GDSl4S9EediU0SsuWLD50LzEvlr73TG5iNpqavRkZ0
7BUOyEWfYpybaS5UVrX4ZeKx1WzKm1TWZfLNDAtwH9lidlQ3O4Py/BGe+LEP8Wjr5buWHtUkxFnN
aCwmwBzIh0Xu67Vmx4S8H4j4+9RZXiSg+U+eiSDTcPSTtb1cYxzkJTLtZ2mMecSYT7IZn8akOgr+
v7u+PJIa8YLFsBi4U/UIkqjxDzIVhKaiEpKyKJ6AuQkINlLzH4FzYPYYvLtycatuVypLJAirLgl3
ww6its5T4WRxLoZsIIw6tMgpdMCEHgDbGvvf/BGhJoVqSSbqye9Thfjci0v4cfV4DIU/bd8Bjw1p
jYne0s72gWoP6TrqE81gb33Jz9hKNl8uh4TZys+iKri2ZlV0JjOhYNt2EabYT8uBI94zeIBhZNHq
K58iaLUH37hbvc/0KgmN1ajjfaWleb652zW5Uxjg2Kc8IEjZawRkaIfPOAXL+aW+cn4Vj+gYGwg6
38gnX3rHnc5aZ8Zl0ETDh5X35AqQETyXFxn2TIoh/7kO9cyOufT/WhPgm6TI7j9MuAcGHclPUxTi
gJwhsCHTgjy4AX7UAdu2nqPbUQb29lE5cCQbka8m31T4pFxfuXMh3hcwCcnpzGWmQUXRPkTuwAyU
6a/WkukNRZZfv7k5eQTMO7+JNtevFkim/UmY73EO/FHOnJwBTZHHENYD3m0GVF+qJOyOyA+Lsd3+
UOmYOcieZcuVzG6RRnnW2AMl8IbhXzXIHC6DxxHOUr1pNnEIKURrS3HEE7Ph+gK7FHuIRS7vsOqg
HYqEZEIExkCf79FXkyCoAm6bLEgRf7gr/6Q+fx83xcAov8KlmECNqYVma8xW0WmcdsYg47nEGeUQ
JJruaKg2TJyQiDn/YA6JwJH+Bnqf3AMUeX2htCs4GYYjmI0G/sCIBvR1XQmLJXdNYzpbEQ96MdLP
25PLvkmSwviqj4FGYB/CHLgwh/wfbclKHYh1ZnWtL2UjqwoiK3/IOIbyfrrII6N9wkONCcWRvn55
66S5PKd+Od/hEdDa6ZDzdq7M+kGV3hWzUaQZqnF4DXJ7dN0W5ymhYBCh9T1cxdumXSWQH7fKchSZ
ZegNKi+BWE1OoNolpCBrt+RiPWbF2HsPJ0A7Jbq4zTbwXIaxd5nlB+xTgGFd/g18u3Iq0NP0KNMV
6yzntrPItMvQ3NcRH/u0+w7JfU0DMsOb/ScXQi94/wWouEoSEH59kje5qEQ7B3vdvmiqQ1tTw8qs
Qt7YLhvWYMLihyiXGwCvAZ1BVFi06cfKSmtrcEnKK0lhqN7L0wpJlzJgxGk/mUkMAtYgF05S66Oi
SwZyFqjf8LiPNitDU8QoqCjCG7WOmrSzdcGa9+zSUwi1dU+QyCxsKhT7bXj1NpWTkwjEOkQwyp2B
eoMXOR851EvGv/s2evdQ8ddljvieHMCGphTtbA+hBCHrjX2EMvz7xGNM409spwCHs56sptrLH7Ao
8ZK6LCecNaXenECydtyRnCNHn0+Iewio06qCuYC6rDqoSe4N+J/Uz3DxQUk41oYug32cwxR2kn/A
rkpcBujxQzRRTcho0REvJeyWlbMY35Zi2RiNjS5n/VgDO5Mj5iESIpaU0S+ghIg0X1y4cI1XtRv7
8GQnoLmWxGICzYHxNbYtPppWdpwaHQGLz5xLGMERFgRp39iaDgzHpoNzeNFu48TjM86fMidHPSGl
hjnxELCq1WmX5ydCtIQUF5aIz1sygtoioCmRweEw56fBX0taE1XSl9JIlcoKPVPXc2HUv7hyUBqY
DUT5UKzWL7dhOMAF8sXHtnU7S5VkPF8ql6lnWGg7T2uLkp/6qmxJY3xbU+wSdZ1tPRezyS40vBzQ
e9i6FZugCtPjtmzzY/PTImRCrkPYP32mchQEqc0bXfVP8HOtsGAGwaksfnJxGNXvSU9RHiaYXFO+
pApBcgwcnF3sUiMTIheUEFxF1wCRNGN6KT+rP2iVxB8dNuk6ejBiPsaaGNEyQtEA27Dghv7J5PfR
CvnjKEdFcrc75QWUoHqViXtlY3xvdAExiqgIWGb2FeuAHDCLYGXJoNc5WjySP8IbNdEI1Hz5Mgis
sLVt8yDzAN2Ygj/3um+WQWsFOuDXDqPK0Kp3SR7k+R9derm0WLVFLGka9k7LIBPJLrVC+WWrqE2j
2K4MKxNc58Lsbp6nGEvBxBqR1fTw+V7/wY70DfR4UHDmJPIAQB4+bxAQqvt9YnbjT/N2DQzLFj4Q
sDU6Jh34xOUXc9Fln2ijgqlVMZ9FJBJPvqtdlQ7MNWbh5njDMatTOvuTeofS8UAnNB40jDVIEV41
NQ1uv3mc7dPE01raoucvib/5nGzQYFcAAG7FsC2TGIjGtwOYm6jT8NJwBe2Wd/qP5KQo8Dc0z8tz
ZAQanXwh+5f+J6nU0FUEj3h+vaNJ4bVotbzzMA+dt0uygPOYJq87bsjWclqJYfSC7Q1hNUEProp6
EAZprnXqhvM4vEEiDE238KfsalgDgIpau2gPxuFcCpG4KEY+bfkdjRkpRG2okqT7qf93ZLFeycRu
EIGzyg1BuVPdInueg0AOJMpy8WwHBXQGjgvmiM+XrpFb0qoF3ncDJS2tVyNdWuu0o5hiZkoyzmJ+
Z0f2FE1OXzKRdJ6ISmKzKhQNjLt8u/GqJi4bP5AQKnE1zPC7HoHzA7VWmyJ0DCKulK69LbgduHM1
sqO9QlGM4LVw+4JxgXKL+Gjnf+pdRaz0Opdi8YIcb38Ieli1ytvZCjikDhY5sb3ajnBQlh8eXv74
3r5rl0cBz6xvF5yN5W34L0lfUOUDDX70XdvwG3Iq/PnRH0jZ/IeXFUBCASaSLPAba0ZS68oxH29f
RMdcDRUpb+qxHkOQ+aBAOTg+ykYAhb+k7iikUEpTtplG+QPNnD1PyAFSvmXQFMAQNhcoUYkR+oQH
mafVjm7ZZTOgmKXExq027X4adypCWTD/ybViZMUo7MXwos0BI9Ra+fyMcAJt+VLns37aMULvYk5l
E1mUq+8jGch7bSZ3TIIEUXG/6BRJ750k0GpZEOZG5vlWPQc3yzUCYdo4uYspS+CEYA/hIwinGqKy
fpVwLhuiEYfcycof1bsnGgMFqM7jbT9SLnSBQj+8KPPruJqfaglR3+m+BNyNuI49B3oxeBz5QBft
3hWxYtOff/MUwSG1JjcL2o7b5DywK8yhMsbtWKHG3TBO4z2UtdiFG4VSU5e9B5b46ASncW6Gb4fA
YLwrCcNH12idZByxX0BP5I6cbD2EiWg2DLRlEjZCJKkToBCxieclnO7hJRmpYskFMDy0rJmsTpKW
fIvMe7TResVLsTqQUdxQwwzUV4VfLoOzq46bTuJHvaImsW1kxDjbKv0lvgFs/0wlkryKhi3RO4KW
mOTAc5N2vYhXqju3RAr1EjSZIAv+4Ycnr5YLxam9rC3EOaB5sTHji7jK72bhH3/5cUInQNOm5bPu
rsS+scPx5ebDSHiDFfIUBWm5hzCbIzVyWtf8aMkJ5ZtMGYXkBhH0sTjZ0pnZ2Xjit3i6O6GIZgq4
oLHA7HAGO8zUPnXY6VRFpWBvOsslsRtSjt622r9u5jqMWlFX7OFLvnWJGhXrERkcP6u1Sipo1R3y
nLlMedR6PtbgnDw0MxJzELCGICm9xSzTDIDevyagDecHHNMXWvBIyaph4xQgwZm87NK3EDfDVljO
JdBMipNz1tHReNBO9trVZ4TYF1Db2J4pCSq0JhW2sSxNHozSHGywYGoj9uq2vgT02hTYPDucggg4
WwoOT0T0ZNgjoLFiHKHjkFw/N+96tDNPCLZY+U7vIVkLD1MaCkipF6VpHdRxf1FmUllq5cJuCZH4
5lw+LQIchh0P06f33cT1BkYR2JyHUlrIUxjhPKbvXN3yFHLdvbLZ0G9JTfFX96pufG9a44sv2bsH
yez9jmmlmJct1N+q3/R9OZpqa+UMtFJswH2Qpa8CK+szXeL3WzgW6ybpR1+Bun4/dYtOTCu4IfWF
6LpDpm+qcIXkn65SL/Sis58kl5aT8aBCctsbFzUEZ23xpoTSpyyRUzoTTGaKZbnVgFmFdzuldBND
zjCSMeo4ASIfA4dRKbKYsyuTk8FRzmPw6XbuRyHLbDaqFV6V+eZveJNR62L7jgu//WRaLMie9IAI
zLN2LPzSXhJoyswJpb77AGfw1Dn3q9swHjbSzqzUObI5p03/pqa9jJ9MRTjuw6A3TsLAt08crg97
lMXe2MyMCtIaAky/rqWabR0k13QdDErTKxMVDjZNkMnBCjeQ/asfOizIM1iprie5PfulwhJnvLZB
X/YJm3uXL8WJZ3TeF3mFejROzbkuTNGUOfgLfDeT91cTFkNXBLPdlBWkOFgoPjMtH1TPRseUCBsB
BoO0n7hQmsnKWTXxgzbj15FOzcgSOwVn6o+4x6FWc/EtaoJyQ68R1ngjGwXt4j4M6LaaIZ0K39Wi
uJKUTyVbtfAavJVZ9EeMIUIFPe9Foujmv/WhvX2cbDuRTcWS5kiXOz81VIN6pIWjK1e+1YwhmFhV
oWchp0gGEMhWEC2EqgrBuziWI9Z03bqIJFmWz4OAfcQmlWsbE+WdybHkuX7a8m1KzgTxfiK9LjWH
6GRG1h2/n598nC65UKQJ/JEa0VoXwSCecZTy5DL1w/FgrCYP9nOV5J+ZJGI+U14XmFncICGTxi+M
rP/FbndHlh4IUstRoUd6BnyBGuOy940z/tRXfWHv+PxIWa9mP96MJgFQ08QqRmfaffHI+d5/zlwU
dGDhCzrrNUeNZJQ8K/Qbn1HNTy1e7cckgp4WbJwjL+ApB0vndO7QpAyLtVWDaGbwuG+85ZY38an8
Hj06njTjWW2pA9mGQdsqyPLg/sasQUEH71u+GhG40Y1l/MrZBUaGLP0XZ/dDSG1pe8u4H8HqupxB
SEq7XGQlgGbb3RzvIbMgaTFRT14rsDjpn7smu7zR3/DTWyEJmCEZDNVAWtmvSkA7HEq8eoK1nsXk
iEfGB8tk9IbQJnVE7zIScoRVpzs48t7DQkxlGLbH0offUKTVy587OaoNm6XhC10UeT4ZETptuQ13
/b1FTSwNRiZFgl2fTsol6t795EN2O4vdami4ehyhp2oHaBmWywLzo9sTDpq4i55A2Z0TOjiaMPlx
9zPy14CTQQ6c71MrTPHV5TN4yag6Mf6/lGYJVVdB6JiImNWHoP+Puv74OXY4Xsnr3BecNWwD8LH0
jZW+TGqn0Bqm8danMfKCPHsBSSeqLY1EkEd9xVEpnjwpMQNqDcVujPqfvYjAmpDT/e7I9LFG2Z/c
HAM/OlttRMv+zpnGDzOeLqf2W0V/UMxUxicE8SqMxcpm5onSJrzDRxCfQ7h5+SUII5ACE+hLxwbZ
72NAzJyGuam3y451shkSwYoI/5sYRqEFlC2yBQm4feZSDoqBIU40BJV9qXTpIC01dP4yyz6J1ffy
BOESKJLH7YQwP1f3xzOaTccLPm4cwUmIOMjktsMDISoi/9lx1XNQrhCeSY218GqbW2PCGAueQ950
VsYaFJuAdGZJJtUfunquYaW3ZXD+LiphlgeFVZ7nZFdBMRqGVy37zSJMjCa0J/6JFJp8KZD8yu8V
PrJakKsmEuN8HJWUGlblanzBbkIQq0YdMkL/m9ifWzHYAE0a6bVjXZUQQgVrKJ31c59BaJFK8v9s
0Z2CKNMowqVl0npVuXGuL4gaUVHkk9KTj+2VIC2s+8/KVYcQ3fMu9DYMQzuEK8vWGtUkPJSmG3+z
ZzZBm6cZ2KB6lQu88SQ6WqQBYDdT/69M/AvpE5CApb5ev7MJ9l6VOscO2JX2gRWR7SsKP+GgIM9H
xOa88+I4I1EKA0Kai2/1T5Ylwv5drZ6gtjAZZS4Ul2MKM3pCk96QEyPuCPwMRgWNmzACXPOjUBbw
70/hGd11kDKeOpOkYWgfCy3QA/pSRWeqEXWTlzIMiU9Uq6xjPquHfRodlTnwTKzFA0NzB34OBYi9
aG9TwSmGwdFvNqg5emTQPLaUq/VXfDouRqF8PY2BPQo6eogKMeErET0kGrDgzUYhZFFygqRmO+kv
fj/o4kTeQWkViDgoJE2Rbgxhh6wVrhyqXcw1tXyf7mE1b7KqXQ1r1LJzAAdsRoMhXylp7wewHF0Q
HfRfGeQPt6wfpN82smdeJEztCCjN8lnThWUFv7ojOerr9oEwxd2bNr0+Xanvc8NEeia1tkisguH/
L6qb75OyO3P8WxO7XXQnl07Hx/CX+bwQCFki4byGTApMZ9lSqmIBYifImIoLtL1Zj4LBSlu8jk/i
QYnAYt7AKAcQZTTtkaeeI/JH9mHTU4VgJxOYDgdZEtIb7tRgJMRY0MQM4JFubNkpNc6mK16uH+4S
AoOXkYWsL/7sWqPN8kSLUD0rW1tyo/J5BrGb57waKkxZ1tjCwVg/wB+0xih4vJk6cfnco0pWeLZd
UaOFU2lPyGx+0fkoZlH36D8+s4w5T/Zsx8XGOezz13MEhGDtmx53BMi1m8/Bk5vNWjG9tbEII6dQ
2/4TgJPcxNeRIK/PnI8l19ahID42fuffLic9JfNXXsKKxzEY9gr5GBye5MiDcta4RfU2jP4ArqhP
RIOMyzty/d1q2TccTGpz17uiCqHFjSSPHrjTfeFFp7vzB1ItttebprGAxICrGdZzlRfyU4jTlfn2
vaPKKarlGOImsneH4ZislgQazWGg76+YAWqKbLATjjvV6GfoJX7YdS+IQ+oHdZBZUIIMh4dHWcz3
UrsKcQChJbKURnpo8DsDmDeOkJ6UGcxwrF3i2c1xOTK4Dza4o1YgNy3ffVWYAWJ6uSlCNCpty9Md
cjXRSjdCe6tPjkHkBk8Wj3UJhq9LABr31P//I8LK9qS6Z8GQDpO+2Xl5Mc3Kpk/eehY864yASSkj
cvE+BuceukzSt7BmqZIUhHdwtbXf7Q4j1z3OsONoXgAJ1RQKfUySwF8H3toUe6eKXKo9Iv7msTpn
Ty2cqD6ZguOGEZgQRAyy0M+AzT06gwnZD3hvS+Kx8Lv52IyByTToBOK9RtBFUxuhh29eDbQbEz1Y
xJ/wJTUM/HncY8qNcwQn54YV1/ygY1zFo7lddnxtAGfwcBQVSJWvdT+jA6g9N/6hdJbKsQ2yk1BL
cuEa0ocWl6MiiN0rZCjq0+XDSesz0UGwQoB+85jn66pNBnfWKfc8YfVEAUHAkdDXiAP7hh0WcXf0
VU1gHdGi5jiAvjVlj+CAd0+m49r8Y4bkhpE2/pNv2BQjgyGJlWBRK9eZ2rjvB5tlESBgPlFRz5Mp
t/uSk5zvOvIxXL39eh7SqkHPnVbQC72XCsGV6JigbFmHZewab+jo+HoAb1c0iSzXIZJm9EFxrBne
roYWE9eO6avInVtJvmvN9V3sE7RAzOC1JyiHKOBIwuoP5fi2UxlUO78baq8sJ53+8/OIlozNhP0d
h+ag2TRvPldGsJR4spq1P//Lz0Pnu9Wg3+ifUG0jaCUfX83OO2iOPrtbI19zSthPCqUSROSVeGMO
1hRNJuIr9WVmsYw5seOIH/b+QJYZmZG8pmP0sYRTYI2UHBzB1w22J3zgAPsmPg3uDZQQNA9vo1nx
JUAWG4YLOTOzYx6Y3AuYGXrAakjVOJ3D1cudGrcLkCXPLmhaqiMRU6Zu5CmLeSv7c4C3B6dpk2sy
5gOwChBxd83bNMAwLhPa4VVFXVDQ2zxRgrDwwXsTTAIBDIOuUkN1MAW5kQhnJQTfQAlLVU2612gu
ytX7hICdHa1rNV5Ixdd357uBd/3u9wDydqgsF7OqCZrOy1nuczaywZG2JC4hnYtgSDwDU7yozt7G
BKhzObw/29hXz8auJPkVLqv12Lf1Nv9mJxOR0yPsj1TntEWk2UlBRtbVWCw8vq/MypZPVVaQCqqb
xjbJtCUG9c6zJb57JQXTPXiPApSA1Ygaxu6xPS0XvWdJvQ4yGYXH/ox5xOL3N+gbfd9+WigAp1o6
oLhRBbOZLRpOoZM190LcG+/GvLASMHbnb8f7sv9x/MRtZdc/+b7NAE14k5/mZVXexIUcJTSSJE1t
yEUQeaseYCt4T/wuVYwUWgQMNDKOet6XuZev7YJ1dWkAiokKrQO/qXCuAEc3CTPzmQGfHARpP3Nd
jTJZPgChmMvGnWQI2SNKbPRRg66eox85xLz+736RCQZcsT6Ju+MfC/8IZ2nF+g7hFtROc1vmJ8oL
K79N5hqwI55Wa5goTIaciii8OAj9iVNP8dNv/K8Ioi0HbcZ+tyjSukJIHsiRDyAL78BBIH7qB447
XTPyTYrqeNFT7/1GMuJ3C9dfHrSCAAl9wYu+Azb6A+pPozugWRVyn0Wsr7aLE/X3RQv1ElziWRSn
OFl3Y0Wvhthsw+8tiEyh/MGteGhYXVtgZLOgrfpmNfBehynb6/7AqEpmxS20pJYJrmKiR2Jyq2gH
X1+MBkYNcQre0xBSje7rM1cVddPkttoUjzyZtN96/NLdulfXwKpOudn1Ix13YeYRfbJ76xV4roap
nJVyPIGeW/ArRsYJCLUOvfEh9DuHnbzXQrpPpQsb3ukvezCYJY6hL8+iwlaMhqg6+PxYQF3Wd8Bm
ue01orIhV9FSdAlbQWDGacaeOEK1mvYc1TSMLnz2bTe94f1kKmImQGCshGPa0se8mwv9nY/6huIv
/+ln40XWtbcKBHq8hdar1cebLhN5UV2h8EI/Syoq1AqIwNNm7CjIbRtjK4iNYBj+NExbAQ7bSZEC
6YUFUTHAJBQGsC2quNpGTnttZGt0g4KnGMTaJBvT0gXPs6ZZxBzRoCFSo9HKFXVIKXee7rUcLEkv
f3H8zSnuN+xENqSbE2/SfTAil5ptCPfWn2F5sctJ1onTZohhgoGMEAQHr1qf/ozRZCOd3SSVpCS5
BStwP7kWhzt1OTww/x/K8JdG7bGwZ4zYpkPTSTYoPkhDrchjJPZSvm2Vlf/HS6CiY3l9oCSl6eek
LELIP7gNeeETebIOC+y8YB67HKmS0HqVQmnU5mAZUh6Pk2OecC96uxhb9jKhXPWC707mTDspWBof
FEUxh/7le6pF8aisoNvvsyP9LX8skxyLGKwsMGH1ZwA0nqsHlbQlMFJN5D3Hfyw27HgbcD4/H81O
3g9RNZ16posbbWmnDqPHnK6ciZ6bsTXiwSqAlE0dPrmllG7oTOu7H+7dSMpYYtUesjq/0B9dIcfQ
Aai2rYalu84yfLm3RSAdHt6livB/cK8vQY5MS7j8Apxn/ygbkiFNYBeUte8zCtAzXD9Scx4nwQvg
zdIdkLYRGXQzgwkHSXPwV3VAZNyRhg+0T9Iai7yQO6fVqimVYcRjJjwTWgggvdDR92o1ef7EFCeH
LSXg2wn9C62v5R5/l5hIqJ0El/oI1DJ4SfpN3hJa9H+Lo4auihUWBmRxhQxSSfSu89vI7vjdI3qB
he2O5sNaM3URyRbQ+jjw5PzwFmlt9Wds8JIzctpohsHGvttYipUa8kI8i+hkaZpmz14Yl9fVM0Jh
sAqvvKUL8T7hRkkB2N2ZjPW5732VnRvVWgLzbGFHHqjdjiSLXri32M2LDobpxndHiPmrqRD7RwvJ
I4PdqOFnYty5+EeqmOSRsCOMCg7KOvxCFdwD16YJeiBXynquE4q1jXL5YDgso+KltNdtihXcaVx+
axpCMa6cEWhU01jU+2QRJVbCrhNquEIIVKbU9bNg6R4HDQoE5VFADw+Nd4DSFbC8nls/WmgKnRLJ
CXKkzXcWTG5YyVkiJizfTZsJS14FUgSKl0FxI5B4SjhTgkoMJ4yHjYEn9fLUG/ggBYg5AbTgwyCK
1ebibRVgX5/AujnXLojpAvr2oCGWXfEoEDyGg/UfhKxGyFc+tUmzhTpGefcghX4TTWCYkBW71PLW
ri244QNBjnPABBZDP3pAc91dn3lDzVH9qbg+gIkJO82JKYxLZ6WIGYZ8tIR3ppHx012wEYV5uZvx
/TJLJPRo0KYzBGv23/UEgekMLH9p6aTE52ohUO+S7lU+dmwRpBvaLl4NKaoQMRHsPXAoHC8zD4F5
bmGIXaoJG6yPhf80a5d2CIUiHP4dglMSkxxtknylcMC3VuI062DsHulY/7AWicdTe5Nfiqq4QM8Y
525ji5lD+mf27bil+hzuwavKIJ6IIiPjj/vdoxOpT6T6zYxhCKo5A8XeQFx/wPtl/ZtORyd2A+zH
6LGRMCyoDouYEVsf5gyG0iqr6JRul0zXvcC9sR3o4/Dpx0by9LXdjeeRq6E+46Sno5LlsrvZRf0q
Ob28hmHjKWfhuE23tnoTykPcpVQnhYVicq6GYJErA6zbxVA0RpnD+aWguz9EAyziFeqCWyW9vENU
CkMa39de31qsk6r9h1CIhDL6j7zooq+XYEhbyWx5zz1hCiYSovGcBfVXRYQWsJuKy61F0kZS7+Df
G/T6Wau1HAuIqGzXcWcHZafp4AcRlaCzpBCGt/nDJYhiHsYusycwMcp6Bt9Sw6OQ++HxHgt1iBiB
6fkdpNL4IRvbXqZJQSpJPYa1Enwc5z9LEwcjAQhsgz4I15C4MsGIj6bshoaZ6hXbMbovQfAuPPZq
95f3dsu2skL95bQOKROO1WSQPEZEfG369QJhEhAusXPUNtdPH5vTS5/4qimfAfwTgxNb+ga+bUnb
x5oszo/53nmwjFkUgAFx+HjBnv5+AvLiTve1iZBw+Lq3C+B5a07yBmu1jTuQ14iovXDNlG2BVMO8
rS0HgO28u9fIrFm9HlwUtUCU8C5BZGEQhzTz+fOe91fpPpJDteMdHUj0UqJtskJRPl2oW/Sz8xBB
Ks30LRE2Jl6trnUnZBPcmp0tIX0iFjDOUFCkEUQQ81UpGqet/H1NQibvunPgamd0LMtW9O7UalyF
GRh5jcpgopPYIlYMkyxId3rjbLDq2Ph2D9Ua4QBI6RJiTGsZBcXptSboXFdO30OlnrtPKie0QHUN
3juLtBztu2lP5ZJHPmOZ7mTqpaPyrvj/FtDJoRUgoIjd/oQ90B+wviYSvTm7doyh98x+/T6DdKg7
Wq6158vhYRgaobomgu7TK9LKNTogPBSqyuO7n63YExnJrmP2YrUyPTLZvBPDVpdDRf2PNj/tuEfS
qLYqz07d8KOKXMSfzynr4AZrpglXHJUm12QU630rlHeoTdSXRFyNGAMadyh6l1t3lZkmD9O8iOz5
hyEthV8MCMv1DJ1sBCvIcsscNKiVuO5cf+YYzGNF2NSM/S+0+nfkjNpCWF7oVmbe/o0zVG+PxYGZ
5X7m8xILwYBOTpdKpRsTYIWh4gmPlMjjts935zri9SKXcrPEhdc1cX59a+qDQLpfn95uxPWPgz1r
g1tTTI5rKmNDpURreh7iHDB65h2Nvi0JxpUYGJ4efCro6T4OD+wbUCCGgEu5z4t7YBQtj2JgK/ho
HZOhZE3i6IzKJ4b0l7AqQSI+TKMmvG6Psp670rceUDeTedUhjTrhRrf7kJSIb048XqGmZjzrklZ8
/gDt/dzsjRHQYkLy4RVAMLVY/oGfgbXZRhzHWVl8jDkAsDdZnhgPRLWtrXGJBm5K70MR+T6xwxz1
ZpPnu84BsQRFe+7Cn3fuGNNzhu7hygwkFpBSg8fsOFIjaMjR0sMyyHVxsMfJj2kyS5Ur+mls4jgV
6b9QfRZAsxXXXeynGeINtNdlJhSMgTKvGjWEmLgUurNjM1qLGjvmKRlQygBIn6f3/fztA2aq49ti
bL2w/OGBNLIS5sZKfdj8DhaDrsdv8/6AGCvJ0ZpJCEQxdTrwFW4oNHQ37mrdc66ufYNrEMm2l1U5
R10FOb61ofjvu9iXCnkmynMCzVKWpTRBC2//TSBWDPo+U3QPJK75O7CpfcYCZ2nk55Xow2KK78IR
HS8FA2NxOAv15W6ITFj3XmKLU45Y1hbQDoYP3yiOGPPU9dMNn9XCiczS82KxENdaMzOx2z/+J0kE
pQig6hiw1wu/u4RtOBiWK4ksbqnQ+kYIcdD+BP6bSr7j9sr/1gFZ6oxlzu6lX5/1Q/zhKvjPmR7y
y/xGLmpkan7GVoi7MS/cVlQhKl9D/daRDoToMwpwCF3Bkw+SgmaIlIogNvS59fiFujunz0u+n70i
cexOC7X0GcxRRi5yEAAmfmgPGO7uvgZ5qyrvXzkfQwoqh2ZFNjsodpsV+AN2hV6yNOfW7o8StW/U
21OKWLHa8i/j9dvMBrxTMUAH2tvNXo/ykQgUqKTijTsVHhK46Hu+Y1euQk86WT8AQIdJRXp5aQZA
wFWwGkFLGvuT5mSJnTQMQCSiJRQVOeHV0OwMrGULlE/XLYfl+Mk43J1kxOBDmaD4ldYvugww6I7V
Y4CdIqnf81lhtcPpRbcNxElAJC6WNjosp3rphZ75l+eYa+JF74y9CANclleYZXcH7p5bBgno4Hvu
q7fUOmZ7o3DqjH1czbk3CCkmjjetV4pzkAh3CxYKEAbMYLmDMI2Ih0guxdWwVk887cqB00WQqTtZ
xDeRUxJ1OybCmI0jIaVc6fbkbry5S2vOdFwlTjKUa3Snu+KCwD2DSyzr0w0gf3BhyUHnrBuoOTBK
5/gMmgf9EcjWkt646WWsToPQobTGefOOQqeb/KuNwyoMUrngnNqBXwT2NsZVSmrQFWFdjVzjaF0x
fYZ/mHAQ9+sIamn7a5vzqGQWaMkZKFINxGRaCwBG/fHxiDReVJapc/mFEue/S3mn82nPN/f/Tsgh
xS99cpRka7vzn8VbR9Fnr+UP5EvEXs9Gh6/0oa95nxZ5+JRgvEgRHmNUlfNu//2En+m438oE/w+E
l5KVIbbQhrXfcN8bxYT8kaoAaRp+xbZ5alSwi/udfHPbwkZVbShQehCAUff0wBfdQNj5sICvGuUj
aqPDXiPu0vB54Ew7y2ugm+QYmQme+BCyMy8+eLEn90zKkEWc0u+N/aZM5gk4eH2wCwKDuHD9fkqv
/Opq3HZpvOW38xuedepHuYi4HagoZ6YMDE9JToBHx1kwexSj+tXmUvHC9JhzcSAjGo5/pBN9lJwO
VJDhc5VwpCWRUtJ7r52RGGon8RIyyHN4yhcgbq8NuHFOnPBg37rPz4m0kVeYKPaQnW2E0yKXLFeb
L+We4yrddICz+e1FCx82UiCSpzyM2+g4KdjwdO4cljs/QPNeONx3d5/Iz5pP1jCsfzrQd0ZGXPZM
LfaTB+hVTNYSI5fgKswkPbwMbw9TQ8MUvO4UEz8fVjzpEvfSHahZLsNpAuHla98rF45Vrm3jikeD
PW60mfduLytRYO5NIlbHgPTBpAZS5hgjhMsR8C9Uselfl6tBOxM9gMg5yNZXwUMMen1wMPYCfoWo
Usq0yJykwGTrD5ndGXnlR8s4U+5oDQ4uXrVrWwSHqZrrob3pgDlZeq1CB+EGcf4pxNe0Redf0UyH
XwoIM8qktoESgoHGK04cF7SyZ0C1aEh6HRipzV3HcubRmiHQzjAMqcf89b7p2lVz2QIP/FcSMU6K
uf4VvMM29L5z1ra4XlKMSP3t/A9fUCRU3wZ/6KCIbBo1jptcapZlFGmycfu9H7+pvjAQ7jclT8ch
6z3iPZadrcwHss0pZHJ6FfNzVSFtelQA//qmFW6g/Bp4//xA5CNlkfdhFvi3Eg1Fl5cmsOHOO9uT
jH2sHhLsY4kDTNjDB8rmnyJry++BpZm2fpk6Rt39kRv66wAD2UtY+9pQai5V0rlgpRebs5RsUzh/
xWokAiukfx1FFcSjjBVJYexNKOXFtm6glhr/zol/mCUpAg7Sj4OOtgygZQbLL5mq+EC57S3nxX0P
gyXKrBILu15qdpyheY/R3pKRndSddKXGlryf8jME+p3OJxOSyLGCDbIjBEMptdxK8TpBSqQBCxcC
BOYoCHUU8NKLhqZPY5X1xGWyq6qrZSUQOsP3K6BDDbacIBdAYLCrgy57LDnYkzOr1wu4rdVBaij+
RV1QCau0ip0iaurfoO+JXo0+1MHzRGU1bfrqJjHTpJUd+b47XG0QMBDe2r85yYtU24OoyUgStTtc
OxPfZAtqetBAdxwtxIDum7jn4+Nb4ybLJIzhKUirLttTWYTdddOggAtZf0Fg/OLVTgR+25JPSw2T
ASyDyuxNKzUhCm8slzs2tV5Ftxtf5wTZDAKSwjWC+FYJ2PTFKzR2bpb7WmttIGEJHlzViidLxsQx
8jdUbAswmpVSi1WPxnpW76WDnVzCGmeupMbjZRPUrIXLCBd8XxwMKPUdYOwceoR7hFpy2SGV0OYZ
PBrpZ7aE0kt7YPG/UvoqHOE4e65CsRkZhlpmPvlTBmgTJZQKdKwrZ5Hm2q5p6S8dbU9muvb2QA7k
UJjIQw5nuF/IeKDi8MihKnx0OefZNdavPqkZGAsXTBHS4uI3e+HE7hyXohWnbPrFvR9GmHjJbY/5
1Lv/1MZxfbGAXHA7ddneHInTz7MAHFQCfDP59AFa9WRGsswsfRBllb9Axtl1VG4LQhN3xxfNsn/r
pznRnkq2hUAJlvx08Hg/8tt0IJnmnSVnoH5mQcoT+y0EaLQDxo8kVPqOJqE+KmfpP/MSpe4tiIHF
n634BJmT8hOsg7/yVbwI+J7NGeuslQ/c4UfXXUcoIF9Lcw53qNOD5QUIttaFqMRSaT97O4kDtpIO
3Q3I6T4VY7fk5VIumza+zU9Y3Zp4l3GNap8IymSfAeg9mcdNt/gksRo+sae3A+cssCPZc+zwZwUE
ouAI4rUkYjH6lCbpLMMoL+OTZn9KCJXedw6DebjY0HO7Rn23+mtBRLAwUHhBr7C42O6Yi9hczfIQ
eDXivvBzR0HtSSUQQ0lU92ynFDCOhdX7apEV52gWSzU18XHE8a6sJ/vDqcE5dNlivSy1EkW5Ezdy
ecoX28cU+yBLSlZFNNP+DzENe0Ubsqsyp8Bei2tgdthnBQRkjR/nJdh+oqw6AJlCaIyfoO4ky3F6
0Ew/6BmJNUQuyURHz4QC0wEX4IUnSwpBgvW82jKkJRZSAFlFlgWOPHWDDS86IW2IJTGPaHqU6Xbx
kPp7SgDCI4r6VmXA2kYt284GElO/HPS9NEd0iELCiatNbvke62xcwPYw/KXBb0WWteVQ4Qusx5qC
eil9l1sYgsYP1ecCPyB9IobexrEvUJIhpt4EGL01Y3DHh/qLYuLaSZm6Tw1FH5Og2WxSQsrkC+zM
RtYdPRzsUzbO7Oc1fgKsDFQXmBcHc4XjYOMtWUHcsS9HZOG+sUBc6F4Ua5I1XQbIys2JQoTgCUaj
auDIm1nl0fZy+6z/ZiGDZKQuiDINrS9XeXBMP/qtvwLCbKMLhAbXf1jtQ4Mmfs57WgjkcVC1dRxk
WT+mNYlSp+4D+IMcHyBCcRgwkORXJChBq2GTGUoijA04esPNaWLBohuh335BKkljzDdkZMYzYdhK
Xm+tLwv8kEWj/jgIFMxa+43t1M+2FzDkjk4cX7KqHyhZNUHUWWwEJ38UPHmS7t1+DVIPvdOdWEXb
boI0M+XMa4b9cLQpVC8oo2To/mn5KpI9jH8aPTALSyz9JNkW7lxROsfGWjYWbNZnzKBU4E/GMMQa
clCeDQFwH6CkHpn8VO5pKbJUadk/3EuYLIetkYKqq+h8EHjx52l7hcRD+g+Slp8n2x2NXfSA2TwX
7BNsJrK5EMBRzQfi2pikhK5wZKps1al7QTAKGATp7xbEYPE3PFvX+sEiP2qiDlYcr9MC7DYP1B60
O8ZZwruI+ghtgADBCaALOsYijjN2COAuX6aSQEsmCmLSREM3El41AZzp4x1YNQVY8Q2rXX8If79+
/5ySR2pBa6qo5wT2SKLO/TjKJZDSW9oGjrfy9hOaHdBlEuvufcbcpV72jCVu/k2rO5bcc8xtYZ2K
cTnq4t+g4paTUchXQs10peoGEKGJ8iwOKAerwS1wUas89lQaanK4eYiI0h4cfIuqjt+5YcV2QTi5
BTgMI3Go7dbTX0GYpoc+utWJ7HHI6TZ9MmisMYRwHDH11Hvax74SccYUd25e0o7UAFUCFG5a7/pn
vP2Mz72WBeUWFS1UiWfJLt4kRKxqzSJWg1jTPzqIVqUU5zGIZrYGUCDFNATSPO8OhPoDFiVrj3Qa
GX+UgmUinSDA0OJbFw0sN3IZiNjcWfzA1PTBCDsBDiURr1/Gu/z8vkEfJl++l0wM3ztzg31eL/s3
q3yq+Ixt55xJLOXVks+4U6gZCEc2tObLZIX/da7Favm/5v6W6o6G4eLlWvHQdajeHb6oGeHvkxQe
zLOLbcOSQA0SEPc+MwdLOLzbFc+nk/rOVCTf+ilbJ8iCHTkQIsenCFBsx+pL7YXcBEKi8N9sKObx
mdmcKJvpZmFJOa3YFzQGGDoUGK+DYw6H5sN9jeE/kOfnHGbeReoBAKj7LV6Ux2Rj6GznGuZDW+7L
5Ci8xdFtepuxkncf9NvUlbf/yQ1gwYWkUu41RSSAzrE1PuAarsk2uKvjXYL6INfYmpI2IWFscPUT
YUzg9ZVIr1V6pWvuK12K0uo1Vj7DCarFIyrcp69lQULKB4TTfKUiDdta+IQoLuDMSh2t8cc9Lvc3
6HfOQF3bN0ijhbvj1mKOIAXYqEmMVZSRKfKY9+qoHX0Bxsr2TswQC10ajNkXSDnww+mQiD9R2lDB
ny4WrsNFBaAgTttnV6XsOxh6VjbdvW5kJGUTcGBhfuQOfwvYpYObYUpSPBOPulC+rQfOL1NawZQn
BlcJLKYz8Rbl0Edkr7TqkcXVp+bLD0p25xDuAvTYaWd/+TMdrWFOD4jyIFvMKzd+/qWsptO8A2s7
lAlnWE2aG7jRhOvm/uGewJ3WV65nqrjguB1yiVzXDdh+v8dCKRbZ2VDmU+jbK/URenTxJgomo7rh
IB5ZYyoFWmJ+3tjh6UpmxTOEMiRGUe3Vh7pjeiYX812iHvumhHieHK6jBBLmW8FCLdPiCA9Zq/21
VKB2Ld32LQb6u68fAVsh8ASgbMHf3mYsrCE0iAg44MzKRXXO01Jjq5sba1QTtj2BKJAreER0f+9I
QczRWaJSvmiDTbwuMD8LxNv3j7gYScFcj51YS62ZxuuIs80N6AyBtLvxm5zUc/hUraOdKR5LANjP
Ff/rGYl8PXOo1uh3anQKSXEcpFvtMYkkFwvaKsPYzUZCd4o3w5d80jdSEqdRtx1bQ8opmza2dgFf
5YwCFTc9OwAZbeIBq9g65ZDRbAjkFZ8wm9D06bGSzoLNVaRD6ixbjBSfKZ4bJXFVpS0a4LZgFax7
lyYCIQo56th9AXgaUbjYOEGJamInajCLfFbE9oEz4zI3ihG2K4Tmw//Oph2uSrOP0ADH/BAYczTB
bKdvTCONqxzm6dkRuaCw8vnKjhxQU3BjmlulJQJoWYjmPW/43NzeBnqWf3G9StUzqdL6lzMdFVPY
C/s1XHJyjiqarNSkP0ZKH4Jg9xZmW6nMjHoPpG1tTabumOd7rk8VjF7oxTH7nULNQy35j+fVMfWB
MrFnJAwi6tAFqbYMMmxOy2N1bqSz8gWpVW5I72wOp5YIsgNhUwxNo+MdxS/DAo6vGgtQhkg4c4j7
VgZbgLAJyCGWu6hCTZ9eHe3kQRCEiNDmY7oBffykE8Z7Yoz0cD3jXq8U/xXkRk/CP1cMNqfWLfxJ
LqGcCqpt+rX+jE4/6ObUWsNvnqa8QQA6Y8pSFz+Pf1YojUPRXdoCYWTaffkSVNJY9bywWuN0Mxoq
H1g70/4e70D8dimIvXyuP5rxtMLmtxbGDhMLkcKfzwz48ujO0/Jzi8dH17nYEAFuFiowJa6UMJ57
RTYy1dTmH6Q8RLH+ogFqfq8k+KTGl+/AdW663oswCIpelsBBwVkDGH1wc8oZRfG7zF9mT1nQH9i/
x3ycozkbl47pQTZkVPjHwaQMIS/mYpyu9O/mKPdyPh/sLT+gB9C0WbjuTb0UOu+B1zSQUJCcZozI
AnpRkgsrTJ51DYKas+8uPit0QnZ48VBGwsH/PoYbIBJYSQwHn6Dja+RkFKaHzibAPH4/1sP/UGmO
X8t2dIvFsItySoOiY1OkR8a2uI27hjIpYxk4kp0/h+egPPHtq50s8sOLwUCYpJJJQAF3eNy6pNYb
JKPcBjE5Fgn7R2orUIV2Hgi/W+yBgebsVuuXBIpCXUqj2E0v5/ItVbCAW2zDYOJfHLHpzWINI5ZX
7DdMuh+9YDHIAv+Ac3p9BLOTKRkQ7IMA2VtwZ8900ItBUyKYBablz1/8PzlwTJ1MhaBZiPMPxubW
glxIvjkT1jltiJTeKocNhH4ZWNLF5k0KbdraAcq6sUkQ4FC5phkhn4C8vxsBOYIpiMTAx+F4ZT0G
0SyUXvZgZrTGCFFSXTse0diERmU4TIRbtul3U3euliBLt5MwXnRUtH5mgdKGlB+5Kozg/jeAzSgk
FNe8C7ZTk7DdToWhvxxiUlL9qr8EPvfeeG4CfMv6l1ZQE33XduPDmw/zRVrqHblADOAvvyQhHvmf
lsoaQWZkZHI+Gns+6h4y4ihMsAF2JMJVfe3xmEDY2gEgy/fFmHz3ZDco3z0T0Z6gaJL9w1s12qAM
ecsD38irSz03gRHZYokuSOMlY7XH1k/aglUp9hTgzHSiTHDjNBJvcyYPUA8Si/Rb7/6HQnwbpAsu
ruCij5ffD4rUxiP49vce3x6CkeOwoP9z7wIPDj0KUDMKxVdyQcgzahDgwGwIMFgnM8OSvRFv/8/2
VSJoXbVBk5Ip2D6oYzSaic0/bsXr46ePOU3jQemXotNbK8zqcxi4jWeTmbjjJFdidZIKMEPlrJpn
qHELWjRyyUkMfp2UbRCs2IT+JnymbiBDVL9Mn63+8dedhmMCRtH6S980R4GLE9sE76OVNYD0vOe4
otNnk3mHbGnY7r1Q+s48ur63v4Ww9k9bp5v9ABdjlDwb7UAvzp5pgS1/JaKeDJNyGhoGHA/ghMp+
n/SBBcAAiYv2YwvdjOEJ1HtgJoSD0LisHniY6bgihAhAPhZDW3IjPQ2UUTIgl+G2h+hOJINcrptd
cRPjOetC4q1GSmzdnySnQGtwIcchcm/1Kxs9PylHUZOhA1pOwdqD6K04dO8ZCzLztNzmlCCp2SYM
e7wx2d3RvKlnqZTYVFGjnJojk2SbvTI5o1uGdVfSw1JENO2evnQ+JSUlMPsZCDtfxiiKUfJgg11D
8wRCwqmfiBCpOwoDS/osfs/ddPHFncNklQ+XVxwEBCXaWkoA2Yxug1MfoEMurR2IOS2RqxlRuHiE
pxgcUCabEynpRKkSPZc/aTqs1DicwGUrdJSQC3GXPefM82Zh11z2hDPy8sKXxyd36yuiiQUEaR4k
NBirBKG7uXtEJIZwvZL5yCwIxv9Q/XqNkCsSmV2RU7M4m6X0McKuxwv4S8wrXdHurL6hdeXsBvoS
HN+GRViKt+W44/2RMvLF71YOk5PKjk01NPxDLxqgUBllVOkTsTZ0OfJpY1Q/shueax3MQawUsu0y
JkS7DYnFa3hQJV9Ikt3hswR/yN1J9Ihfi7drKqHfexNIyzwk8/5oZPpi0z+ixHJGvKkRn74sA3D2
4SYhZFLWnnT2AMeCvjyJGjxj2j0lI/4TBTN9q1SAqGzydck7ZJiZyiE9Li3srRKScLxSJDU0fB8I
Z/PuzsZ4YT7JmaApL9JQFkbIWjX/Lahc54D2xkOFkKjGsVUVr4rkVHv9COaOwkx8y2Lwk8DZ+3bZ
dYc8bCNqMPlWYjQ2M/q1jfurHEGt+WLudJ50b7iGXYuPi3MRhang09ncOOhbuQxSewOueQOGVwr+
jTvtSB0BplKRGTXX9cFUgpH2fZW99zOYzLlFqtX/wmQaaE1TphZ7FNFBMxuxcckEY9Aa9xIhiqF8
lfCsf+pY+C5hzxm8rmtgb7D2B7NtC3/TA5Nxf53TxEFFRzaq81+Rt85GFZEshQagxzEL9yJFA9jh
Wqn7QbI/b96BC/QMReApL1XHQ8hdFzy6DTKlrzgE0O5Vfcn2lqf21T16xyv7b17WkXKhRGCxk9u2
/QTnxaNHWK61XgYs+V6Vls8Fdi89SAqFv9D3nGEpcfRrWI289F6NV1wWv6tydRS0c3a1BHy5VzXQ
lBJZeZx59T65j7+B2Adn+Tv5KP2I17V768WLS937qKPH1RadnKLb9tN2UzHCYVcYe4H2hNkrFJZT
Q+sfLC8vDMRTd0ORWo6D5DhQv1vPJGuIIDkMge8KOsEeg1sBQWd+q9Nh+5ooOPZ4zIq/VlGEcx9y
eJzmgZVOhQ6Z/6HVSPTciGdGOeBRLfPtajCojf9RvAU1uPTYjR7bN4fGmRkf95rZPFa86Vl5KuMV
nJwDUEnRNySO4CLIhU79e7BTPbL50PztR/1NtuiJXM5f0b0LfDjEoDGTYOm82NyAiacEOm2kC3Is
jHhAD81wGcTvIoj091IttLsJcwH/ovNPQTHquuVcmGr2AjCl9Bo/j/sX82GNTCEL7iWxazK2XUiy
AoUESbTDi/bZfoJzX4y5ZJXgBbFNpoyKBF7ZSaxHxWQYeqSBMAT+X31hd/5YqjWQPp0GW97AL/GF
QSYexauzjElJ8/rmI9eaIg3N3XWi7O3iyQhzVlIytkM7bakT/XYBnlzlYDpWL6K4/LyWI3Rb/gjy
GsKJ79X4xOYZQwp3uyuNMZ5sN8P35tGz1WGLGQBmIhdS6fzRplayro5POhrT6dBt3nDCf93go8ew
JqmGLTQVEqbs9gd0BiE+HKTCweZJ32YPxGnT4YNm336dKCCkvGeB0R6Zo6bYD3Txc7UbchxO8yyG
F23FJPxmRCuZ4O8w5sjNbvW4uAfeG06tuEIby4d9P5FjXu16q4Vf3znixNaFzl8BkH0iSUe7Eikr
Sm2V5FH3zsm0LOwtEVd7iwX3NI4CTiyJrBV8BCDXC+boG2/XpCWvsWU0pj5aX+xEtUjRXEFRRbwg
OxtcZ4USI4OiNGSP2QW97yiT6FN2uSh3f9gEhpWBum2OjDlO9pYEmksGLsUfsnfhFf3b08HAaVh/
XYm94MB7LHcqpf3anct0k+oNhWbmmQr8bzsadI8H7lZiX/UaYC62d+/bDLUiM/jByNqIIJG/YlDn
NB3i4j1RdvAQr7Xra4ZMe5A4VRISVidPksQCIDGTg5DeFZEFd7Y++QucovKePPIDIX7ad2X/59dL
118FbogeZIs1fY+RzV0IbJQizX2c1oNcAAMhscHz91ZNDmdA8P+y4ED5ZInqTooFu2P9tFmhtq5x
2or7pSBGtanTK2Bey3YJMbX2CivgI86YBJTLQEa2ZbNQ8zdlkxZYIXZlsvS3pDQB6iJgluzBWMsb
4cwbnAM0hi+D4NU5gzsXH2nNbh///3apnN9dLzZzUHWo3pViFvJ7lFWlmdhaJj3PSm4OAvAx58qB
b11dyiKNsFOpOHq5DqzCpoRSjmI+9ZvpaM4t1m7AGDlMRkPV9/WfO7gRTYuQyyQIRpxgx5qdouqX
IC7LqE+MI1FpeBeXxRV+uxIlFvgdDvQiL6YdYWknz8sIA/EHUqiCcHu0ocJOblv0+AFnA1OjvD2s
oZnSS0ljqUwwVmpaiaYNjjzyoQDTiVN32bdWNtwY45pM7WUhFkc+p4767u6+tjMggmhOuHB8Gzx6
fgfhrIqgrVfXA5EwUMvedlRLdFY/ULUfiwYsUwCkLzsO68VMDsez4pmH3Z9FqwWc/Rxjq8ZQOKWA
yHf9wPAMNfurersQ6Mt0iNqkqaSYteMGq7hzv4hNC6x65/qzP1mrIR7N86ZKHtBvLS61U5dAUvZU
i+Oet8J0fUSNZUhmQOz51Z0RwxuWGH/PcGkD1GTF1AyQsEMvLD53hCkXnVoAT6OIltnfBYkLt/YK
lstkI35IL0jugA5nP66lKHM9+M53dYsxe/EmLsZxiaXnPhhliN+0SMgc/48QPkgntQhAorQVQe0l
lOXeXl5N5LdfAT5mxQZWLRQrO/ezPEzRDWATKWfOKetbFZRRTB0hxQztg7831PZF8BfVRqYXhsD0
9TGXlOF8Qn4qJTWXUSapSPtr8AxN0cQNCwanny0NiLWCvCs2K7QcTUjBPe69NhxbTpM+2aeVEUu2
/LxDZEoLybVGobMBM/7kJRn67BJp8RDQCtVV6vf8EvBqWsG33m0jpoAlzvtWiGqG2UHFiS9RO3Wx
rHIpLASq1taPLVQYAp/UaAkanekPEzBgQgj/gefhI43QzrHkmRu6GoLaIrO6nQLLvMShR4m3dCqe
Hbat+TIvdsOy9jFWBpGJCr2TuatQdsFnIlEtTj0XwlYpB3Z2VagrqMzTjTa/bhjjBmUA7C/z8qfL
Flf5YSLjIdNvN4pTXFAH+haGAKYiOOTlzS5WuJTNSUSxN3Kwb7+zyVth0gQk+28P7YWEASZMlwlc
nFsDqU5QovdSSMyaeenDBpi+8WPcycBOkPs7FRZEGXmyWzEbatA7FQVzkmOd+FjHQ2xM2iCqCpma
6YBFcpv63Eyk0ozpR1b9fW3Dw4mLFKz2m4FNani+/6zoNrRdKC8GfOsHjYQxHlk4tSursaJ0FNap
6UFCZWm3ik5h6HQDNlfFZO68Iewtj6d+S9dpG+amgbtevWe3TZ9sU6JfSLr7FEYp69yHBDe+75Lm
VqZCpSanWXzTMtcpo6Ddz0mwvF8oGbGtfAdsFfMeCmKOIN01JMidzamtw5n4TCTUwDhEszvxOGQU
qRYBFZ02Ew7jpkAVnKvi1Now2MSQazlTWSovqLjiROT8UkBPQrLxwOuBVFXJOHjiPDtyPTYnV7rK
uzHrf93wyMV+lG/95dZyc7paPXi5Uc5LwdcpBFQE8oqU59UxEvhy/xNnpbIrv5asU2EEcR5eTUEe
Kwh6itYeDaZ2l+tpemrsWtlymXJ61tlcVU4OwcSAq8URchJnV57J26q5/NY7tCyUj6iSOw/+qdi0
hH4KhSu+X/q1dGAD1EPQkZaw1m81bmcm9fBnaC8pWgHR9B8n2fqot+HzGqKoS+SWHRvAY2Nev/vo
WRzgj4ZB5tNO/lX90o+q6YuezI/i8P0PRB0/c4uBLn2BVCHfSuUVjCm+kq1mCcOpQmQhkxa5cNKH
QHVp8K9LwdH8N4lIl+Z+OjK646F0yci0S0kuaBZTSW7jO0zehFAymlrH88Cl4vtPVLV0M2syWNGL
qeSHx4LNp4+W0y2EgqhG5uuGJ7o0cVSmAU7svKDF10vb45DjFMQkcxJqO5bDJkhWR9QYcH7yn5eP
/p0rztQzPzB0Q+7KTIzEUgi8GdXfvl552DtuJZ77F2uCwiNDMvfolBl/d8+SE3nODCxhPvNXUqQT
i2XZ2+x1qymSFaRsNY1ngnRs5CNCYMC3OqdampsdAeX2726oVCFn4cL5byDx0GCLm6pU4sCd8GBo
YkKB7Fqow4ROpMjLSaROQgu/hlBQLbF49s8/M4LGEU4x7WOafVnygrLLKxHz8NHotqQQSu5EdzmW
56SOJtitHUw3sjNKOqH2p9iKtLtC/z4o1Sz4JFAHduE9LPjb19Si4jejNzyiCgQxUoZSOtWvh02R
iBws3M73y/cM4uE+WpVrqVyK74t6SLa0Qde4xnDcUouGYQkvtXEFe0H7kXhNB0K1M20ttd2jZ9Jb
1YY2ghSNF81lUJFcmP0c3NXmfFxYlV5+mPclRpRbXsFVBRAwjSRh7HCR3E2u6JeLE3l1wZrkdsMB
rrWxxCr1y24AZRhn5N4LfxRX1xQ+wPuNHmx5GHmXZF7LbUPYsMwh3IAjuK0ZHPMOIpdnIG2Q2PLC
yWwsKuVdYuHqn/JSknQg/YD97NLYANM9XeCoXZyLLgQoJe3pFqhd/Uc2OxkyzLqe/rJv5Itye4mx
R4DfVmFtFjgsIXIc51sOi+N3QESyrmleP/xpFiNZRKTgA8qlrYEUSrCqx5dccvZLBDDsqFdptqfQ
TUDJfYTjBWcHa36ZvU44gpagoqa7RUKiOQACc9jZh8URzUdEm+6nwmbjsRZQqABPY/ZZqx/hhjbk
UpWGhwQLmzzQRBX51HnAOfxal/h8M9FAi7OysIUOAL93xOqFbOPIK6BUpoYwiQfhMNvvTdGVGTLF
XblQB5oSf82PqHqw/GuTKVkSEs8iGmzjJGtxZtzqDYE+KX9Q6po95JIu0DR7Famu8QFfTkK38U90
FjuVG1ebvZ6MDmc7ZUSy3aWmO1oQDOvcBacWvw62wd7wBqth7Jrmb92ZOCkaCmiAyvGS6XLKObKk
2Ly8BysaOglraNKfV1EKJ0NU75jTLJTpwI1a+bgCm+Bshis3pCJMWa4FZ7FYtb56rGGRvpidhfAK
SoJRPZW8wqlvNPg3qhVgsp4364aLFnxy02zq3Np0nzEAfDvlZFhtXQ3cjQBNXS7sSzA8gyNwq+RS
OEHi3/NfK1D3CHft6R7183m7RtMe2UI0NwWsdIYCxPdhDIkGAaGtCGRXWRLwIzo2QNbKIVX7RpK6
AtVRmha2xczz6z3CqBxJ9LE4q4TeQgLl3dWwh6gsQo7L7qvxU5XnrGnJ+NeLXVyI07nyrsHU2CNk
XKg+k+O4lOsf/M47jgC//wjcQhcQ6YExpUmNpBYnJYqaiFSvzN3o6VT4JdHKI9Lz3Yd3PwQVSY8A
2RHowwWc0Amq9FCOY45nTgmguRmcj50hX8Mvq5DjPdV8LMGUsJmzibwShjr3yvZcdRQSLvK7v4LF
tl5uMJ/6f7NtihfXAO0/xoAS6fluaq9G6uGDU8nIPKarOyke+imUh/PRAvyxFjzFcb4AHDYorpVV
OH+cl6jyqlaS9dZ3rQyRhhA7bwaKsnV8wExuRe1tNLdFpxPt2MIIzE7iKGMOD3/NneB9HV83iYyX
ecH2h9FY9Kmh6d2OJZoKX0QY/Bv3o1MFLB66wnk9U3gsmc7YCFjnzQna4O+xrA6QUunaZFA/z4nZ
goictt3RbC+lXNblzoSTRZqlXJ0WFQpsNo7rmEsb9dCZukI2BKLyP5oBg48u7m4bF5CYGeI3ycmC
GBw9krYn7YWPDDJFMR/nzD3uOWxpCBbxLZpgty/bCZ9quuvWY7J+3SGoK5TZLv7nAGVqRG22wggb
eTAZUbTEBNihWanytagfpy3lPOEuhP+8oOd0FJMsLyCvWVzvO94pDH0pKk+Ip6bkuL49VzjOkMCI
MwR9DroG64MvGyXjVW2cMM8HMN6DhU+6L/DZtndQyP7bCeEFKUCVoQWSqwjeqICNdfJh/FiHMRU+
FPW7HMaN6FyC/Qp618+mNwE/X38e/MYXDWYgM6gSGtQqtUFHC3HudqYifS1nTnjcH7zmNIZIMp7Z
9AI0jvBqLIhHat7HLiWC45agrJOcuPPkmcE8c2eHjFDUOrRzj+IhPnYhpHJVGIcOG6E6CV5dOPGR
NWNDbCKweydRXNSk5pRm7p00zg1pfb3/07LQM7BF0I+1anWCC62hgxFCyKe49SpIqSKS2HGBsyGR
2OssP6lNawAE7RNn8YbR16e/9wevssZtNh7Yp0jPvpWHiPBj9IVH2lAzuf4irdZqGSi8yU20KYoP
RqPIb4tubDcMj1AS7+hFscQRSPrRxQ5Rwbin1chTG86I0BCiepi5qSy+LIP5PilpWprpL4RUsG+N
AmORLXeXqPcCAOgsTIvyWS3myQAWLSfDDpBaCsS3SYZujuaVpGOdJgyXzlCH2F87OsxavAQUjU2C
PMtmRhYDQXAQjVb2+FY/fX9wr6D+9yAiPkJKws9ZqPOzJL9EIRqAEQqec90t3AynMY2EatxyW0zF
eEnAbqJGHEDEeWuItGuJ+6ONYkfwo5UssTZL2oswiQSK3EFutrMPyRqltsfWRXYyHvpDJcBykxhw
JvtG51j5141LrF7+TO7Hgat0jv2WmaDEbt1iWRWmFpH6Zrb/dRA3CMIeARrWeMSk7lmmCxEdNMmO
PpAAPEK0vGs4BpIzpTnIB/+A38jD3XbJTWaA8Flf3RIpZt04gkX26AylWjYIU75ZC466iK6zWj/p
npEJUlBTDkXkf+dTygVNzt2ITdg+CRN/WF9c4fsHHqkZy8DOqeqNsHG3b3//sOHORtEU9l/M7W9U
qFm9BMSpkcK/8mfiFF3RdOQ7Y9PDQFPu371s6g6gxTK1Mvy5mf9pugUxEOes8zPdD7QbemTvD+uv
2Al0nF80uzhc4PSGjgUBDVC7A81z5EPXVHiPzLVbLIY89itgulFOWNpDxhfVbeB3IyHdgfyWBQTj
iUsQvcDgYwCZ1t+V4HjnT5Jc60ZSahOJ54g/xYEo6iGY8sG/wZlBWM8IsqBnM8dMR2nkuu8wesyk
AGWtisDKl2nvg0GCsdRjUboOVJRQECUfnO+lLMDrDTggfxJNxtgO8rPdceFLJvk/9nnqSmY2Z82R
JUjC9OAlsIbeof37zaSH11tq0zNHuevbnMgu6bZGIAQ57SwoJFVhyMFXpeo/44SWt62ySNg9Luzg
qPhP0ZjAy24EViR/lBrS4bGU08cJ9ic7P9w6brR+5k+vPTDcKh163dQ+nPkxnAtvjodfDeJD2MMA
T+uZJ0rYmmtLYmwsvMuYspulu9iw7L2O26aWOMv/Hb/+rvnRhUD+0iGOAJ8RvSreOJsN5RKhEIkO
wKuDnMHxLavra5uYY83/TYt6BGjf2+QOyHiDF4UG2fdmbCdf4tETm7rAVNDT/Ld4DjRD26wVu1Vp
ceSYckib7HjkzxWXJ30NCZLmEAq559/7guutjrNljHWJMAJKVKJPZ3w4drwl93qSd7IfDsTdQmfU
JfsPuF3DQazX9khBFynTYlGR8wZFfw2AWGuPylQ0tQUSNf1znFGmObcwU8M8Juoha6w2fmeQgDUI
KTHxGMQz4eLrvX80AcPxv070sdlEBfVk888OdZHvgkgYoNCojkHxa8NScESsragu7s1MyGsWcPnO
4epmSPcHW0W+IxHwuSptbMJaxB7sUZ4V69wVtntmR1mdMspZUlBl60cp4Kqdd1joMoyWabm4y4/4
vemJDKZ34cbS+3XHz3i51jPM4trUb1Jc84BxF4uhE2pY3iWaG0rz+kT5PHwNCGRKZfzIJX1/KVvO
d4BgAoMylK9n53JXRV1FbA2i9lWUIr4ffHbNESQd/FSXTIViSPmGEalj4Li+NtAK/XuigwRUP6Du
1en9NtN+v6pOQ6g8SL1ZRB0M7hxi23GFICHa2eRUY40dTzdJfAqnQpWu2f2j5IpK2u2k46RpMWSX
2zttAfCdRiqprVn9vv9MtgKf+HZzEuNJqrLq0Gkhfy5aXJv7r2HnKkFTNkCgBgm5wTRJ4p4NcgYj
N0aQ0dDZzmnsVjcpL1dU7M8z6xQKuBKSQQvjMeqGfk4hyRKaBOUcyXQN4iK78q/iuT3DKERCfV8r
ShUekQ+82rCIaQXuUZ/98UoXDNtVNgdH+m0IGzDoa8q0YvplME44DvlTEt4ZbT6q1qg2OD/J6hVQ
kFti5OzQCx3Lo8JaJvfcA+jK1s6ocWYt4+ymd7ypYQPlx3os2zc+u8sF+/l31EIbX5t8FDoJMwua
gnC0f0p2bSMjcRb3odPCaQRXuizrUb1vwhsRuYkPtCa8iEz0SfeOjjwK+KzNQQqQJtcTgQ4wLSyD
LOlvXVhxVR1xFv9+STGEx5yu+CTRZ4hK/6DiIxC5p1IxYXt/UXeJDGPlmDH2twnRN3m+sLZ9Fc3h
ZxO+iXxUM9cyZ2fKBmVU6NgqQbr0fNTPSq47GV/t1eDK5tQNBKXTXAEBGrqbV729aAl7AK2Zta+l
bprD6BO8SatqJQ3V8F7n5UBjZfusTqCjdwJeZRCFH81i/5zGst0/CmnzFNGfJNrfUe8Y//CxuJwB
BS1E4GDCtW1nZluyP7kY00tzQ7n57IgRTHfzp2JdSwuPCO7g9kvidXpru78rpA9iR6Zg0oF89Wmq
Z2+DolGIQb2b6ktQr8oV3zKg7FnT/j1cbzVPkGnbJKNq72UL0vNAghN3dlXi2sd9EU5Tmfbs5Xbf
CemxVEhDfxwpVtqWEyGD+3RLnPb4C7Ah1dYjSsr6iPdWAdniUhKVNTmZMKsoEAucANEpwbUzexWr
z+RfvkT2xN4Pm1nd1dwFwoMLOXsrRCTOrSWXy1ymmf85Lto+RGUAzROwmh5Wt+iITSfeVg+yIwwZ
Jyj6RpRtAf/8GXg+4PnDWcgFFuQ9tHcTyT29LPUWAvgZvFKXjNGVFK+ikrVWNVzEpqDmB0IuOGWj
rg9QtTV7JpODUx+8qvJLozVkYGPD8j+xebREeZnTB0vn3FZUh33FEr68RGNlNhj6+qhgKEmJDI6D
XpF+OKTWlzzdzAcUwMyVttzqNOK6PnPnEGL5rbZTZO4azg0KIlokUn/8oUjERbPJOfTF1J7rkYO8
by5b9oe8CslNxuLIvOBsDIVzFHmQkr4bhtvT+q/FrsOzFHrdGENcx19Pfi0pDzc9kn5WldKsy/uN
apMnheeXnU7dxbkvYtOl87U7WnMfL5jHMSbxBK2gPGknxwNEtd9sBFOGCvdwNyGt+lcIUkWDzSAL
2Xtd29kZRIT0w9G13t5VNEti7to/Bu4+e1xDHW00bGyGZ6anKFDo2wPrd9PmsyTgn5j9HAdZWEtI
drwTyEwaM12tGRK1TVoR2C0sRqhMsNRAxYBIx1yO9cwY2v7xOk2qY6fQ0BouWd7oEFYWiRPhnAXT
iSJY81akIq28ERicVlQtlOGEvacpDTtRvQKQfIXRDL4tQmtaRUMWAGc2oMyDRR2ZG4dtFqDQnAf6
SI9XoUAPDXpcHpjIa2WwDyTka5Q5nI6jK50TnEBX+IMvdHdlEqZisIGZ2FSfje1r1F2BZiB7GzE8
kX9LsaqR5z4Qp30KZL5xAGelSpDpasmNt6Txl1fkvIaH83PLqx31teda4e76vax9wx8Gl/dUaMS/
O0Uhr1q7mo09OjROVK3N5VpcR0CbfIwHX78idJLWqvNr0cL55bP0ZlWPjL4GXqSnlcg2EN94RvVs
nRxr/jUhMMU5Yo1srcVIXMPsMLKUYNTLYs6VWgpd6rQQHRpozmetwIhAWS6HTHCfXngRNSJDu2sM
tS7PqN6tR/vklWRw/6B6adI7+yUmZKrYlm4bVq4nbkWJbZLm7+Su6MvLestEKB4s6QzHXJUBDr4z
CBkVnWcbv4nkX+oCWY4HnmzVUzN5ynp9+2v5K7Igmor1W7YiKymef3svqDjcanuOSKbb/UIPKNZM
++BLiYYKXqH3PP8gbsZ15BCvQe+XFqZN9l+NvTYhxhbeOp2fm1zMxECSUl/Pme67WKr7nEtJPone
FKeTkk1EBRYaDCYN0SGlYEFkiKvLDSaUs4JEwXsvsS/4fABrZnXl45TYpin1GoN+RNvFUVdMmRW2
TyX2vvPKQ4IBeuULlXpnKebC5GVMAE3yxkSQtmJwDN7N2lVHcj7FmMtpOW70mk1j0Ivao3gkLkQX
pcGPwirm4utBKFibM6qeUBWSmce/JJb3KQLQSBBvYBJphRh478XpWW8GclslemlrpC6IPnwypnzV
I1vgLfZFkWLisKlXf/NosRdtnMelsrXtrd9U7Rs8q4bSw0r5sAInvRrPsWEmG7hyK8rxOcAmrJ3G
ofG+q3ajqV4QUYq9giTXlzTACwymTvZqVqPHeJO5fO664YqFHyyuv7BmTbkRc4gXd7xT/u60di5N
n1jBH2dSzSvLaLhw0CrIiqAF6H5l2wcbF5k1m4ga1nNKVMMT+bqUiMOBw+tvsey6EdGbLPKJoeE8
IyQ4VdKAwAsl4trqrGs91/0I/6Np4sITpdcyZ9w8B6vsdWpVy00sbAuLwv0RWXg/mgU+KCceHayB
KXrbi08TA9jgAR8bQHGKxVfGio1Zr4OH49ie/VRnemV/qfe9rvyb6Z8A1ttImWykPHYaFZ+iFU3U
MvUkPMPy5M7S3zZ0BxC558Z/Rr+jGdiTzrq5mJfc65yefHzm/FDsxJxY1XCiBAUCp6P/r7t+D7kX
6+7yzZbZ/i4igHCGl44TZKGmpW3YG+gpav1hZIFq6Ko++YdnRvFz4+N+zjcbeXtsL3cC+DmToLXs
YHNNV6GKS4BHgWjLMkDTT6GX7GAvIVRHs8QQVr5Xf2wDBowepKUDLRILVZ+dNSxrnUlmFQbN/u5V
Sa3HSFm858+Jnl4ypVuZiYsI723gwfGnOjj+6nDbBXSYxdTmHcPffM5/yBRhbhppgjiCo/OzGv91
bY9gLSc1VeXp65Mn3iLTxzn9o1GeVcu2lrbx7CFuugszdIpyuE8fgUxuQFH98vQh8LRRDD7lEOLB
CBfDuLZjMyBhvgLAi3T1iKguljMhhwlFYOmOyCDa1pu6qGLWLGlZ5vP3naeU1SuAsibak+vfZYV6
OlvEtnfjGSy/y6f44jE6YoLObhEQQK613XaVGKJnSHuaJ51SJUIBJJ/XhSqTVYfx7JXE3HOmqpIv
NzX2c7OxaU/rVwxPRGsw0mBal/5J6z5KQltueFB8KSZx7gLKZhWmuwg1nLypEcyV+G4zWIHuF0Nx
VeRxjWPI7VI3DPZ5d9yMhZaGVovucux2A9FiKH1nb0mR0zP8PlU02VJRUhe/dDnGbuOaGjG0QSTy
UhnXbxxLbEJqQ+OG0RitMYMc9glzdlcRC5QFFxxLwRlmVcDeEhKALuzYeZL8oiLeyzGyYGs0EYhy
mgLceWXzTp0QZEkAGIjT2ADvvtfwWG2zHF31QWdsG0sGP+g2MeMEPv9t45z+z7EbwQJXhrCKIkpi
khuFhTVP1yRcN59+sntILS+Y/AMMHG6hJXZvKhZOzSIbC2C5KpNUNEoJPD6J7ZatqN7IZjWW56vt
PULXi00FSd/o2ShCqMQswpg09IMvx48/B8BYlieon93tuiYuXQnI3gy6QJ6SDt79oLfbrsDuqrmt
6KfigE6b4CiGJTeu2+ReaP4ENgPALqAlC5QW7XyTpBgOuEVqs+f4k04cCl8zGJizDMkN6k1KCpWy
uO98ibneWC9ebZZHe+5qRj1B+Tm7+bpHWtRhrSkFFarjnA65khAkNpvDsHWYGv5nu/llnOKfzmqC
r4d1fWJGU00iVR5S+V+3KdZCovTvk4LFR1z+LRWXqD4B+AnNl6+kIqwfTFtpSYm1maNgKM4DfBFZ
YZTG0PshNW9IFcUJUKAuFz18Nn5MYzVwLl6RQAAlw9RvLzyS6uukbNl+J0yQxb8Nd4O5MFBo9Zrl
hDxLh0d9DVNwyKQJw/HnrvFn84IYR39aaIBvPhWE/dbNvniXoWbAKeo5AYi1vh0GSuv9vQ9or7kW
PuxKujaD1ZSZ6kMUSKkgPYmHh2Ct34oN5qmEtpvHT05isn61dmsOl2RK2cLdqTR4FO388k6VDfKe
L4+qhelrxcP81004MIfT08FiuTK8hqRfDqS2PGMjJ7ez9uYgt6xRlbxny3Yb/ZQDb+O4T/7QGXi1
8rXwX0ft/1G0EAj2Ig0/lbev1LM2rJ/H3OiWf5yG2Q5EWqzEyz2DFOe1KtvhbBRhLnNfAGGcSE77
nWZdHcftEtJjZyKNeiKRXN4e2Z0un6JKl5vOFsgvR4FrRzB1ezdz/5e07gKuowJIDN8Vz7lKzyJG
D6nPViWj7VwH333xRoqN0pu2fOPZ/A4pVkQu7D7VDXaJEq/AYk8jpqKTLTo+K2vFeweFBEnnTug9
aES7Ymbn6c9gNC0rQQ4+opG+Iucwaq7gSQtP37OVsI6oMZ6d9d069afBkarno2GyDf7u8e9ytVky
O/hVxxwgg8JPqKjtGyUmb21y4oUBRIXXeGTmIsYPpqb762ndWL31U9JTIcMjKaogssQDFUwV3BVi
Rm4R10Qn2GVIwIdjTyZY30Mi9BjRyYKblmgBvJAbfkVFyPNFbRujJCXK2HyiWD/MzZfRIOYTWiI/
3Q/luzO9sdo6Vane+gT88LrFZHFO0FaXrtr8fVg72b30Ra9eBjutrnGe95qZSbTyDfIqEY1Tgvij
9cAjbQG1HGSmjeUOB8yxkP9wRLbnm/O/sWr1lhiDAR5m08H84lKDNNsGSP73B0iWdPXcqY3JlHzB
cyR5ZLSIAnQQnUvKj2xhf6bvapRfLA3NrulrsgjuZq1JIqHcdTuVAJ5KOzBLSGK813H540RMD63e
QhejnN8R+/Gv7inKXj1X8g7zSG7GenV5GSMQJvXeDQusML2q1Jd00vXUpXlfd0dqLpQNYVvKwTlS
1cy6y8qcuLfaVjq6HAdoWrYxbBCoKql9ZbexWPHbxf7lapffYCRw9ant7GqdPqZ9qTFWXLl6ozME
MMe4lRDVGqY7XA56fQfaryYhbvGF3HSs0W+yOyS81vEC310akWrZQ/cX215MS9PM6X/TzJ7h7IWc
z5SIt8iHuhU+oQzw8mPUyGIkqj/BEGWVyg6jgeLdLdr0AynwM5jAyJHgQ4RUX79ucZMutCQOV92q
r+WkIi7L+Z0H7HBhWwbeSRcTLFrnt7aKo8wN+JpLLqB6/sJkye2RnxRI8hprNG6gsfPMZTSo9mkM
5m/W/RIuTZshSINOhfR2RaWa9fG6sEfQyxcsX8KUwjqt0m/C32yDvmNNb3xlNAFRfBKmiFSTfu78
rbKV1UjLgp9O1m54DSHu3v2zKiqfQWbxaGRVCsoxEUzGjm9HnJjIAZv2l1OILmH5v/uesinxy2zb
hxjdLw18XPmPbzqrbPRZ4VxdOdGRPTdUvlRTwirG9+ftNQAbuYSse4K3oRbcUfy7cNJlh/ZXhAS/
zHs9rhot3vXBEMY71xfif1gsGRAeKCD5dc/3goJOTEIhzARVFF/vZDSOyOSY5mfTZRji1LeSx0BE
uXa6w0/OAjHawyLXh/VF25FkDb9A2MqfPe7bFxYwGdsdwUxVm0uWbsAz8ecVt79XnqZB5UEk0jw8
UQEVPY7W/7yVSz3xK+rRUWhTWZ6tAZo431xqXpOX3FPvto6NFK4NUQkWrrEZEusVP6Udbal6gi6v
VpfquT+AqZGAIIIzNsDwf4ZmGImDLxOZhLdkRCAiXasJ0/XtQ78ue6LJt/Ve7HcI34wevkPL4hJq
kx/+vbUDK2nC+ostz277TFMaf3v4EzvdNhM0OcCLdvI7xj3TmfgjaJiD0wOipZCISjsnfZAAjuWq
gojgWHsGeVvfiY/KYrNjYnDdxmZipAfk7TVqnkZTuIpELeSn0Unebw1xT5wAZDw3gWAZBRUjWble
14FT+RAt5mfe/AOG0aE6LQE2+yCkqrk6Gy3JFsI3KX6cyQr5c373q5kioP8ha+6YvM6fowBqGDZl
XSblfAS5E1VXOg1dlvapnJQP0PcAGOIXXLippQwX+SQkcoAI5aHQZYnRa61E6MK/bvs40XLYEOnz
xsCOm0/ZUWXYAm/eR3tckos03jwj1i3XuPrvRZmNQSNSSdw4Oj88LJZKtRq7qwgc8o1kkqTBOpqC
ql+wr/O9k0c3oGmhwSvMqtKJUwFNkkyC9tMIFYiwUWWR7OMdMexQpqwEKaMROSYQJGHg9hWfkCCb
CsbLeHOApDHVGk1AKBHqchentkKbslIHAU+N5UtyTo9fZb3+SGlOlyeU1ZSnmbAVBQfjTwYHrvLO
zR1eqZyL++HRz/yCIJIfTJGL8TTFHNzHkYIUezMKKjIbFy63g1fCgvhNgjJBOMrLV7F6L+eLXFyY
0LmczJR4rDkvADjQ+nI8YHMjBHhJNF/L9vEoPVMQ9JV3j+RlJuZ5cvpYDKoDvkq1C1Qxskjilpfj
3TstQR6kBNJLdpOaOEHBA2jbiKK5JhRiG8XJ4L5JMiIu+ECLsMe+D7qOQHBatqQrZo360RjqqFJ+
Esg/UpLP6uabHw371hEeLwljMn7W92f1kRNDymAMWZtz4Trnzg3ZgX0LorNWuS+BFFuKHx9vFYEG
XooTKWR9iYBEs8fEtQ/BOVfa6Lg7sl9tjT6f8nSUdTK+SvuoE2qbwcmZ7ktmV+759AS5lW48DQCo
bLvGPkF9XiaFRFVWhxdmA1ZsZwnVk7n7bvNMfjxD52SX+ADpqib3eSKVaMkp0OuQ0NK9Lj93fygA
NEgldbk+cZxxhk/C3U0CeOkNIlHi5t4ohlK1HtivQd4Yt0hRyrhiq4up5egggZbQlcsT+5BTHgNP
LTX06v9fxh6zurZT94yppGchAOWDf6MQBlcYu4jtdhTVj/53ibbgia5VtdBvEl/SlzoXUcM69NQI
7SPt/XRHQP6Qg3JceTB/S9iartZopzDIYtRDrdYvRYf5Jo2IsGvlvo3xhLp7RJv+IDt9qrjwp59K
U/ySXe8z74H6+6aj4Iz0HtiIUWsY+W1hWDxd4TckFc2Zry4aWGqqa7fCi9rSjeHa9lGlvRVw9+a7
24pZtkoP6TlJZGOX2ELm2cGxyeXRpau2uk9rUVenQ/oISWDC+C/ibPXKtfblD62Pr15BtY/iI6Sm
Pf2hbYsC6c8SP7/h50tcuScShJ0Hs+A9N+kqZshNkzPfHy7wa21HOZ9jXxeAY6kEYeKqj+CMdz8Z
0HQoHXvqQvOeE53U6/XBS1lShrUv5ixb094E9H8JjiKJqmxHJ99GPqNHKjGAY4TeR9BpB+zEFqZj
kS9i2rPDcqpNblbS/b9woGWFojfP0B7I3VOgdjZDVVvhPHwBXcbhJedDQhQMePEZxMUvvC5/oh1K
reglBwbIN1Z7BkDOzxFh+5/pvixhNBUueBFPv16YGWGy+TcSms349Gjj3l6OsOouYBpd6Rzc2Ygx
+YDyWP436BeI8RLlxahWs7B2RSbfL8yQZ6zI0kM+l4e049jbZq5nre5tcgi4aCH8QCwKogwm5O1i
et+EFvKrlKyxKie1qUjY5EIe4OXytEEa157SyUQTkmNyAgnz+Rp4vptT9IV2DArUx13bXqeSzWXQ
CGqGvaG/uzib3qcY1IfgcygIt22j6HMG6Xw4Lk7JmXLVItQXs/uYipgX5j+O+REDBInhMij00OMe
DyEyHuXdGkkLF3Nabt2bawacxu9qx2lP/MW/4+as/ohT+7xsCfN8WOtuas7mqRq3HehzvixT2MoU
H8prGx4wvJNx3JVG9VNpKJtWQbwhPlwCfImH2QsFHye0ziFYlqPARVDNMI9Lb9D38VMJEODjzsqW
bXiHEto2Kx73YUSIMPvIHwAqNpNETQESnTXGCyvK65U55OPm7AwfBKji+9cyHA9FYYmMChj/H+jA
FEJcrPGHv9ZzVhr1Q33Wdf/QZ1Ybcv8pxYbay8imKBr3rlbRxthle36GAUynOiOkyT9A0v+N8VFG
XozC4sez9qOXh+JHrrsIGePaQazatbX5rEkrN0Au1WtxbShiExToc/S6PzRjhdKFP9NBGMQo5egz
Zzmub7RnYFwVJOZkuDG5O1eyEa5YMKl0QKqM76HtKK/KGGLmxfbvtPkFeN/qzVv96KfAF/eRPaR5
VEy3t+JRPPFn1UEhQ69eWxrC/cx2Ue22bYWXSPSBYqycDHohnXy67IHgGWZuYVoNAxWRWW4OTo9o
FaiFmR769rFykvgJNbl8IYz9Bs3/6c7DUuNo+9YyPAHbRVdfA5yChx5T2dJFaAjaUkJ5cMJut3K1
hjHl57c7FKow1PHRQnxW6ZuigD7i6zQTLo/npxpHpp4R4fG5lTD3uQ/Lg6Elu8FHfo8tqAG0Ahja
XqkSmc7ygupEB64zf2vMYpHHmaJDvhwOipyyFO1/7rz7bigdLz9WoF9vY1jeqCIf2qW8uVZ2R+jS
mRuwLoYuP353BJdgFY+Xc5CuptP8VycpkwoUcMmmnkaZltiDqExu8j5P9DRPtw+OsImW7WZQ45gC
lreJOoP7N1kywUy2roG8ooQ7d4wE69pud+2WpX0Qa+/xolmgKqEMl7MQNQnwOC32WpyDt9IqgTry
1jts5njqV6Kv0GnSUcfgW2GGpNnjj6IooZfhhC8l5+ukMBANWFk+5/whXE66q0agWiSp8z/tSqLw
I5ksNMEt/NP2vg7nnsmjeOKrbkRT45PceTgUQTy0V3Pfe1NHl2tELYYMoqVhiqxJ8/rMvWt27XBZ
d0vazEMu7ndnGyjoHkjt6fPL4i/HoEGsmFHZqiwAguq0jS0mAjossSIxuiPsdu8J+yUCOlx0T1VJ
NYEu19jh2gau4PcS0DH3tbm8ZT9jgunC1LrIUEPg2kBoz5bKeACfWWIW0pkFmKMusW5xm/ulJE95
IJggXnWrB3LsFkMxSLTkSRK6GU9DS5X1LfP+0RYuK0NfQUS8TQVod+LM0OE0xvJtoq0qiBScySZS
i8V9Oiz0rcb4wCx82knqQ5iPMEFr/q2sofpAEeGHUfHCilBoxIt6gvrpsLGnsV4COKYCFXQQ9wVR
5BcbPVYRdsu9JKe7M6dqyorVZRExYprI6zh61lAjSW1uXpfjefSx+iIHk5+MHMBKTnuWqnLZrSI6
AT6BNBKRnBCXN5figBP+0vFFl3VzIXCWOE4K8Kt6xMKvtKYz9uRjNKFRWJiVCtuoPMPmWpwZhIkP
A94VY/024hrbko+dl0clx3q5QX4VKsg9okvME71ev+h4ySz/5wkb6/b3vxsy0FY/K3axmR5+G8qs
S2B1mZEuSFFdHQnma8mmYCNcCGbVC2WdGrPRyXtl/A2M51DOi4ED4wlpqo4J6oP6XBDY8aM0p6Rm
Ko1cNPS24ZQM5l5WaLtTlzNG/ojEUkpIxjcwvqZNhybRLgvqq2vR2bhFl8ebdwrdBeWTShHdLD6u
OACTRHDftXSTi1qXtutn9fAp4jXf+kWv8Xif5BuIwokB/F4seaJilDPuXxLAL1b7PIpDdsOq2+8g
SPWPfbsRIe4Ms0HXvbYGFkK3d2nDxSXYg9558txAlTwf8i4FJ0vBP9CPMjBacJr4t3AAbIc8BPy6
vFpYvakMc7XbEgSgTxR82D21FIk+90xL1dATTGwBZJN3lo0+1zxFNFh4vhzr8iVVYgO29EO5sh55
q8J98EHDPF6/QCS0KwAlYnlWObPVFsXsGlNB7+I+DgU+UylbIiOydKHfYrQ1qly3ElAmx3I9dlXB
XswWYugIPQe7gI1DJuL+lUJhp6P7tl6VBSQuhXCPiMP5SRVZCms0GAFydCnyOFaT1s8VWa57RtBE
T7CovG/jpSZGNe6Wk9clgZ3dwmkW9eNcaPez4nw1a+/VpoSfS2NDk53ODSn2O3SM5RsF0N8EFtSJ
HFFuqRZ7aaX0Nhbjs8XKONJ9bhS1xwV56lsmW5ASQX1zZrei2ueP3WcS/kM4b7uYeMLbYh0aXkzc
L8ecko/QozKvAU6BelJ/Oet3MlT7PBSnyc6FkG+AuC1PeZgA0IzSsjhAzz9KsmOxrbUZj8RkzdTZ
CayrObNnp1rOwaZr2CftyOryFyR58+OorI0qlpFBj8J4W27clOy+u200CmmxBBBMDDRxEYew0+Aa
yyAhx4rh5/u2tX3kCOrdKkMG6DQUreN8K5b6UbRY2DolV3bWljdoxNKYcaU67qLc0jdcQQNOPFlh
MV/arHBRN5vEAhCGpfxkaDQk1m80MRHV66pSU24UFPDqNuDQGQ80E+A4a3WhyPly3z4yNSg+bOmE
5Qxj/bv0mG5yTDIbar2FJVhB7wkQYgySE0dAvIJf7J4W6EozNTQr1y1q+12M/dnlmvEvUSIQJnnU
5UYMQdu25T63iBzyNl1v/efGXBgn0JuAmY/UULT0FQDVwt7I/a9Job9Eg44rrhM6PnPniLGx/BJu
KagLhE6OCsGZTj/RGce3FkOYuuUE+XugcUSB9UCGl1bB+9kw7FNp4TMFPUZkpUb10JpDXb96XkRs
wTwlr3se4pHiIH4mMSzm0YWvxtz4kY1uANXzGprF/gpVb0Nv2MmPNqXASkjl952Q14KZy+lSqnQu
i+TFPpDJHwEvKMX0CnPOwBHZSCFfwSxthU/CLIxspC/8SLYlZL1UZEF1Fz9vzD5laWKEoqc+AxgE
mD1+h9QKp7+lw50xHe6Ntrw4UEPsu9r5JrAmm1YNo2E0oHXPpUGkOZi2rfKoHJLBvNJWlx2S2KWx
+j5ccmMylNVTdtp7fxUW7Nx81UxrDMXC0EGdDtceTmgG/NvaBOmihFthMtemk4Zf/n/vL17ybFBO
a3hGllBZIUOEpV7aPccDJWL/oW7Tzrt8aXGKIfSiXINe4Fd07coZIlTNf34cTN0Ybl5szNke+JWR
Y74s5l18sAIueu6cngUsGtq4FjIHVt2/1z3maV0D+eShYcTcg4PSwJQgYkLceoxTWWWjNrUpQ5Kw
1eM032heeiayG2Xzxwakm1TN4eyFa4dCYDtCrziKzIFdJgnHXiztnVCOKSvp+vroHJ0lwBvBXbqN
IZCXF8SjC6IdDxrV2YeKer/ijiWSkZZ/6Trh83/crG6dbRlt4i2orohbvFaBM0+ujKUzkWvnKFUT
wcXvL018EjzGBahMq2rzruxC+3J+DH3RgbhewdWuS6PWw+de3iu6UDb/DCeoJlJw7iEaIU/ijaTX
U6QmQ62JSsbqTh1ELmRwhXM4goNaxeunDGKhbwKqzkKn46jLOSWy8VmyNE8zthNv0hdq5xGJKVy/
wgLlvHPxVq0P/XdAsLo/sIzye4AVDWAroAlJpAFN+S+ECTC04Fgvv8mB3bpIFv6ShhYITdeIcG1L
/zHsZobh8Yj9IEmmpyJlk57nnZ/hMUimEvEZUbGfUTUrtsSvvycoH1B8D7iqINMCr5f5Fw0tZ1Cv
IZlwkLltMiPZkjw9jDxHgsAkoaGovikA2Xs5z1LK563md3VOu0wWjLvSD2+wKNA8JsoOanb4rSc5
URWaL6d5yQBG4irr09qM6aaTNepdc+phQtst4JQnvcaprQsuNhSua4JDZL7hExz9D/Ml1pBy0Jxu
Wv0p/qs+iLru7NqEJJycb+VUUpQFXC6KUMFVIDAQk+Lz/4kZwD2YpewMEEZ2gAu8PsLgSYnYznCn
0Rlb4gKpUUgYmrr6s213/q2x/o13JzFd3hP9CT2AyohLkP8KICpoR0BG/HNUdstKEmP1eiQfvxZd
ZJj5Jq41FSnEkWkD7e2bhzwro39V/DydbPzn5MRadxkpeEGWaus9fw7/QOr4dnEmIlZDQLRC//Go
PESktnUM+nev8rgy8JtPiN1O6LxkT6dPvI8/inmVnl0KHv0GCUCVVqH2Q17fox8XGgKgjoavalgZ
ouqTSGTjFOUE1Jc1VE5N+aIss0prbmEbZSyv+0My5c7hkI3XpIPl+yEUFLh6+zGNr2SBohzZ4ph1
4I47YR6OJyCrU2/SXnTa3rec8/dMN+8Ta4b8AXQ2Mma77DrV0DRP+us01WxVAzOVHfgFTDz04E8M
Y0o+PQnmKpH1Yt4QWry9IPNdfa2wtf0bEQ4S0O4eQSNrIzb2jlO2XduCJUPvi2wRNFh7cqZjPCi4
nI/VMeCjpXCviWQKv/x0pqwXcy+PeM/nYCtTyPbiE3eKCWKejq5KwtuH3leQ7/CwIw0LYlWJ7E5H
BJcvUM51I+/hnMAphpoE2diL0K2eOOP/IfrF9SVNUmeaZ8R5wKglKSTVd+9RuKuhAK9vsuLUHpf5
d2G2QuruxdnFTzpCTg1NLk3HOVfGCRLrRHb4nEG776vNyFOjKcj+xyotvEVAUPVcryV+Bs6XAtne
tfs3uI0IEnu9yGKUbO4JSCI/k+jAb6RIygM/GCdL9f/ROQRRWx1AnPj9HmQEk0ZjuwTN7apaEE7O
fm0xGplRRgI+4rrP/RL3CUGSEaI/jkQ64ZIh5ksz8a+4A6iqqCrJ3z2SNXUj63XxNSKfG/sL6wVf
pMhzJ8FtXLwhqUDplBhIWrKq4yHNnDy0iYyt/uUFr87HDUYUrw3hGJCloeWZBi+udUPSVQLFShde
oNb3nwLwq5gqQgT9Hka3IBCdr6TFH21pxyymMS/9lgOU0598Eu8SpJEIBbAW39T89NEVAeucCP/6
dJMhjuFVsWojMwTrQUJSoPsW1GUE6tGp5Mwjac3Q3jMLPJ8OSyM2Z8fvsfodtAjDUUnQfGfvKOX0
/2QmLrTmuIpeaPLkpKucd1pvtRYTQ43iLkwFxaLj2GV1T7EChdJrxlxC7jj2mnIJcssoYSCb6hbZ
1jG4EDV9dxvNXSnoI2ALaM3KXaXfwPlOtuFDZ+Gi/VQHxzDzjgpnQf79+8eD4M5e67vpr/c2K6y/
kFRjmDVZ93N017iGT4u3eCOf+kTUq2/JQbBO3ODK4vyzy7XU3BydtdPcLKpk6fPBrxs5K7ayVMcl
xGKLD1BBdRK5Q2s9TOrB4w+qcgcRfC60km3VN8x5P7qho4Z1Jp8Vrh8Q5hZd2b1fg8lXQgGNQiQW
bomAI+0G4FjqBAQVUs8TipeMPX0Hsk9KxZ9OUqNoo3vHMrGEvlddjLCoMGJZEx6mOiJ9fvFA8TnU
mRLM+Mj3uiGdZ9gVWqWyOd6SnzKk4uFAJbKb1SDxNtrQqrF111OwlVG8kwoPXFkzkd4e3bPBheqd
IBdnh1HFUZ0JLq7LepLtKzi3LWOp1wJG2dI+cnS3UtddxucCS+COsa1x1sWlT15OYtEEjk0k9LJa
7xrLG2odkIJAsLmKYk9CYLojgH9Uo1B0avI/ZiwlNFreCRnlbFfJ5KtHa7rAoTEURvwZLOMf3WHB
ck1MrIXFBFAU9WXlSXdBV7eCXlirp6D2M5NPTv3RibqIXhw6qyB0xtlrJZpOSp/p3aLoGw9cFD9t
pwrv1b9Le3bNZvVOeMICfkHYbTgYMIxTxNBGlqL+EcaVGQpN7yBf8dHRvu6sGm5kjR0+aCMRv1ZA
1UdGpOJ5PIPv54jObfvV41jbVbiOwNfhL1RijHsiFS+clMZtoM+zuunwCIWDbWmb4onM+M8Kj7ES
/4d4wGdJuKjhiBHqQsEFrtgCjgHjK1juvR/4IhjrXQ6+wgG6RD2ITmUr/tkrToTiZBx59n8sI+J2
j5DLaSfzLmKjiCSF81v4Wuo3QpfwRsiMP3yApuJhPwAVXd0jpqJt8rwEXMW+wfRhQtnpe9mrvuRR
9xg6RBANeVmuPqvDyDIGr1Vm4fEfhme8W8cwAAbNOn1VVmfBmqFeRN3UMII/7D0U0GFdldI6Z1rU
/7CERqxCUbd3T6NmgrVPsR/8cT4xW+fZ9C+l/b6RmNaMIMMKNdja+oWcKBcYAzKWap51K8EMoVyH
fqSx1sv0Hwd1HqqDRRDDbuVl2rnzbLtbjuWjEJFXMAJaQcyvsUPdSpYIOm1SowFmdCAQQRzlDINK
Zz2XCrYeYjIgnh6QMgfBIaHeZUzVhpnVXOIIR27MIgAAFO5BHIVo39P4FUSVM784lK/IKMsV+xMM
9UscJlplITgHG1yLz7vUQkKQNdv1xxXJP3lPxQs91wsSA60Kr1hkUVixSQ3bW6sD1rzQgjLPAuva
//PWGkoFeolYZ9t15rmgtud+E7V10ghCYAtJjjPbFTdTcEBh7BCSJU+MS9zgypeK4uVlGrzMX0dv
TPmjSW+KMr8usyiH5ujfdVLQRJWP+104sK3iS9b3nDjo+sCHxLHEUpA0aQjpmkto6bR9CzHRZkuH
De1r2fbT7iw++1Wk+BkTfV6ELVX9nNTERNuF+TTskMh57vKdBoubNFfjHvNWraE6YnlnmZZ4n5kX
0VZ9g40EDOsmSsawFZ8FuGC5E6Bw0Wc4hM8qWxLvpP2p/AHIpSSNiYlBJHUtQY+Q7W54YZdK90fE
/nAwbW3bE0wB1U8CyDA7YtVLUu7WUGIywNVM9JXNvVswNLoVRRTn1h3oApoJnUT/E6XgwT4TPuQ6
FzMhfZNPQUN94DH24Gh3KjCdtrRT08QxnhPalR3b9bp/T90/lx4T54LWi7NZWEIINlL8vEgQSQmj
v5UNQc8kUa9zqchoAnnAZhoXvlyQsVTJQUBiCLM3AvMJYprKAPXaP7wdYyxr7ymY33/ZOoToHJQ1
51SwDE7TkfQ7u/BQPhU+JwHeAMuqjMn/vtyy7rsqS2TxaKs38H/6gKsujGn2yrHRf3FLEEiTPu97
zVWhUsfEgldgEzyksSqXG9y6E0ZLFpiSj754cenwWVNpT2S0/QSQdCRVlYoDfyvCMh5mFUnUgNvm
mpfBqa97v1LsPaNzFxrTF2Q0weRV71M4U6+7Dp8Js+QuzVTqjGwhkCCk93KOBX3Vkg8KfOBowRU/
5rkMuqF+hTCZ78AAB/vH4bn021O6DvGDEHZ+b0tlBD1tnpKKT8lEmUrS7hgipk3uwmriuAyIwkd/
YsQaz+qcBpxwiGwB6TYf85HWkPR5HG54zPCxjh+0slboEv5GjL3N9XvHMBJUBuYp+TuZ4wo34FeK
fvMZhQ0j5EPIqh57jV6X49tZIMhTVazcU55RPma2NqbrmFjISRC4h68TaEYJSZitYNCQIRSo91VY
n6m2ClU0UPpIbudXyA+oenj65jEqDWUuxcb3V5vnyK8iT9Ltxw3n/p7rd6qkLJXtuEib3WR/KQq2
EWHMSAGJE0a+4CiQrZwCmjJoQcMKuPOcxmNeRYV6tacppd4b0UXxO9USonhI23aO++f5ixFXH3gH
+s0nREUhndP9IndqJTap4VUlK/uWwfrwpvq8t+4GJ9MlrQ+tsZ1yRKL2J1IkxGk+t/zjiLEC42sX
LM0P/HD09bmgnFLRej7JDK3OJ1Fzl3tDEdU05n6xxqKtFfJnPR/HaAj8v/rOTTFPgvy4Mz6wtkUE
+lfPx+WnXeGbGe1QKbXfulbbeWrw0gi3mabpLCC7P3aEzRp3fpmNaLEj3YuctEwshIkNJX/bnv3K
T9QvAzuWCM9plVY8CMxy4KCDqrYGEjNNSzsRMnhJ61ghLSVlr5OjK3dHbRcYxxIS53xzmSYt9IV0
R7DDglrVcsakEFp7VzDv+MQhckvs75cdIYs1+zD2yDxU2ZqR/98dJrIIDM6DK/sGWDOQr+XsGXb2
DtGhDV+q6u6m7taHQPxgzJy/KQfnlBE+1M4FhAupKFGE4TvOIWlofBRTF04jmia3w3Qm3bDnlDLJ
HUubXBMHWOREomv3lX8FBBl94Q/QTGAr8uTWiD6WSoUp0c3KzRi3kb/NeQvibL/fDQLsbKw9PcS1
HkdYw1S63GTQb/EeMc5tWjCYQhTDjOE6t4TJfcgmlUwNv64TlCAWoNgadi1CuR23Y+Cd/Rj/wO8k
UoYwJk+sSPYe9Tiy6/Mba1p1DEDHW6aaV813pWV5OMHcllxdjk7Z+9TlDDDL3m1pNXgA+DG8h2OJ
TvOswO+ZeFbTOMOYqQ1S2CvX2pB57nlNuvsZxb9Yztv2K7Ig3J9pqT3T4Lyy3uk7t0eI9UPZTqY2
nbHxJPxVCRAtxbOTvZN8H8fySNQwWGBWsfwxRULjaDxH5OBwkgtJqiBwKsjVyfPFz36s+KUDp73L
BsCi2cWsol+V7KtBatlGCAvvCUMH+nk6J4CVUqgj4gb0olxCtMrmxnCImbOgekEwmqNYLbhylOBT
t+E7cHbhYuqzj7lIpf+WnClwRoQYtxLK18kVUaylpBV1RiF+62QqRegnpGglP4aququkgykhKKjm
gv+xvpUlaPi2iUk+LB2Wy+BxFR7vUXLaeIWCIlzcU07X3yCTQura76siedlh0MYsq5k6l0GkOdSm
QvJm2zE7wU0ePQbPRt1sPh7kfoYVZk+qfPvSIcun0QoO7d4Pz+CKfLtS3wX3FfiBgy4tTAIWA415
bsoVADjBgDcu7pBosj5NJeM6pv4i2ofDSH7h2LCAc9r44mBA79ImebwIeCWoT1WPYJZASom7INE/
NeylsjWmt8x0I6enTkBBBlI68A2XoFyNgzN7uhOOX+oPS/JlACwu+du8buUxWP7TBSehHFVgL69V
PY2sTqfjB2y8d0lUFdM4aeoSj496/prfAEKOQuQWxbt+0VAwWw2MxAIPrZxndEXfE0PAbkoBNs50
l5ZMtQQP6vvGrzVIeWQ8MeEU7qhs6gRWEhfoYc1MgF29FwMUjIK6D4pAF5DiPzXWTi2zc4vFW1LY
DZ3v7sh41Y3H2GKNcouHe2/uqaraqNNITm2MsFzQaM6DG2zWDy32YPs3ha4Jt8fu3iIwZD0Weot/
ryKIqifCb2bGXXfjJEYm0No8LjRITHCKxijNHLj8Fx7JkfrsrFF0s/uuJOKhdYI5LxxoNJ/KLxZ0
paFZ+izVrr2VXo+aD+NS/WS00k2s3ApJAf3WB3mrgBUeHnMvREE5YzbUO84lytvTae7PQTt1ByqI
lcOx1ySNTKSvMv1IVVecO6UTLf2gFDv5VezFPVv7hSxbzikPgEwWL+sFJfAEIUFO6R4VMZZpgKQq
TvxUIURIObXra6yeUaVnyd5+w9OeEc57ieYzJ24XuKZSUl2ShkeBoua7CfzbY5wKgKLOaUvjiMyG
vWiXzoBV4OsZgiGgWZ+XvFxHLxSY6EkApLY7Znz+yPdiDpXEUbaT6RkmJYgKV2B8KEGEpIXZub/8
a28e1RoPOZg6GqR9q9rrHOAAeQOXEUkiNrjipat1MCUNznfa0QUym4dRmWZQ8rDfTX/JLiPP5ejN
WQd1wgQB65ww7o4vKpeR+yYKl3qONhG8A376n6qZIk3nbRBPtXDUvuEMk0kLqglojJPXX+gz/Rdv
dajIyPhlazGtEGClzhRQ4QlE0B2+BOOWjS/W6ccoANr+WdDj35WzDYOevUIS3dwzpjQFirBUSvlj
gGSfwFQieU+EAmFsC3ID4qUkblUspMI+1QPBR/j0ozeAGMzQEKivCASnjBH47huQAUAcL0uajDEz
5VWl47wAjpLGTEJ7aLPq5lDUb8aCMJ45zqx7nW/e3y3DBaP2GnXozBJalXOoMh2D3qa9gdl1ql/I
p+6au2ox3K1EV45LcUwUF/2czfbGmpA1v2DUR1Jg1Cg53PWqvfyqgsIxO3zzAPhHT4dVtIf2EmyZ
nhTcP0+RntDcWM9wg5NFq00F+pLR2a9hm8a2SsGMhp23ge/sLpuirFPdsCgAQ0MUjuBblWJQ5h0Y
jwi5fNODNO71Fsk7Ex5dmjLnesBYL3Fw3Kx2/4ZaoiHnRC0/UDaVaT74GQi/kofoqlMSwh2Nc7HB
oys17D3C9HugROS8UdTrt8ifddHwTAbtCgVYzl1E2If9CbOe5ed/6pfWzDoHvEX/sPg7ue0uge/1
pUH0dV3qj3ZPEaNmtVpX6cQR5vjli+/uzVf66673zndKU7zGkBqtUO/Mx8bZanYtzDsnOn2YdOjt
naRMRsSJkwYICj0ckXD4uuy+0V1slzMdJwSjNgcCyDEyBksPEVkuWMX3AHdLwlSx4MNRDOmOZ722
cY9E9d6MFRpcfx7/v3rZQIc8TU13hGGFG3KDs97UxOVYtBatqCEhioF8KhMLEVPsxF6mEPrO7L6x
Z00mg4UoyLwgASbwzhm6JsYk5xUrXL5B6Ob/3Hng9Ryl+E0zH8knmirEDL4Pnu3n1emzWgYcbTxz
GDpIYw9kG4TZlMtBiMxf7C2kruhdWkqoAVqx2kSRWG1514vv3Nxlyz+7u7lcp2rOHazu5EfHXFGd
Fd/p+38v+se2F/RhGiAuKD4xI9n8oSUzJarqfnyOudXkcF3w/qT8GHTn6RGOMqLvy5dS+XNQvgfE
sjygKeeJMx0dhvNAzrMsLAiCtIaBS8Ri4jOWbi6VoHZJk/a0nX61cVMwank85bipvT/8bouk2GzK
Rrx+Ea2g8H49uQVE35S59LDdqOmoIxgPDHHnK/f5V+2AANIfKz5fIvqHtMN/8EcA/1blyQy3OVOt
BrgOXr/cM3HK8WuBUQxwDTpb9OJmaHrqSY8C8vIz7IrYEhaktDOVbmv0Rscu2jCHaUWtC/ShCpJy
z1NUmS84+Jrv1Fz/axb1dEhNVGiIG6G8rggpi57rb6EAYBbpMou6vwMQwm3ZmQdFGPbSkXeNXjjF
EtcWfWfuR5QyraTnYmfaF05Uw1mT4niHW7jREgzHyhoS0gbyXonO6qA14n8SS8EThCVfRasjlP8Q
SkpGhsRaMnPdqVomUIE4wWN4+EMw4Q6uBrnsePhCYwiLHbph/VmIPoC4oVOrskxUpNnCAjeCAyo0
wjE6jBAk7dNCOE3LhxrRMXs72zc6A+v/NOakIAU/JqTnObzGNWZyun2MQRRdgtNDGqVRPfFW7G9K
259XGUsWeOcwncSios5TlEHWtCI2SHVaGQDi3INWsTG1MK9FsYlIWxqJdVMtuVf4cJynBKFk1ITY
/oaSCHJbjB52VCcLcyiOAoqN4OMx1/oONtOkT2ypy6hwwSJy07Th1fX1LP3czKd3tjlYa7VczeWW
IrZiCJQGEtEO5HqG+5TR8iFSgFxUuINlWJ14zczYCLvkEzLDPVoP3CijS+jdtOXP4p3Zd/n/QMjh
Ihh289sS/a76YVMFhXuqLxjU4BL7Urdyt1MtEt6DFPnAv0er5JFHoFOcHEqFDjLTIGkzYuCww90d
EFfJig5DOEZReGnkUllUfILHN1MyQiDbWjvQC5M5Djxtxq4mfgeWlb5Ma0SOIYx5Q25mvbCabhQQ
6IgW5kqsDn8cQMvn3347XuQrTiGzbKYd6GtOa94Nip4Mdw6WqUI1TPLT4rJfzJlYjmmI9Zqr6HZ1
WZDwdTXTP3KQB8iT0LNcm2Ov6fMc/FL0UhYuSFcCxPnFNSyFItcIZi5617Uvgfk9fDycffNmgbXU
/S+NQo4aFPegaDGP0p3C34L0KjWjByrMVssINM+5VKVXaJ3ny3M7uYWZoWJb+PREcFzkEIzUI/rc
vw07rPbvitX7PMoTjQ0KkHZdLzNbWLgpqxFPfGPMiGwhrW246ehVqXTe1p1+a5ilhKum1EEISs4z
KgrZ2xVkK9dG2TpKsy7TF5DtvybtxdHrTXlStssoSeaMThTm8Xpt0TWhgR+EL/73gr24Ho6aqq4y
Zw/ohRozQO3c1nQpJesCy4QArXNTKkaJ0/oLmynEJrr2itt/+4sQQkaoGAgKyLGyeQ1Vmhc6CnbL
evw/nXFugmDSmMYgGlXVhIrJMHvQf2aqTauxe8kkWummo9rBfh8zgpAE+qtvnC2srjcu/rr+fnqG
/0ywtD4FnxcgHyGaDK/zfk03/vJaxspbCb54APXSSOaLajLS1Vp9Ayk07ux0KciIrGku2SdxNI0g
awnq9vaBd4fd3BOagfWKkKe2YZ9lzLiO+G3FWNDM6mWzvk6KPDPfFGWhUtLVfqLsK69Ju6mu3qkE
TTgAUPAneaeMV3spYFWF94EbzaEecNJERuwd6QvRa3xVnLkr6ca3PZ1JmGXB8OLFNa5/vvJl1HR+
kOnGaxpYJYzx3ICrYFyKL7JoxnGEesP7MDMAabQ8JyzdtrupIPgXe/Gx9nJAHfoFkuVGTouwyMNH
XBisA3byGI/LB9V7gSMDr+mgdKM/w9xZbq44PmgLUtjJ51aXcOYWk373Fa9FQi2LUR3Pa2uEOaon
hT/Z9ZSJXnkocdi6Nj0he5qkwSLKz0oezJIJOOHq0ZmDPKJHA58iTN4sMISIiBLbtlHWGW+nhJS6
OkzNAy16lMgnfy7Y0h1maCxcbxLKafDFQ6dai3wKn/VtyRLFO9NHhpahS6BRC3SptvU01HE0YSon
tgi83Uchl6BORpQJUFnVp4Y4U7KA8/QUXS1Uq4xpRrLwDzGcw2JEwKIDzgG3jVI0+EJpdBqZevVQ
AgL5qFtpRvunww2x3H9/+EoFDFOJ66oFPAQ6BukWEejtUNfvuZy9JmLZv5qS6RlFSRIGbdmMhwhp
HwpdR6RW+N2Ld8wvnqERTP2rAwILQKipNmJ6MzYWi5zM8RX0ccmezB8bCiTcj50i6DcWiABul8r8
KQClhjmGd/N1tdana2+hT97LzB0j6lpc1RD3+C2MfypMNkX1tUECsYyL3WZiPWTdjF1DIRCDEl2Q
jX6x1onzcKjBPHPTkdYtMPyi4R2+GHhX0hGwnoHrMSqL+UxcOV/Bni9ql6jIjc5srvwgeVSrV1yj
HLvMYQlYmCRpQ6IjF8CnJavTWpv/aLRerZf8CMX2u5AuHegYx1Tba9PQ5SL706HUmW4ic0qwRbzV
ddfF66Tsc786Po9yif97R5PVGxv2yXCskJvXSUTkEvQARGayhBj5nGOsTBKJ0cXlCIXWpTy+73L1
AhLpsRnMLIEuDBzvDxl+ndNgt51wcYRyvMXK9Q6bFHGILcWidS63tVF5zvmsqaPASJ+62koEuYhA
G07cGcNvx6173Qh2TlgbBI6Ff5B73tj/cFbIeBpiRYjYceA/ZnXG8pJyR/GAwqizcVblT3PZlGg1
hU4htYyT9MsFNtJdF9kErFnoBcVmXdZxCe1zhForR4rSGfAEaXusAlN6vuGeLbmLP0qU1wp27Hc6
UG2y698JoMFRPh5P9biIItNxl59ggdj6SWV4/02gKwbNn/Cypdq8eIkO4ADNZpjXY8P3Z56CKMjR
XrSt+5Sk0w2RvewnVOdUnKlLptZvS16mVjW1NGJQlmboaO+W8ePVM28/ABqjAronsaG9Ro8YsxSb
OVoaE3cFbtbyzMnMz9CZc6mXCgOd1lGxlJqxiVOlCxKJF8qLIgU5yWrj1NVGeTIBrZfozsnOhZMk
PGZi1HWDT7VpxaIK6zMwjxr0sLozWl2ovNkg5ydDtcffugmF7gqJRR34xhAuJJ4XPcfEHUCwTbsS
aPU/p3siraHz+MmLDfrk1e2qpjS+jkj8h+3DV1h1s1t8d/AUT/cHQTxZXV8Y4h9ij0GhBOP0xe6d
iz2w/WLnJ1JcBU5vFal5RFJbutwhIBBxF3cOvzSBMOMS8IsqVEtpo6Ytb6F9gW6YvbC3hY1YSiok
T7YqZeN5FOGbkHuSuQ+XJ3fvDjUc9SD+Eq0eiItm7wKBpMV5aIYvmD/P99Gi9ffcncXHQcFZJkpI
RJ8emMSBjuOkyOy3YgIlEjnkuS8uGJlCFVeBQmNMFHMS8Aekb6LKweAMSsBaBaY0kHSEMoh0q7bH
cc0RggqagGdXDyYI3wsUwZytTuQYPQktSLxuRwNQxnNXYC1Oz5j1uYN04xJxbFre88kpHlf7TGlk
ytFxRD23CX6ZsIFOvEEhwCK/7lqau3UjpbhcoBR29MyyYlg8Ibl3LSrWBHfeEpD7CO0tqDykPrXG
Vqc5FN7z4+Zz4VPkt+ix6lPnCtomYPkWR8vBA2N05gcAp1Ar1QKAUsCp8anGIsYZvrZguqSm6mzl
WTZGHWLHL5o8CpQudcnFRQsTwWc8OU4yDi+6z/uLbS9aWYYu0HiXALKiitmy8hFdRri9dmUvRERf
VZ/SueolxPc1sWNHFfrQivC5oo5XLcaJauI1WP839spS7Y97XiftzNgQkekMeRxejE0nooiGh6YP
ULCH6COspP+vr4gGe894zOlzhdqTRo3kR6MOOkr5XMe5nhLhk3jZLRHERZ+nDvGtelFnKp5PeZU5
NF06F8qinGRAQ3zt0mTidkNhhK6gg4n8IqHWDA7Qhxp4qthRYTueHxer/qOswN4lZwHF6cwLIsCg
yzASA+DsOpO176g391dj7mUU51aKL8P30xO3fgndoaDR4jCdhkq63/onuzszGcYwHK4fm7mOzE5g
aQckNGglA7Pjnj6E5yAl6wV7ISa9+iqRtRvNwnf59hCFtHl20iZdc1ZGMJnP3JtD8bGGifPmYJfJ
ABNOEI/qj8X2NirF/pVlPDUwvmMeOQXs5C8Y6UcLATq+2RGMsrCeqGnb/h9CFjKcfAMPwlH4ZBeu
RDgu1wJqR91bCbRYnYX8pgyubTmT1Yutj4YL6WcQW9O7e+a1WE5YJeRvk9LXRbMwmbkiHEHEQt+F
lisv7Kw5ez3MMWoGXfO8YSE2D0OdvF99icPXKI1mlfTMAegesNHGFoiPGoUHeJiNSwGaMo9zxjMj
3pA40B4nvRT2sGaNik3fvXOquvLxrMjA2HBlWJ+04sjm9wjc91Adz5RcUiOD0X5wU0AdK9aOVbps
/vDemra6FmKfrsgNr5N6qDbEh/b6FNJeQBYNgrex1zB+Ks4pkOt6AIdAFcRBSKnA8+3ob7wkXV7H
adAVnwpZDbzFgzZ9c4jyw97QE2TmSYYg9qsaSxhcmqEKuwOyW1rf3uusiTkVrblf0RpvEYcjAilR
fDgz3iJZaQSH2AIJMfSoPOLQRmSe+GLdnXK9Z8ZeL7FGjRrYCWoYygU8OLFxPd5iQ8W9dWg07Ezj
wSjFbozaOXZug7YD4ffsDRxI03jpsxK+d2t2i83Ve1JNzz1xcLiDdXq1uoOOYHFDj3ovkMsFt5W4
Q1mzCBimWzlDgoZziID1rdiHxO1yFJgCLFV0+F3zFDXL/gGNWfznX6ABGdnvQ1RQqFQVkI/DS61f
yDlboBiU+VNFsqEYNV2demAixcUR+7NQ4DwBgoBkMXIKWKkU6PTw/wEiTgcPMwaRWzT1e/ndyrKe
XGx33SqJCNfjnbYtK2R5Qf8RXZpXGlTiCj2up23e8fN/ulGwvEUH599fEjs2aCt/KyntBUzFn5yA
ZslTVOOPemWAvDuwKZ5oqD6lRezc3wPzT1bhX707MOq219PyWMGXlHh80ZAk2/3O0RpXW6AD2c5Z
UcRntrCes0bafItHYvrf5V0OBkZcJJKjmMqZPbRnRV/Ser57OBlMCIvwg4G/cSbQaY7bzEpLWkXR
cUw7mUrtOpHrR+pzrdxR25IaNZZOsC6z0g4ZTtb+q3LHuHNf0v1tPOLBPtNbObYabsbPq628VUni
1uKh+h/RTUW4x7IJp/6j8H2fFvTZ+I9gq4EoRlh9baY+YvXPyYLPUsi/VUOb3MzbRexKWZ4wxmlg
KsDBLJ9vBIDDbep2Ez1+rqhUZtTIzNvcGHbqIKE/nDFg/dzw3IGzt5LfhpUCsGSWiLYm5HSwwLoV
fBrnEWmJmmVaxGnyTQyAH9z0/+SxRxBoGAWjbO0Lsg9dvqeVF/5DE+93dqu9UCzAVfY5wi6Hw8of
iHGljZO9n30QyOpWb6OcCc0DZWsdVtf2lBzfex/kJV70fk0pTtJzXOJk5HXNDHA4x0C0Jj/QcCjs
LpkXBoYmf4Ek/EEfDEzd9VLr6UmLiXhu8hacvUE1yjfMeMHw7i+nQzY4aYbcmkrRhFkANqIDe1bz
gE1DfwRibGDsMhz87HQCoConI177+tX8Fh7tBseycqeVLfjgtH25GOIWF6HYB1CWmlSgp/ZpRhz3
BN02dm4aW05uy0a4IcZ+jxhLZGs6ns+sOMsI4gDpjDFCMMxII7q4s3TGhWPKFJbX5ayhgmbxT++6
Hu2fiK49f8RoKWmkMSg71TN2B9E8xJERv/yki23oGvTTKIsTHlJG40KtzjOVJaUjXpET5mQZVXUg
xakQKD2XMk6TlAuZp0IrsFyUjUXBJVYOtBwIFFvaSyocKxe7p/OasvcmD1+64TbG57QedSZklsQ+
1zoDb+cIKQK+2JjaQb5HpretLs7g+j9mSWRoILJtdEeW+tOa1fItwYv5qQutUTQOAnc6PBRRNwII
sDgp5B02q8riJ7jpk496ZjY5v51SStV+RIQxG9xI/+jmg4hE1/bdOUqE9f4QZAbmGUt/JvL3m3ax
7cG/JTYlCUplAHXLktf6HpzhCX8O9F+3PVcVWic4MUF85kQ1qUC+QxYAiJLyzufROHd+ZrNeH9Lu
fETjBqSGZsbN8qeqCkH7zJb6c6azNN0hTky/10wG9Xr6YUX6RO7tQZYNUiB0WtbJCQ8Ei9hj8Yyi
595scURIeRWsfjXFQjPWEOYpAKNOmCQ/cwvTwdgqF8QIjzFDtWc9ISeeDEdujuKN7b8oE3yweqIf
HBkRCi9B6poqCsQpfDB8fT6LuPoq6V5tRmte4PK7X9sMl1kavPrVl3QbWNqicGdg1cAG3X2fX2LJ
d7EKueHlTD2cmF+PcAcHawygoGtTMM5qMd2+cOegr+rLUjJB8yrcpuZrae8uaIorN/Ojm638oyyt
EQNOhrlLON4biJhc5l4vH3ApdnQurfaD37q2ta3u0N6OwPaGQSScgthewKyVMMhpZ8MUYOKba9Sf
WawsWX8cQfbKBBJagZdWMigQ4no+wqjUDVmU47tapb2wQadmGXZC+1rFcfoC6jHEkAAGjtELtIt7
BvWyto09nvl4f9ZT4+OyhiC0KjsYyT2uV/kP5ECanyuAKxZjiQxZkZ/PdB9S5MgbOO1n4n+mymNq
YLFuLPPbCROx+hr0qI9CeZe+55gMhsZwc1Of9ghqfLrs9vWNhhtRX4ffbJ2iHZhEYOtbjwssKE2m
7myGQpS8bcx16heXr6AgfzN8bFXAc7Cpea4Ffnu0jF8TPpxqsdl2MBhRCQHzgDXMXAuSFweBTQE9
YqgRESLSOnvnV0SYiR0q++yYGxEZS++yEujSbleik0bmQomgNuiNatXVrHQxlsZ6S8BviYTBOYmx
4pcIPmSVDw8pZgV4K17Y6R2xy3K3JczI8XfTRhnbUopK4cUnYTs5QAtMjcoHHXm2L564Fy4JQed3
GZlbkd8AR7pJuA4lL+PyOW6dpA2UWE+doYjroU71Dy9Smmfs6HviA6dL+VmscuDn5kiv6Q0qhEhi
f2/Psdo1167JMiWBhOByMFwr9Fuagcf/B6v3fPn/Ia66lxkaMieqOb4FlEmZ3cif2injR3mqM7Xg
v79nn6BIVfCfrWEVSlGP3izAlF/AA1HEXuhSzZYnmHoDO1wwdiFPTxisf6uSa8j+S8acZ+W/bedR
YjLEWGS4eEHtnRcxY/PMCOHUX591nDXLmaWWXglllXnkiUPI/SjkQgvJ+gKKettTFqNUO61eHT/M
p7h044e/uuLjgiB1wGLJ5EG9mZYrjOwuKinAyQVwEE5z0W+i8dPgYPXELgpSRIVSon8ytvmoGmje
wcJKnIT6quVVOgs+M0GI54QWZzHL/2bMN2SwuwLeddGHqbZ9+Nv6DAXJIcT5EQyYFVAEdSlJlKwo
w5b/NliMp/J3rrmJdVXK+YyX4wjRmDaMK+Ocx6Zij1eRVMntnKdhAOzKohSZ4/HLC0m2UEWuHVvg
iHtvXecmZ6qfMbu73QBn7tRWHYQ/HWvN21cBpHK9ocz2HPMHu3o/UgNrbP7e1dwpvvO1u2TUYG3d
OGZ56doAyyaj2g0pAS5YJpNWffjmLLEbiHOpBCYXFNyWETukvjih/RZkVEKhos20HhN0mOrS5A0i
xMe7lOkGl/0Ko2/h3NTWTd5HInm54q5ncjinCBFGzdWcJjL/LYicysxl+oL9JuhKfQ8RV35lPcjv
53UVS5J/RN/8QStJJxcMzEU5o3H40J0lljTehN2kA3qtlY5VMxMsTgxpomJRT7HNOgNvpNrn0Uc6
YETho0jLlPXlTGTeU/QSBzDGbc9KQhL4xustZ8C3oNBORF76K5e4vYE2Rf9N4o9E0+hHb4ggfOzy
W/rK5gqB5voSpqrFk4UeTgquzoG1AGyqm5rzMyKZ6Yf/9bR5foHBXzBQzRXQdAm5gN/sMiPJvOkT
zUcyueAgsgSr3vL3oxV4MO4pHO6B08FwZSuP5K+VZWS1o8upH839rYZ4UodMuHxTEhKjhwmjdbYV
Z/PzLlWXlfY7CfoOHuBL2QuvmE90YhNAasEKkPjcRDPLDArLmJnsLVv0jHhE5jkcu0onWs523mcC
F9772Ts3u4KMi4WIoyepTuJAK/pOdRx+l00zfs0Z2BDHBuuhxRXD7OGTadU9GDkS++6NvcgUPYm6
EcTlO3VQ8L9yn28YTYZDbapZKSGtnhTv3oZxqO9eg9qQL6DLlQfJxwNT+qFqZMhBJD/IsTGOwIR2
NICvG895SSbgyqZaOa4PxpPk1Rqe2c+AuVmo2D/fCgkvDHjgiNnPzKJ6eesREu5i9MrHsr/qIfD0
RGJDC00vNayFNVyyxGfN4rOW+sGBwf+bUaTll+DZXoMAoK7nI757LBlWZY1tSyEPh0SBR5Q/4etw
n0XTkfbHn16+WtPCw5/9GvfK29jCToJ6U9L45F1vBWJ3iZoUIuEjVkN6R8PYrD34L0V2HSrdfghk
vqSbG6nugPSOuEX3Y0D2yEBy33U4K9Hx55HRhu06DpH8pebMg+RAcDSw2z+XLM2AfuuzZ5UEmwgW
pJZHpzRIBeHIyh9sD77dxBsI4yz7KCtaAQiMRJfnsyiG7GF2cSo6OVyi8/uyCNVPX9TVtk8NKVud
8+gCuC+J3Lnh3ZB1X+bWf7R5zsuSu5YZ+flRMIkHznzmDZyj0VNoUuA+1ZCRj4beGsLCCGWjAp9t
wu5Ms3DFAaB06jaukgobAZzmsn4wR7Kq0kXEOBddsjsJ/B1Uo6xsOvDLE4vI7aC2U1LFI8IND0Qy
BZx6S2AJwONKKpxLkRgiySLOrak/WRQehMz84hWxoj8fiE/5t1ocQb/qXvWrxLbtMzFwk3a1zjSz
19UqQyF9erZAzZlO2PEAf+QPui2Xa5mbx7yPuA7DfqAy8Nx3JkerIWIdECsfQ8nDW2+Uh0os0qC2
5QUQNNXeCQsz2BvrWwtdc9XFIJH68i51AJzeWzSiU+9FNPZ6XbHE8B0rhg2fXbajo36yDU9Y4ILd
W7hnKFgoExtIhDIqGd92DQo0yg3q9wLueZykErig6IOCHBrPMopYqIaCKdmCz4WqFs9enMqAy2O+
EGH6YyWfM9qpqbK1lhcCx+ScC/pp5l9lf8iyY7xu/ceOYJCVDpcbZY6EbCX44LYXVJ97z7kubGOR
IfyRHX3uzlbgAhKi+z88Zs+tovt2XWu4mk+5tuvRr9Ir1sWCXqMnJxpI7wbLW3zBf5eDSQw9pZk9
ps9xLlQdeZLOq+Hs7K7M0R2rUpIvLeV3hpTp0nQLWtNbzbZ59rDeEP2kiDlHYOwjjbbHXEGdJXlt
gQ7C5wx4+/LDnYO3bj3z22cI4dKBUYubU42Pb9cxw70cEFTU9aDVsV3Dvh7gNOgkFhZGcg+j7Q8B
4fFgLYrNzNuL/U62M2RH4os0FxA0mWood4kmxG1Wi6CBsrYkVkaducehko9bLs9OFBRQ/bxxme9c
KrUMD77bVHVCPNMnZjK6FJ17BEk79o2nH/fXLo92uR0VFjIA38kdZQWgy9NN/wz8w9L0VZUOVT7Z
MWcHUQRW5W9GNIRA+Z5z0eAifJmPaXXlttz/qlFQYpVD9XeBTLVLLdORyuekt5SZ7t+nua7AKqP6
SaCj+xhRnxmZxbN9HIO4vuvMzPSQy1Ej+PH6HU+OUEHKSX+SD2uFkGfrPPo7kwrn3NHgXEX2lFpN
uiD5bXHjQvBdHNyYOxhT/erjXrl2z8+lrhQT1u4uqittbzS2o8nIBxj/tV4aGQeVuNgwvAIq6CDh
5wcbcHtdFD9Oi4qSjLLNHgMUReF6WWPZqJ5URBRnbEaJRMJRUeUPF4yKzOfNXljwA6AmHiICJlso
cEsHayrMryGJd57eGt+e54k6nDk0tJDNSzyhpthQ98q8Vre2efKLmAGTzGLapaQ+hNUv8bTTgl4S
t91/8M1oXQovLcRdPfRxDjC+tuA3ERC0q0EjGRULPjHJcQyyspPr1UDXauFBuweu9uNb74cR3OF2
Al3f4oZO366vesReu/30NCW09Yulw24SYjwrbD1fDzmwTj2wY5MPYCMYjbNT/Ww/2bmiWYjOXrU2
OgFUNEnCuQpkQXpg7/dH3dBbgnQ+EcNcoXmy1aBJLgGmtUV8M5Kv68qe6hgjxS0UJlvK95Nd9IES
pZflYF4o7tvcoZBv9quKld5P4PiWzlxe3fQdaaDEEAH4NEdPSWdGGgMWOEMdgAn3nXryb7Xz4rnS
xi6+S9bOUBnGQgJdtiqO94BmenCQOFYxl+TgN/CWjTuK2RprqJA2ry3PyCBZyFUBHoQB73M6vyN1
QDRItrRNjklH0R2X9IrkNVeRA2HL+uNrs0wJFVKGs/ssSpU5M/C+DIg0mddPXsqNkfSw/F2oP63H
Hz72cA69rMeiU+TWEIUkwDSvsMCRb+ni+DTFd804V3z0gjOEiCQx8/WUbCb26+WnxDCaIZm2V991
0EujJ+rD8dfT2jvOClf5yGwoIPXW1I+VbOHqRdhi1k1IVGRC8/SQOc4rtokroP1su0SwUL4oOgWK
L4SydgpHKEUyLhGoLAd263hKScoL743315iR1LAEn2hPQYzCvsM7pxQGFDuApFusDmtMhEsXSLwz
lq91/xDzqm3+qC5fCKaPAsFekUA+FMJ3QMN6xoHkJ1mIWRuwyF9MiXJVND6z4MuZ2afCAC2Z5s5n
FTA2KyuNAMwZ1P7M2QGwLaEXaFsyF/l2qJwMyfwRMUS1EYSPbO0sdLiNAR1hbv5FRksuqO+lwex5
buJ7dyyS7vOgGFfolKN6DaCubvExdmB8+zLsmPhPLoQ4umdX3q3zCd+C+9p94GXOH1PNFXgf93K0
8ytLeBetMGPYTGGw36UAJGA4avmTTIE/XtAUQuxvTSyBnHzA7JFTrlR8FwVnNwRXAauTpnoHuzEG
GKpWzi+8nMaDBDPTt6uA1GoiUvIh+ZfGihbdNb2pDKQ6ah2v7E2CuOaDjr2+lIuB1fP1egi03+K7
p+6RoUUE2cErFfD3Ix1CWElfN8jd6q2gmnmJGr9Z4CRqEgX9m4dtHxITVwpGxp1BmSNFgcBOFY7g
uyDK972+z1teA2JVKb5Neo2RFB0TCBnISwyTobySLmhuiCpxrQ1ZP6N5J194ltpsrGL0pe05z50Z
2l6KvMqhgCM0eIvYNbZjZ8sEzqDvpnhdsFxtHoduRk20DUwTiu77GHkyvo0TQlC8lEHq6IOQsvLa
Z11CG9wGG1QieI4rEi7BDnwf0lwcN8hVlTwN19hdMGYEvalJ+YTbo+D6IGcSPT6a3MTsn+hOQihI
yAAxO54NdqlEC1I2J0aJP5ZqrVen+aNOCmUY8Js8USDBV9uDSa7Ancr+YjRzg3i9VKgkYOqO/454
MmH+wJkSpz72PFSnd/UAxIe++ihMXfTyXiqX0hxLRyqJbh1Lv5f46WDuee+FzcOi1nO7LVrmpbrI
9AhAddMnKHrmDT5ksUlABnadGWW5hqBay2FsG76tki5hIDq8sB8HpbHapTaO2DGEV7HYGA5rBLoi
ZMmTpxmqvHeZZL57bsoGM+i3EcrChNglOPbaJdjHhJaB5kv0rHWCLJAFxcfn7xt8khiO7nkP4DIR
BZSZPCWDpez8LRjX2TrUsSAjtFVlkTkvnPX50xgRy0/5F5xuahVaFVvc7VFrQTDpC9aBxutO1p44
cUwVOSi5p+ozQfBXfr/7zOp9OldJ0hvYpy0d+fWk3wWz/fRYGSQ1+gepq2JxhJOdd7gYKCPl/gN9
4a1bcnsX7rr835fwHWmJzeEQmwgMBdMqzlSR20pKCvrGB/hJ8phDQ/U2xK/bnIMrTJms24hiuvVv
C5M4RM8ahkL6KFfIzhBZJ+Unkg8KaUCH5SfeQkxn5uHXMbS+ihS+7Jc9HClrAOJUveZIwtieiGbr
nY20JjwI036N5pV8k0/nCgtPmUwxZX/RNN64SYO+EHTUz5+PYTzlVLbgkXLBs9Zy4YS2QCarYGYm
INqtNQVePllz6rRTLEvGGG7274Nx6fCbNfjMUGe2M/z6dm0lJpfaLjpwbXlXmUNXILMDG3GCVUx2
2cO8HuIxBuSFs1C/2/FkWEaaqVh+qRj0dxQF6B1umaJRyChxT/5DLfjG/EZkFI5NC+/trpAjCEyS
olox8G8Hnnra1DXy5MbiyY5gwcW3l2OB8Gwabt/z6WBeAYTeJcukXAzt2WsNF0Ky3ay6AU84vn1F
PcZyq3sq98+IT8rT9d7mzH6mQPu+aMptj3HK7HPvfZk8K31NHETebwr8Rc3p0n4OMxXdjWiiS39w
xhPj7vkgJi+11bT+G00ZFxXn66NlpZIRxRe9lFt0p+wsFcXbV1SwychE9GxRj4d/AR9Mn2yt5B+V
c3+YfN09QY4U0gALeLQIv09HNuxXZRgX1Om56EXEqvrOQHHOloDwzF6TnNeexCrTnVkYi7npBWUC
T6RQLPedBSuQ2MSych6O6n1pEx+4wreNph6T4cyXi2QtHXScYIHLWQ5dG5WLKCKPaqaQ+tDtvNZo
H6itR2K1vdoyQCInydZ+A1sqokL6lnp5pHNvf6eJw3lIqfgEgM1IIlyKyeqvAi2tMZpAUr+kq77s
0oHY2Dke7XtCE9ZgdyPU8CSByyG+p/T+heAVesbp7okI/ysXnq/+Vizx4ImHXH7V4HKBAwQozFzf
V3omrOMVdhESMRYAICpjP1z0rTHhl10tMZAWe3oMTJTv8Tc4Ys6DNmaAwfEj5AgJPJFK4qktKSr4
2rq8P7+hG34P33XHmKyOAQmTeESUc6yPIWsc03alZxLfr8TY6KNRK3DySfueuhnyVDUcIYhZ5402
SxRTsnJBSeXkYsVdDQgwfuS2k6QIsFBT6IPrynDI+yYHd2XtJfZ7YFS4sEuvWBBzw/Ge5GNXMxSw
H7I+8ZIWQv/cX/E4OXVIqIwtgady2/TbKKPmvNExDROr3WHyUReEwsyNQIozLNt3pdSk74z6RHDQ
C+h5NLRssLNi8nHaeJRDcWjr57e/FPC/wYmtbw25KfuyE1eYYkz+b6qQacoKYizw/8+mMiEhr/5m
b74oPUJlH2AwMndGqOvsqC6O8AVW9DYN/IMHa0ZH4pjSjX58FerpEwcwxM05W97SeI3KqawDME1g
IUSD/8YW8VAeShjW0kw96kBpC5R0ejJlaBBq9PTeRkxPHig9rx2ot7B2bPXey0OYYNNmDxPMn7tx
0Lnl7nCYLhwPDVfT9ffOxhF4CH18/mLiXGIJsQL8QxpHqAlzS9PoLzcO2G4qG3aCX1eNeP3Q3COb
FVn3isqnxuHFxHd9d0qy5TAA93HBZ+f2YaWmLK8gTtWoLyzYeh4Iva5vrcQEZOUKtt2RVOovlLFk
Ta+tL5b4ewA6RpVJ/ngv5p30UsrEmX1UfKa/bvzt1OwI4meGh197+4wKWIxjaJmrTv0rvbDyuOdu
tjxFtFwPcW5IUf3uKUzT1HnE4pXgO2R9iaWzeis0Ci7ba5H2EpBsvxfxFVbIALLEE8ScvezTotWv
9fTjn8cUi+bTU1GeR3R7p33ZdZNw1eqDGGFDX0jAJcvn4QVwp2huPq8O1MKpuBsbwMktVESadh8+
eD3r4mf3UXpK1y1b+B4dzr7craYmx++ZdspJ4oz6lrvJF096ku4WSMbycK/cwfU/Bu3CEI9+PEeV
AOFiMR/UT/k7yxqrcpYvAoExR34WGZxnxf3WEwS9P2P4MiL9HyBaK3GaFAjvPe1QwRGhb8OV6Ft5
732j+owQLGdBMh8T6ZPoGMVcxPDdBtv31mmB6G5VqX4+SSeBPnpOTQ3rmTMp1rEOFB8Pu4SthHDd
gVUMkk/za02yXKJbuhfRs31QDuO9PLNd8nqWCyj6kOf+zs8R7OhIgn1N3JFHf+gtRwrKMkv0/2r+
teRERM4gvp7DqiweyKmu8r4tjCHCl6lY8Oe7twBz/HajkH9ULOjTMWpU5fg89YYQ9cM2R7gDMrRX
4XyST2MlQvZwS3OHHdKRgCE/G6dYtcI/CulspllCiUxJO9aLwMwZVBOR3XX9kcjH4218y4kSvR1Y
Isf1vqa3gA0x6I7OiJgxgNhtoWhOnSlEQnosazSJ7CXztY4uu4w5bn/csWi9OXoSOO30nsbcey0V
dcEIYI7bNmVv38pEapuKmEYNjoqX+mQgH5LYvujcXDqRMQKXtfdAlp4/buLIzYk1e3Jyzsks923y
bAdXXX4R9wbXUMtb/bRTZAY2HS2vlmug1yWzurZANvCCIWFnPDJ1ysFuqSpgSfrxcD5F5AZhGiS+
3QoECunAENzwoljiPrv9VbRE3GBpUeu4/rTu/GtjUGQ19uSVwg3BaMQrVT8yPssNH3CgDxqC1ini
kaqjAbTAWwjEZsj1tpKttDeKp+i4E8QGHujc2XJO4n4ZE5Hl/D2VQRI5hxdSY+5rHlDbYQ42fzTs
q3Nl3rej/VpsxLRro/qwxXKgld6MUVUKtmDgRa3hdkSL/cm8zlYYwr10Wgj9A2v/wrZ6lUUrk5gD
YwXvs3W1Sr0/zQZDSalDk3poOxP6gS5uZZJsgfgpd9QPghCU1InSGE7lox97YcwMulC0pwLM7xdX
qzBCHVfb5RWARQNtZX1zxn4IoTJgKlilOsnWfGl31nV6bs/FwX9RxA1FkeuPL44SQ4ZEu6K5qoCn
Q499ef8EF5Sshr0y7/T6QIltUbP81gwyfPwDmvq32Ct8qPTyIT262aoKfyHpgrlJAhtAsIrRHhPU
JaVQLPYyAaEw+CAHhhG178L8tWXs60DyQm5lC7jIpfp6FhDjYtbeSBNJ4Mjy2Ql0DgUBz/xNt3VF
OYBUA7cb8EPDw7Cwb0ysHfjK9YwZqvYgWKsPGLJYxD1x3UxO0EzDpQstyvoWb8dnomOEZjYwSxcY
C4f+gWvbznXUGjYfvBdbed9xk2JgQ1qzhdHJdj8TtjNMMAcV6YnHlKAsa412nu8faK/eNLr52pMl
uwqlw4s9ZExxUDzdnlbeLMx9xtanZNVZ0f7t9khEbOoAbPRp8yx796Cw4HxuOBEp5GPiG2HvGb2c
pE+lPFtd+NtAg1UnRlFjC1tBojsY1CnRflOOta5FdmvondCnR4y1I5O1wzXrkW0yhUhtdZT3uEQ5
Z7BuSJy7ICrpB10Xr0l/meIMQZ0xm/AyMuk6BDGf0BmCEZtp+jzsa0Avv32+5j0oXJaghVoxfMxS
hYvp9sDSclg5Jl7RIIyFx+6OGyIysFXG+Qc1H+0ramwCf/4jsIfffHM9z5exj30FpyeFC7NKh2IW
AmOHbx9Nv56znxV+ZGzefZdfzi8s0Bk2WqqoILgptRR2Nl7NYyWjtPaYv8IIh2bPHPI19+oWPW6f
hNGaxrpA2PqN3E8PhUaDeVgkR8Sk5NPONaPdPhGO5cUCepDDa/QyypMjib0x3lTNerjMaZDldCnz
xOOHCZiBDwy+hiyleTBdOijRVzM+nfBA1OwWLBJfD1vJSF7GSP5N50eKsYoufCteJ5r256DRW9ID
xx/WddnPPA6jT8RcG46Zkngm6a2eIqifrCSnc7P3VNUlGLh0MsGaao5NkNK7OYrzlHRQhguJEsi4
I5G98XjFABQA80sV9JQ17YEgDYuZyW3CU9MHFBTpIuXqz9gxV37RfiVWg4zWS4WNoHardADswe9w
UB6NzUmiHP/TJ+/LnrKuBk/lPg1g2Tz19woonkgfy07OsaSgRNy18RFklULkRqmV71yA3Rh2u2Mw
Wjfagk45Fob9SCmLrPaIq4G2PX8g4+vWYfUU48/V/HYFV8CBbnnjYCRgCqurWCifpCNTpwDWkbX5
Wu6Rh2TsbirfR4/tcHHkFeCAL9ZPhTNSJmeTLR6KqmyMQKl3hkMw4ZlSAF5dSha64Qw0eSqneohv
dgAESMEQZm9pIq14w5bDXhT4ErifTPIEbDyGyrqk+L22Az6t7SD9OIevYdnwghXifnmnskhmrxV+
k9mkykx8KRffouVN+KgyeqvneZotokBbyB6uw0N99OoxAxdcpIYInVqklq0E83YMu0y4XOjNXyW9
dVDwBswLdkgvOlWkm8u6gC2cCXkBu1ny5pkxU2UQSJE/4xDbl52ihcifeR3BkaloY1iQzMjuHT4b
oFID7NTyVy2ji8RU0f1x9QH5f8zs0tNvJPWfEbTtc5hk16s0FpcmxQX0h92efDVB7VqZaDCD5rcQ
472/5JukZptPWvDmzmPjbLBhbshcVMZdixP+eKUKLvh3F0PqWWs5dUPSxVUNPGkuxfyuA+I5IliT
NPtxZXdaxphV9nBAEwI6Ln6QzmDWS46vGWWiwJl865j4O7ZwRVswQETDTMVR3Yl+zaxwkqf/DQ1D
v+SaoWqBH1NUFxwGVqLG/q/9TlUjkPDy3evQqQgnH6NYm6xHYfFilU7efYndoZfdFKp+FM6B+5lN
ssb0BszkGhb2QHVNC6LkDutsfFPIgXdXKZLcwPq/p5eQF8C2kDTMulFoga8RYkAIUfb5Ybzxzr53
tbErRvV7sCF7VtCFw+rrMZBxxK5e5C/2OJSU322JOLbTiu1wPoQEYAsRWOsSX6B9uwr8uzcP9cWj
soQSxQ+B/InPawJieZBfxs6WXS/bBO1QsGp4jT6E5rAp585ibSp+vHm2ZWUUW26iNX+F3oQO4KCc
d9LJiH096yW0j26bSecMlry3PStQ3kmYaCNEIKPUvDcdxgC9G2q+zxNJTKzpkyXIf3Ltllu6vQ33
Es143J7+t2wrPKN3/eRF4O8cdy0t7RGDVfzlP11mtJOOyU/RET8qpH0XqXrqTK7EmPch7y8Fne/m
Rs68sTyV9caDzI+6R1Ak1Avd6uaut6nDQMRgDEwMjvhUkcYGeRhp93jlq7lMj9OjqFNszDQNOC1P
7PHZ6Y3xO5X/AiuBenkXoxdQ/Gl6icwEBCuukP/OjRorVRCcIBtbmK1miTmikxlY7OTRhlrQ5wzc
dPbYtnXGwUDPloPg35mByaqCd37qeibonynRcnUxl1XQeL9dnL0ZDCJF5T1hQTdLRLId8KogED3V
R2+lhzB4SGTgBTH3Hnev/pJHqA/sjmyufDoEUmIzzhfJc3UfcNFZthaqh7Q2arJ5my+7oQmJIqu8
wjGP0ryZ7P6EMf0Qu51aV+7NQaaW/qmYRxuYMOgDzPr5b/7pLmMTV8JvTKjnqvwFDCNHA//7iSlv
jXdLMXPOmYkZnZtsAsN/MfHME8wZ4u6ABWS943YtM88NNwEcimvGmxEHaNxNbUsAjqT2lHPhEUHG
Z2Nc/XGkzAaLjAwnnVjWPMWMkwDGXIgm+rDMlTWA/9V+Spdf5zTljcyIL5TzsuTJ9t6G1TqhvjrP
a6yUsH79ndun+f4k6/LG74BYxi21eWLCisD1RvN1wvabEUQJJHSj3tQizK1nzmga0OUiBKI0nnh+
zLtL9E7zkNuXG1stdE7jBCPSCdLVkTWCtWXJrqroReKN1WCSDrM9sNziwjR0vnlIZ9Ggtl0/hpwB
CanPTxjQKRMS4ruteNk6ZcwbQbhxDULJ2dOZk32hfZM5EQuFm4FV0WEZHgGS1ASBY4SG5VPzcFLM
e+/XJpLbnKNO5CLA5ti0/VQ5SWzVS7HHaibAkNXwAVqW5hvJnFyYD3MnMNTlhTuLMrjhUt8SMUq1
JkmPAHXc8o1ZBkbFFTK7CL0JyL4sGxmFVKYAB7Ge3YvTFoptOMRWF6wGPdNz4kqEn1nPbtrue/bX
QAeirDgj1v8wOXnUV/SD6Beed+iduIkjF7wIYZKQlzkmT2cXMgXILEKTBP25Kx6igGygVQE1U5Qb
5FI9S4jy+9+0XhXyIN4chQZiC4vJygMPVZ5TV+2hGJOM6VcdYGnPqTehlqX6kZltICcVR1aCzm7W
truZ8MsGQdzWFEOnYMjJI+jaXLx6L89XAWLD+urPQQZM0KcREpI64z+agKjov1Qfsk0Wvzmgsq6h
HLNYqahHeIhLXh+WLmmFXKBRCf3eem4NZr68Ya4xT+6SZB/iJar43vf+BZjwmDbSMKqhmVmq3VWq
882NYSptk8duNpU8ZP8dUxrWf1lU6CbMAuntZ+kn/irarh6yzx4jU3RRt6iO6s02kLnqQ8QiCpy7
iNlWuAJv6+PyC6PRDCEmBJ7nzGP//+D8b1HjYHdX0Aq+B1KENSQO0AUfEG0U8cSWj937tGArN0Zx
mF3eCeVCV4w3l1BmNCRsK6p1FXdu2YPK6mtFOcrAlnOYxuZd56sCNdAy4ZsOB1kWFy36eu9gT4Xo
spHr6gito2Cu2LKvGCEB/ltdyqPz6MYMb8lez24Uxw7oi1AMZbov8PYV7SbAe18xnGiil1EfcuSL
Yn/Ge3dXF6XAxsD80r3x5VABkDxYCv/c03mda3d4JfPK1V+Q1bGKLIiVNxMrajTbIN6zyiRgVGSQ
JauYz5voEtEq07XxCIAVtHW1eCCoBmzpd0PScC/uyDMkckDLEb8333lVNVQ0TlGY7q/tXGqvlzrY
7ce0CtWgZd8tkldESKicBvjWwDEtqn7TiOGYksKBXi5LeLbFadFNvKMeJ8wlvE27HFPiyR4nUVCT
rs/nYR5wMpoIP/Lz+C5BRl5brrIWbSPm099WZQnjR9Gru9hM+RGNYO7fhYeUlUvhHcJ7hGDmi0ze
zPGioCPPSVDy56Cz9ZQ2qbmc9YohiD2Er0kFCzFJYV7nxugP69XLMa89nxOjPInoihdc7Ti121ZX
N+Bj+Z6ma3ago5nXjvchzahNwhfVCf7ToK1uNv688DK9EIyeQkV9ZPNz3ECPNwQTeTc0rvAhbSHo
ZR+jEiDhHX1CIZceQ5r7mreXVopeKQKfnno5q1mm4kFyQfeDWLkIm5dzlVAvB+hVDPxbNztuqDoz
6k3TLpwwKBbGr7dys+W3wdbY9XBaFwfy2XaVNj13ZEhwagqJ3N5JYM5Ixl9olCQHInx2TdCTM70m
urU4G3i9241qE1lZxcxQGGAkc6n8+Hd/cum0MdU45iw24Oshy+sAkxO4LkLTadKwYpF2B0esaJRC
wZNK7IBhga9jtJqkU0M8LVxd9J7tnpxTHg8Ccr7ITakRaI09Lzla52zOsIUfo17a5Bqe9T+e+RC4
i2BC2rwzwhcsOk5h3NQW2gLBKPUre9qCBcm3xdRT8eUs7zkGir03gA/enDmOYSYcvJae8jmFr7i6
LksPc6zN3/EF2mwAmH4ZgZwyk5Q2nAembo9bjdbTvpiMuhe4MxV6GuINNQs46rez/qG3lb9WMFvx
30K/azJgot8QcyjMR2ZdSZ0ojKfvkwDTAV/own6ja+kh3pYFi9/2Tf7FTakPq2dybZUiIoRXKOod
rtEY0kbieaGB/xSBoBGC0Mt1Ll6JzXZuQwS/cTjF/HK7HQcSk+L+VDIj3z/MVWDaC63ZrO4cJS/t
k3D6m20+U11jbfoCS2zIOxIh1PcpDdDrYgn+45hZPTpNM7Hz34taQayE4Wifes99morsSMYnS/+A
YN509kwgrgooQ7dC+ufZWzgjs1rURiwjLxGoA3z5G9wrHRauPX0XzCc4T1HHubhgKH4eQS9V5SMr
+BtLiTeyYPzd6NbDQOUM777779cHTp/tt1ipqquOAeZRzACcD3mSQ9ZtegnQmv1M6ldohfaXkIZi
JT0IzGzxpaSQGk3/FM6QEfWAO/8SYVHTF6Vi2P849H8ZpO2SpciMP1UpL3nSRWG7P06m91uK52fQ
hr3yCvoBeQQYkbWAz3qXiq8diZ7ZWAB+j9ajElnGdQ3CXlP8SJ+bRmwUeevAZbjjOIU9ZaNWYfGZ
hIp1xrOsyuMWH+KrijkkEj+MoAkKCh6vDD+6OqQvcnIc0ZhthCEJypGeOTTrNpWzqNrY272ydu1V
kOhKUGt+msUE5YlKeSxsTpBrFjKSBmThIkwJaPQb/ddvKKhM2JHPO1rJ86Af/srAW9V7oFUsCVks
s+IawNlraTC673VgHj5ihhaaKnRI6uRteGLiDVVYYXxPs68WTF/ZwLNougyTpc5ofx9j2rfvdDNQ
34GDRzTDfvCjKqCfEb3cvU5h1Ae3yRhHq4FBxPM1oVGKd7OJOH3Vll/Nfp1ozBxSVhFRghLMbfXw
MpejxYIAsNenuCogQjqUREq43kgV8d3JCfi7mDSEqOFP6/GrbhWccj7X40RsJbWmieMHmWKzOQPV
MJSigEkI7FFf8hy8jhL2bgv4zswJjFZhuxE4N9R1wza/Z0sjZB8w0Rm4y41JiFL2I7BOaojG5JJH
0WunTHqvHRkEsbYxA99CWE4x1FewjQYGR3TH8aTbD/SmK8jDoGgRqkegcObq/Y3rn6T6hBdSOEOA
Dyn+05hyr90IcmBd0rYns95zmiHMD6huaJk1B1bov/tl9kiF29iBVcRXRD+7rRxUvQNgq3zXNfUk
W19ZN2jEYEjDmNNQWf7rmTUgTMR2UFdHBnJ/2WAgTYVn+zPQv//1PkIwc7VLLF9DfSzWIJF8rvel
EM7AqXKPopW6uqGgg5Zmoa3CxJ0G/r6uWbBlkHCNw57Qg+5Js/7l3ijap+C+ygxXrp319yvWM+/j
X4zGo4xMgAEr3x1AXQiDc15PF2PejzCjXUBp1Ge2fEw7J9LO6YSpAv6gDIjunJQOGxJaacKbtZiP
EnfUISkfjxtt//XsxD6rE44KV6XdFtCzzuUhIOGsw7OWqy68TqVsS1WhB6haWhFhR/S7Pk1CmGiH
rkEJtAlsN04jehXVtevmuv6a6uhfaGGA4ESu63ln2dWWbPE+3EyMXhm8tVtTsTPNQkGmgpM7TgeT
gJxrdSzYzPGNbnQ3Go2IfvtGfyy7FGubtEUDTCsL2dch3s2KcQ4imaoSIchihMawUzRzyVIvXHdk
FLM/5NsIqtuDVgverrVbF9ONbAG6joShIkIZApnVPvwAXYSw8dp6qomEHLImo1BPntn5O8FsBO5i
919QGgbKkKJTLH146JQy+nBG5q/TiM2yxkm37H6RKgEo9GntMZl3CzQOTX0tIwCqyehWcTRi8yPq
Ar1n1jB5EHEGozIfkbU6in0Vnwy++/fMvyJtI3COiFLffuPE1dC0SGhffwW7WU05V3Kuv5blKJBF
aFqTC/Vs694Gt3ExoctmHON1qweXX2IL9sY7vCvKaY3my+VZyPC5inIrtosObeeG9Gb8kCuhQgAF
KrKC0m++QKrdS299Yr/W4VL8xyA3e5sd2HM0cZPWO6RwhUNDXMMr6b/y0eNJh8Iinkc9c7QQqCbL
1jwmKLBHY4Pboq7+5fvnLpSKq4Rh8M1lcb6oj7bsIwRInC6VceKrCao+VHv9WfrNgYf1TQTiiGJy
Gc9/GInXFo6rhpmYzpu+4J0qaJWLizY+vm+Uz34lHoG9kQokPOKvPSSX0be6K0K2wbt+V77swm7c
HxJ/3ji6MdfzSnv4IxS5igwReIzD6CNJlINHlHZPtueyFDOORqT1zXM1KpHODd9Vvpffo3Viq4m3
zdUjatQg8CD1Cgjz65Xz5RIyyXyW7FOs9w8B8QvWsYfKWqAUDFlG1nWp5RE+Rgj6KWF2hNU8FoZ8
IshQIDFYl+07O4Tk5F7SPtUmXkXm/hQOF/M5WdUxHEYT0K1V8Y5NQXB/PP1Cv6qlYH7IYN/22tud
dPvmc50Wu80Nb8T+H+XQTlj+TldTdzBtrfb1rSgQxpmuLk+SuHiWFNGI2KH6ZDzwbRtmCR5jBfag
unVhekT0AzJrv+uxW5dFRlx5CvQZoL724GXA9YvN6/3MWC5ZycJbT7vPB9KB/AoFLxIN5DxzUgAy
JSOBK4CX0PmeReyJbJCTTKmOT2MrwelqL2EQ+3JsnbwHFOhS9ID5l69wOSds00zllNPHQn3wqwDK
8vwdTS+etzzgnHKwSt7WxwRdp7yH64D6npnNqv3snU7cfN+3Q8BQj40OEZxQHWFd5C4Uk5Eo+r0T
OaSu1+7Ur9Ou+BQlaUPJ7jcz9euJG1899y43XqTqvgL/Gf2FZb2u9wCtKLmH3IqtFWZU6Z0Unal/
7qKIZas1QCkZEMWRAx7q3gbIV4FPnKe/PT9vZBliAe65C1IISK8mkevx4e1HX4RMVR8XQLhuHDD0
kiFjy53qLCgChVqWfHtT7AYx6azn9OTz2O0alG7UsiyAA5Avekq8ye2fYCJ3HWMkxZo0p0wah7zt
7vYhnb8qUfz5x3BwYv7lFU3Dmdl1I0e6YsEU8fKhVcM0Uj+SgP4nf5HwvTyvOcDqLXRK8REJuQ1l
LXcIPtD4/vWQS9D+US9FKGsFBoBF3x9jiimwOXttlYZkbjY1DukzzElgO9LmkYYCJUSNJguYnYqQ
bYa1R8zvKcubRLOhlAHNDpLeopjIyMKZigYhj4lZWMCoip3TmTQf6ov/E8lx9qleGnx8nnKA8nFd
J5AlYJ4fSlxROaug7yLcHuBsQ+qKKrcjaX03C/mfTDF8tgt8NVQ1/jWWL2UBM/4ouyZAw+UjoSsF
RxdNAE7ZXEJ6TTdDL5X8oksZkIlP+q9JGvQQHpqXKmVxP8NduYZ1PLzFUgYvLCtDAZS0+6XHxznb
F0bAdUvq4CV2h2Q99GFhAIPPd55fEn3gwkY47Q0L5UEz5zBT+chIdMpn+Jt2lNlc0KzgpCXpZGNM
OzoLUCDthabaNc8gQRqR5JtcB18R6miEDGyQ0k87ZsKqAjjELMYdlTFgheAlPwEtvq71Thk4Cknu
UL2En1/lQLgoBRda+Wn1x3g23d5fKrIWfoW9QOGRLxzi3bJ4d7Qt1SCW3PAiXxc4bC6r6ql5pcRn
fBy2nWyQNG53oEiYRCuxU+6YB7xJn9PZxk1nsB1wQrJ2Rv3lWzphiid/sTKOsLtEymeZs077afKB
YNewrfxfRwLgJqnpzyOjmOdPgs+B/foi0oe8NL8pFL/7j4T/CNpdsfBbhu+2l/SFKuYBl2nBBFz5
d8Ovn6S0LB1Lgh2DATdEDju3IWthqwcaS9M6g9fASYND+7UCwZODvKi62FhJGQE8PFli2LUoWa2I
cpLDtijohx76mxOocfIRWHFHBRzGe9l0S1zFlSF86wux/MfpvrLW1kaRT1ir5cOO4/WtxwScZgNS
ahAKSI7dNg3snnAFR5emue87juOfgCFufyTs8AuoriYNOYOAZYOmb/SORkzBZxyNNJoIF36aPLR8
aNr/8sVBZLaFuswuaG9Rkdx9RoIs06s6XXFDihZ79rAz4N5yL5uKJYb7QIrNUcn4HMWxvYqukGPx
p6X4s9gRYBMRamJFYNLzk9ELWCq2/siu8AcZe8WtNUHcsnbTOMklyS1Hh0QvNLXD9NqRW9BQmE09
5MJH3662SYbytgFTTlxNBW2E+8WwwY0t66Qy69wHOfsUZixpW4FxIQ+jTIE2EHcTND/STNrv39Gd
M/QZJV8c6ZHFSAZ3z3fckYsG5fOyqrO6P65xs8NCWHyT60H6m4gQolLV2XNQpQZnuoO7k0UqAk8W
EZq1xxVCvzRglcrwhGziIMRy1n6XhOdtiUgz+XAzIm2pfuwUmQd51Sr6nNT12ee6V1RP1dBynnER
/LN9L2Cco8xuoP5Pj380qObDmIGpYtH7JY0oYSPPxJI8ccUzKwAREVElHgJqyp2aSesEUrQTYOyn
r0BW7U7stRmUw0X6IgzJVnlFJ0qt10pLVQyfWRghRigV9NuX3DfzmKfJj+ZK3OAVpv1vEAk3K2QN
4e4b6+ApRXv8hpLMHoKA6+XSoS2hABfnvF1Lzh9pGeEt9eejV05Na6C0QZUWAlhKc1uSELaYzr0k
dX25JehzM8fp3UJoYS9C9eDI6yhKyfAzFoQ7Sm2RBOTgqLvkO4v905wCY8G9tmef4ro1QmulMvyI
IYCPkSN+vm3fVsiGDublHhi5J8ox/qxUXTw+TkpR0rJzzmDW5P3IFiK15Nnt6smi66V8Pk0y52YC
XaJw2+1mjkwBq9n5DW5QsANdeK/mOGpat2NkTjcpYvTPkGnaWnD3l8/FrLewEboXUsS1ktvkX3el
jg5ZKZ7RtfY3kCjQ4xoPIspvrOtFdiBIIJYVRg9MVgMM2Y39OsAYXiA/XnNKz7CpRXs1yFOTSEzS
HhX54lfE6t+UXSHDJwa0tA2tdtXlYHWSwHktnUv/GSlsWuDp79B+9o5eRDucXu0e11ACh3NwI3Ny
KgGWnjnRRGEfgy16N1HHxGJho4MYb0Nf7TRDLY6Kfzr2tq4wtuSgW170edj7XyPSUYIbuixOvCuw
Dm5k1X59r50peC/cAT9r5EGWXAMkQLcoOTArqiOImDx2/UPgkAYheL+jDIFkHqTcRSXxWAogJB+L
tPTEG8G4sdQsyUVN5s9h6DLA+HKbJk3jdjZcoAvNUqflXG9F88Xinas6Ci509aVzfIwB+2aHDNH3
1MQGca/c8s/KGa7Ck5sPlUzUvBidqfEgRur0DaLRNk+xljczW3KH6s8NC5LNsb8tfziBfV0EKsIo
qWtoIxE1cszQpoV4HLa0924cAXGRi5X0lPvnkBCsAz5ZAxCIfoRmO7NYDSIkfFi50wlVTY709SGH
X4/umOgjy4rKTRGcPjxL+Gbvrl0tQaOG2i0OdMvABzmEWYb68yEY0qcP7aLrUGzvrrIC/YecN2QN
H6Tw0rCkAMjq/JMpgiegjeE0jDKhS3Givv6w5p+qGEPJQPDrsLRqDZ/ChYCcNp/MrADwVf2B4DYY
hbaf8zp7uY2p9lxyUrL6JY/rHRRVhI84PSQE7zXHt/HsSeiBXNNVcEFjoVaMSRrOMszo8UUYpEbm
iUODUKfuWnLLxJK/xBavauFD2pgc9ruKAAsniYaOi2r+7pBVpYBfzpa7Zb+ofoc1zuIZYUSiecmo
5GSDE6YfUvjhLup2Jgngz95Bi8nJbomBSW3u0qSjtPoezibmJECypLED9oB0wegHjt+HCyESjJmN
+YIDFSnc3WPKzXwLM19LrC2kn8c4yD0qEWuMznRBccffXNFTCG8bSEpbiwy6kO4GbtiDSXR32QE7
PjlOxYEZMbe/HDCZ4B4ji7Ai3QG9JbPSbyigCpK/UYLDEArfQrG8pMI8PfL7QpyQQ38827wEKJpO
hujJdxSFANUtBR8etDfbTSgo00oCaffwKMHDsr2eei8VfJvlexVzdcgdEq+jMYqLjnFoLOghUGls
mpLa7OC7dnWBemAIp75S/UuM8o5h7xQrMsIvFJ9bUgum+VTesuYTyfkhk/t9/SBsc6iHTGosbk/H
S8XiyAHJZTOUPKqwJqK0mYopOeCCzmkB8YXVBUjekgzJ4DcCAhpJtDr3WERVmL8Xhi+AzR/ohuLI
P7+dlp+zO89tmGljQU6Ol4a5I2ep7GMnw4erT45Uy08LBa2M1TU+TqmHlGRKU5h+JS8RUP9f5cyC
B8httLiNjpn2fweqRXqK6D+okcFdcxFISR89Mx5aIIhm2bHKb6pXOHsOMeq6pxDlknTObTzGJyCE
dso1diZTcJE8KAwvcQ/I1YgyjVGM0ptpPUNvKy55SbbKoLOQkPekowWWGpa0gyTMnP+JKSu4xaZM
n0wSqTxOOy7bWuAUX+ze4FzUYtpQzXYj/dBfBa2/WTjyAVrsiigGP//0V1ID/awsZqM5obsNPMhC
n0UH0JVJlWomjJOBZUDdmISQod5cVqGwXeAFCdwapaVzgajc4xSGXFTy8fCWumNa/IXz773pYmMN
icdqamEd9iBRLVMtpi6wlcgNO6T4uvbigBpJ6yNJq7UhR1GsEHghXBLdo+6ZiCov0Y5P5XumnY9g
BGdCPkIw8R+hiA9buDV8AFHHLkUYY/59k0/BYiPoWSlbLLd5o+gtUxKYJWePN5v0JQXcO/PmwZfS
BOLdV9LnpqxmE6oeO0BGhsl9FUyI6JWhq20Y8/knc8jvkwFaaJPrbFwDoqfD9dXeGly4S31SHGe8
rUkUV5s69Lzu413YlKSckDcDeLpPmK96hji4xXh4HhZJhjp77k3ecLxdiHqAU6MQpdnUpx8b1yhs
ucoQquO8sq6RRxXlx7uVFuSWSoMkesoFI4Uj6XgFqRYGOyCAY2uJOnsksBEG298nmWdhEKRyk325
ZMFqYzYz0CxXU+X52QdTZAsP40eD5u83NPAACe1Xmql1jdzoRDMnuwjLAT4wBA6/eyEjcbl10yeb
qTDymKStMhHE5sETUWyRMzl2BS5elhePt0VqLnNxuHnGE6UwNzQGjASdvk0X07L8B6ZMWPUT8Ubb
jPE7WqXnLdJwqc4071xR/OxZH65A1fJ2HJKl1XmCJc/68U90vybUynmQ7qc16rnwR1jun2+dbtt8
DrsNaMABYkghamSBUQNYRRUH4uX4JtAxFkiVguiJAkA8DBbAKItgeUJJ7YKbsHH2TmNO9uiyenui
cXOR+hELPu+H5TqP48cNzBBoVMzyp8QS7Sn/JYl/0rc7jfXvm8V27l/LCmjTyy/IhSHAh+iauhJV
GCdQAWRbHg79VkL/HGdOo+oa5jFACmOCv88Gf28Mc668RU9zddpKxmJ6Mp9MHp2utjNXq5Pusxx6
o3o6q8PR2RPf7Hwukl6baH0Qn0eac18lwvTjwe2T64J+1gnemJeYZ0wYgdUXJv7BVM9FoMb9XHKT
zMSIRfD02+Q9D7FFIZnuh4OI+RVuvd4cQi980+AiEb3OLLRLXEwAQ1n7SMtO9WkOoPjb2Bv+oHkE
Xs1F+NkPQ5GRagnBkUtVQuHpS0rl0vJoI6GS0D0Sn8OedFpJSqmVyjezSZx6f39lWk+l2wDw/I7S
a0IZxx/qbF7NHdHHgXWf2FrJyffgUG7xLWQg62H4AZ3LInBrmaYe2xvAtD9RjCvcAAaL3MGOqw8Q
f9p8FbF22H47buKWf+QpyQZcn4eMBKSzhp02dbpI/BTI69x736gH8XgzA6lkfZ0OWRzpr8qjTuGn
O4H3AwHrj1LEniwP2m6E8fzXyszho9E31z+zXdCVdGknQleYz/Pn+OnDn14qEuE/WbCd36vELXT3
Rm9VLJcecHymLKujwIIt/HCFSQD0srPgdla1w/M6heReHy1S3MNT/FD0UTEDQvlyH5MD1ZOyJlK/
wB+LA2YhMq239BFYY2WeqN3vcwb6gd6De6eJQQMS3rDwEGgeqdRep09tqbee2WZXG0RxjsBqUAuf
1i+BOifd9DQul+8msoNdBCe5cvnoP4engJr6fjXtHReAviocFWG5f0ZlY8C1qutWn4qqfadKiSXh
Ywf7SwYVtGWbbNjLEmsUfVjmV0pq9abRQ2WJ3TeN7ObH+qRBcb18tfeajRDBnTRiLjZ9PS4YH/3I
FQb4czMYlsL43yROx0kD1shQdYwU6fbT4SVIj+DHfVin1TMMEGrIsRgAjtSrCX0+l7RdTj19y6nT
hISmmWZ5W//Mw9a9d/ZHks084yJGQPPmX+UroqFUZ19ALy0MniNE6UxWAz0JLyj497KHHuwQX1LW
UOXJCf9B28c277Snrz0DFMXUW5ZhNSe+GRjKNm1J+wP8bbRrFHGkJE97yNzmgC0nzSJ+TfmZF8lT
N0erkncDhQa9uDRXgF65zMSXlqywEf2hMLp/7ufDU7S4YXb0hAT6uqCiad9EqK0zN7tKAUyRG6Qn
yayZcKnr29oBiFL3Xgy8xeas3ski3kzG5Px9NzVPlXc3XvOp9nCX57HNnGBAJBuw44S/r7MZLZOK
3iORajLW+IM1IpMsAhr/Zjib3NbokalWK/RWQFA9Za3QO1qLkeFebLGkmm8912tTIx05pEW8pz2n
IB+IIGUy+hqTf17BPqivwtBqtjiWgokOaC4zrbq87OSi1aznnsiVhi4oMFaGgZUgqMxhB1ZNP8LF
c8il/bw6EYvwpNL8gqkaZMj2rQoClwAvtnILWlFA5bGjkwex4pBgt2LHb6cYIFUiI7r6aIe1vTk9
vwYFasE9MxxHEa8f8Sm9xI5Uta7HVFgzHyFBc31vEN8RfK+8Zqi2Yd0VqBbsOr4iLaiWLs3z+Wv5
LdbllHyYtXcOP0m4Ufy6/x1sjbEydLORPJzwJuv2MBm84/vFpmcjQA7f9XyU2EXVWy+8qw5Pptt2
CgV7GIr0bLLJg4n0Ls+9rb88OkMbfl+6QtTKrZ14QSXN0x9pOOtw8ymuJilZN9VlK/8eWyysGccx
e0orh9uZzm4kb0l2XbB972fsTh9je8bL3aYvBibQRNBjtkEELja+VYo6zzDdC6hEwqDp0NpBENaW
6BMBbwBXQCBD0GVGl0XdDAafPvHk0CJ6cszRoVB7WwHxF/WPZIh4kS/FsZ3kne4Mq/3XMUHQLioz
0kC/RmuCizjTrkPYrydTwS1/fwTURVROOmd0SbJfRjlKlUU9KmFlP9G5jUgg/Uou2yY6kg5drybB
hNcs0AY+NiGSyLHqAc0RR+46x5a4CNiazwxA/Ms9N3E4U5mvkA4I/8nnIwEGcVL6JGrcTy9pP0bT
hNfaub6mhl46sOJJ5AfAPX3M/kgkaaxHrMh17F1b4FaR0XPSw2MYax/JLsyRsQl6tS0Z6XoIhnRY
JbzDPJ+65rDz/JmipzOkiHhs/O3jxj4bgu/IQ1b+3SgKZZbiUtcVvquWINXQ/lathNSKTW6Mfh3h
vE0ndHjcL6WAbJHFpaa8vhxY++KjXQ3pDu8+uswXLRTlQuKFEXs/uuLvlktUhVUnuU0s95QgzCMn
p4vMVTmkkPumqc29UJBZp9A80EYCQlAbUbu8KldIi6MRF/ILBO2gjJhWkpPeo1unTj4Ivt4tKOf5
tOyH1D6mgTCh6ZlIbPdkulWdkPadDgMYYjymFUBq14vZoKr5UCIQi2UjVxLzcLmPk3JrN7fBPRmk
Vb5WGh7gXx5I2hiDfAnA5yxSenEFZxWU/2drz85N7aJWaATwsReIUA4avzucnCzdseXFhjU/4YO+
2Cg8vadFTaEdOUla9MXVJV2BXvhKkY3+Q10w8TOB2qgzt/0O/embWojiX9onbiBzkGOA76ZSBrjE
mjRSgHnsyy9KXxnddB4kthqmcpXGbD0AhH7idj07x2kxP8BWI1GLBD9LsGBIRzaKn4/1injCbJ+b
/mzTW+wpcHXwUEP4poTsB49qDX8Ci/IcJ7PrC2gQdP8mjPR4WjeNnMu5ksds3P9ygBvMgTXOZvph
1Jf+5b4SzeMqDWcU3BS2YwhFumuRbw4EW5aPIGbtbRcxYC/6Z3uVh3ChXpWDT1S19N0RPyfLtdRX
I64LkAEjpCByzMYgaEuHy9HMmLwgljaxoHzdjb5gt1GRhKV73H2Pqb3P7H21SVTY5fN5nDYB2Gaa
pA8HqELn+1M9TNU+I/uJtp07URq6YML9zQYR0VOu1ItIokirDkwXqZ+CsrtgaCZrfUolXdw3/y7G
wDgSRiTqmUABP6ZG2poOU8+aezjzo2K9BxSRunTpRt2RHImeIim3S/SOO2RSAsTSkLhZDZ7GpdLr
Lg8D8P2IOOXx2tClAd+4SN1n8WBQcgrZ4HjLb0pRHMSg1DV8CTjp451PP1CXwmkKe3Ls3PgycOzt
bhHKlLHjRQBotZxikPoCti8xGjJWNbAIv43ek5IxMhJqSqQsVt8NG4EYgG9Ssp4czRwEZnb5NhbT
Gwv24whaqM1Vsy/VxT8VSMjopBYE0YYd9QKIz2EM3H5vLxDnvfs488ZbXAot5HkYmjq0vkbdUMjW
2jQ4d1t2icXyxQvMRehYYRXNXqEYTah0Itz3MMvnwHGUPTwBACzOK1DRFFGGGhpLeBIOaSyAC9x9
6Tbq6qcX6ngpLKj38HsCY8LoqnbX+lljLTqYZa60kwlELF/BPMUE172YkDnYzVHaiHVGAfKzqzyl
k8dN7SWVR9YYWXSmOIe6Jtk/h/o7AmtAqwyCKMBadHbGnfzQtSnNnPM61E3uRYb8G0Cm1eZmzH4m
3ah5wIk5o0PhC43bdMTDLyA7O9nQoO2v6iI6tYcY/NQExAG6ak+y4ikOvqZEoxHGmNopOVJDnnzA
5NzD4cWwGeOWT1YSHctxXEtoYw0eBCFE+wDRipJQkgLaLvv7vP54zKUOK8XGqzc9D9OFjBZV43zU
mmS9li0NEietri4s5T2YFiUb6pdKjghHfh+q1WSvB4iDkEaPsD/Lpalar+EGQArT+2WIIkerqu+y
ktRQ/PLIchVo9EFcF7nxi05jg2m2vh5fe68LEvVLaVrCCf0/dqO2tj8nLhh9Rq02Jl+mrs85PrTl
zC9W13jpx9ln8MvFU+l5Jf2og2iuxNLRHoxdkrxNNy+gArkjlP3500rUvf/Q2e/QgB5AYt4oWT2s
4cZTUqciMRWiIAy4qFiohSftlxHjdqQYKEIe8Agmoj4og5RMvMO98D4aXBNHBHhbwI3zIeC2h+Nj
f57cq8uijV+7+aimrowZcfAw1zFx7NB+vS03YIMKpuovYnDIi6IQOhf4u/huTRKuQbMnGWNQgV1U
v/07XsR6f8fD6gBUikXpkoH6vPlI83PXRTbhK7rKdJGQUpd8y7zg/YDibWfohniBXHbsXd7Oex9e
AvW7y5ZoPnzrB8Ka8fu9ehW71EbLCJoSfDCMkq6r6qURanI9euSliNlIVuYCxed0AHuXn3Mf47nq
EaWsfP6+WV+qWAMDS7VMSLMkodc9NR8thfUwjN7ueQFO87MEBF+DCVxdJ8RwD+byxaMqWMZpfmJx
iRfvm9FYV5dF7/bf2cZOH5ZpqKO1POHpPtFJN6cQVcOXrcgQH1fKEYz1CpNo3W7dTs6QtIakgJ6c
C/dIaGjGMLdX7p2R+zzCv+huYHj7uDvHdHnypeMVmxI2I4xCbNlx8sdb/Rk/f27jiWJ66Kmq/98n
bhIA6ZaVLjgWpUdPlKK/A6JC+vV+4rgHly9K19+Ts8TYOjT/b3ZrvLETPHkThYp8WGQMBlKIPdUp
LN1VBYjpXaxlv3ZgAJIhyuRzueJYXZBT8yDRY8ruv1yKcA1L4Kdrh+/xvXQ6Kf+u0sjOrHDBU7zn
u0Iqi5qCYQUlpsPfVHXWEYjWDJnNtgsAeYgj00LMkRTsv5DRFBaEt1nZWpkuJl4gG73BfkOoeobC
vzQGweYnMjOfrAdbPEDpQn6sjaoeFZO6bSxDmjawIreOglF3tPOWrtdwrphAT+RDhRVk7MxhOjpF
zIYKtJ6XMNlyUv7MOveI00imp4p1M+ZrvwPFlc2LFFNIWzmtSZyWt+JHhrgc77eMvrMiFOpwd5i+
9ru+i6Yhhzn3XPX0tYu6FzI8wiiHxMVi5RHoAU7kdyceWB3qeE+dr+SfrxeSdC6V2X9koDzODQu/
M60VvPn00rZ10+9pYGXTPK3wIwA0zBYApy+ypfdsbHW10sKzUY0RG3plNUov6e0DKe0JGKijA18c
qqgFsNATA+54VFlYV4nznYxaiqUqU3hHvzSDTsyHJcRwUa+O/s7WgN4ooXXQMRMm8E9YMcdnGSqq
HT28RYT/nlOGxPt9Bn9xHn1F72ON5+1KQCbRg43mmK67xqxKjTdmp6ercKTOZv5alWBvcrc3fgrn
el17QBCwXQF3fsgZGng62lyP0sui2yL9BqleDwvlNOd1bT8mmDuNPX596EHA4aw0jqJRJLAthNUd
VfJw3/n68II79ZRoTrGyMM5ZIce0NPOdFDuEpgQxq3AqYxkpkJljNI+77w14gBUpJdZN2LGPkIxi
4rTlV9AEHPhcPWcm7aHfI6ZRs9PKsBzAZaGj+8VBuPGyfr9MkbFy++T6Rtod4Lt85F5+jmwksJi+
a1T8jkxz1RvHp2GvfuriOhACglHR1LL9z2Jql8PrJIRoVujdG4nqhMBKzxGCTSTbl0FUEUt2JTxi
DQpcu6plkwGFiMSXgl/eQCKTiTpdnBPgKO8kT279vr9dprZ3I9qjuGl5Xwm0yIrbBz+TEUZF0RR/
Uurvq5pPs6Zsncwhq+hEGn4MnBAmP3+rK8MGLLyVT0ScEQ8/6GZh1ucbncHR6zjPi6RTR47FuLlx
TRutqjFqUqXbWFbIJ5LtwGCXHqiI2+r46ccmL9opxPHoC8KGJROQKz1t28m2a0HRNoCEB+jekJVV
koQtDQFYWHgxYIEcf64hHeSytB5uPBl2ivVXvcbbZsPM9U4a7Ls4wp+aAeSZt1V1DDxUo1b0SpvP
sm+3HT1iBcxlq7qITVfaATvOkq5Ym92ALoYNbHlzMzytKq+kFMp+Ee2yM32LSwvlTc9k1ZLFQqYj
LbCxTBkoioT5eq7INZPSYZd+PE5wPWtGml91QvpXIR0he2cF3GRPDrJBI4aAlvLvf64bNnmxgvsH
jbv7BixAxE2QAtevtE15NbRJJhJ8+4SqvjPDHvURVL+iAT4xcENNzea47YlHUftX7yCPGjHTADpC
VzVVc4LElDjAfE7QhVLFgxvGkh9WvfV20cCgATAyyICFu3TquNxF0v0QEjsfPJEs/OXXUTbl44R0
RIY714SpqgXyigK//WG5+w+mgVXGLMi3ySYgPfUTvJ815lGUnzDz9IQEnh5ArD6P4PhRZCW6mE8h
09JCU6HKohp493/+KrUSi2fP/pQ9GWY3g/mCIMbVWFVqY3QgVJb7Fp0OlE3UnkRTYe2Anp2cxCYr
EyL0s6Fkv1zZY+B2fRgApaBMZVpKSRg58a09O/4SAqKnZa5UmILPpy82TLYJvq/5rrd4SIkwkUDs
n3qzUJgtOExofRsFTqjITSMkxpI6uBvcnF4YJd/DJ1xpQplzodwgdB968Ln1O2deWoS1yGejF3KE
PYqNmH6oKtozEx3S3g4BjOt1XWHh64iBDN1DdhjqZknqF8+AfU0DyjI4tIx9cXWEVpXsivRa9eWL
9Hvt5Qil2GSZNxstu63sbp7Ox0HwzMNLMJzQzbVFF4hJMmIUgul3u18TdR+/a913UNDe6cPBBKOu
8foPPjlzlWGqEt6+O+TngIZ7l2R8yCyGOI60L5/M2Wln3eoHqsiM2HREuFgtB5s6g8s0M+5friju
aCntHzXk0go0wB/uaJCX8wQEwR2LoNKECXQ+qSMh4blgdS6Xqxzq91SShfGVewl0X31tVOCX5fsa
oWYCVpIIqWwJB+8tN9JP5ANa4zzhpRQWM9nt/p6DLfFX8Nd1cVC93Fb7vUOIcEbqLp7Ih6EL9ZA+
sFUcq85RhJ5/GXtSddKEcOR3j1gekxiPFH8ArnazcPfqE3jVmblk4vw1xN/XCDuAv7JIZHIdCt3+
Ux/lRxKIYMOk0N9GgNotzy0mXQYuLgV6Ifp/iRgQvBt0PcjPuZ0rNmFRj/3Cs+0zrh5Gc8FnuG9S
2AbYTaKFSHDiAHW+OoB7ACAsJ+jOQkUlHcEmIleUHuJk0J+DXd3S+T3nnp42biq8jsb/7TH7Sdz4
muD1JOoA7c0m73pX+9MCmIEVfvLy5/k7Ytb18RCDxrtMFjoNbfZoTA7wmV0kwx+HbtryiMCs+XzL
8teXFDiNXOjPNSXXZ0hhOYZav2nj8e/xUj0xWnTGNMVlH8lqokylNN8BGzLDXFQCaG2DIS7q60ke
PxK3Tsv6qLsFvLscEfoyQeg/Mw+tyACNGqmPFX14Dhsx9YgngM7CKyWujjTguuA5XsNWN68alUVG
TYJ48lXrNGCxkTgTcS8MnLqi0FQaL41QtM/hnB026S6eoI2yPPnUhnoJmJ0zpO6i3GFxgFuwP3zN
28mQBaAGJtxy+e+zCiEVeiHllRTw+Vj0uKR5z3qknzxz1R3NNXjBBoN6Oec0bvxK6MkbP6+YU3RI
5vAqnecauS0rUyn+ysIXpACwcEQcRAEElXvmxrteGhZhx6zrLtI0L70MuyOUDtutGMYE6F5o1xvN
zctoZ/SiUBB7tOeg6TVXmsgd6zen0EkK0OwMyyLbH+SO2NF9W4QjTJfX9wQcJHvjteo9lM10IGbY
/PuYaSP1zw2hOJrNHZrS+A2oJGzCWObitGSx0iHAPWqXtUphm8diuAZc2Rbr53/XcIIwcWeV26Zb
+Q7TNmUoDqKUHh9YH74I4HJiZlfUlJ+07l2xGjbNs894LT9Jy6U3qU2EhPSmJZswhwWJEYMuMVCj
+PKTlx4rxuEwX9qibdSOuDhK37i/sLiys36QKVrZlxNag0UUGZTzZXg4kJq4xp+jeFGz+v8Adna+
AXN0kf+T4oND27ovHER3H9vg/eu+1X4/yDkWXku5x6M+05t+1DOGHM66SPKY0KOU+yJFmVqojVd5
rr/yI9kIFPLyIdOUY0/GnZy4XdZk/2abtVvMuTTMMX86XrpGI9fUJE4TvdhBhC7KT56M2gFCv+S2
Gu7jf+gZQA/tXnM7He/DfEGbqmH43iFGu1w3UDrT8utfaHpFto9k1xv6XIUReuYEExbECGwu6Nwz
P3vlEOv1iHN241hpmspg9LS/JMqIdSf1oJiLkXI06b0umpcp+C1rA/RWLM6Va5YtIL8N+8UnO8Qi
CZASNxhNpGruDPSH9pqn5ew335bVTPNnmV3Is+0R3wgfQFUgXCEZ8YQhsBDI4or5w12Fh7iQYXyy
Ig4uQZhydohLNEv9SdUPNeU7BxX3dkcdEA8W5RvSd92DXQMD16l/fe+mG2fNr7VHEuVWSnM2jsSB
y3cAWADcbGlxHEQRlbJ0q3RNSwXY8ubiNv49wJIrFzGZgw6KqK98Vq5EuV69IjBOpBC4mrRDP2FB
o1tWZgvJzT4G+Nn9pQd4JngUz5N+uSv41THk6tzlAItqR6sOS81OrIqmzZImvZMjIM5md3Bg9ezo
Ld/qlJ4qpbA/t2PJCJHAiBAZqtmtqYQpW/9ZqFHS+Uzvl5R72ea57ia6KYmhRfpVSCLUcS3CmlpN
g+QV9vaLMyoA4cVuOJ8UiFvwN5sJFje4rxj0KBPKWxPFnv/gu9G87k++GwJPXz4vZlVHjEUcwK0/
K0r3N6xg7xZucom88lKiOmB98HXBUgREFCzsMxIWMnr/drp7i1PYmuhIh4o2gew5+pEaY7fWHh6F
jPaOdAnJkhqrnVsNADaKXWcYjZ0qmYgIau71S6Fk/vIKKluI+MX+4dtwiQiq8OlUYggCD9IIruY5
eEo1PQRaO/9GjAKVFwic1Q8fpiJ07G7Rz5QwGallhfALNXVSLNw0Waa2Q4Kwm8qRLD5GmG7StI4c
obv0DynnCuSP7PGlp7N2q0bnyuCFTGc84H/WeZN0uXt4f+ZAvd/UhDVeTp0Olsvr1JXJGTdmx331
VMkdg2dzvpzIX+SmjWWkGHX58EPKw8NXZcBO9dfQsXRIavzT6v3fCoNYW80QNw707yZymi1PH/Sq
BMr7R1VdFeOpvvI9CDG9K2rerKO2VG+Y02/CzzN0HHm2aCuADzWNAbRsteXj/BzikZUDcjAe+Uza
Izty8/kxRDKmqtJN53YVdIIfjStLFMZQsu0K2IoxJlslEIQ1Ojke6cgOqzTU2ZXcbSpuL95ob4VK
m+Kh7I00ik+XfR2Pk3QxXgmYOhH2BwZatNWqOl7vdYieFGj60PJTI6xqGWD7elRM2OyThOdF57ee
dDAoG4NmNIvkALbkQkiXKnyht/afPgpKw/a+QsqJ3WhidgQWkRWTiHZuQ8aZW2fMN1jgfHBslnSv
S99Xj0iGBinRUkZrIXlbpvXrZshAwMkdYC6HGExtDdgCvlZs0v2hO49f0UwANlEsB63iJTSooP9m
Azm0o+xI9Gw0mVm/B+gXWZdxpvCKattfewyTzLmLXIOcqBOuHL1Dmq2DG6XH8xYBOHBsdDVx0+Wx
wPxK3Q+zpBNdNHl7/L38bzkF+OOITEKHktL3mQh/SL8Q+dR+hdC3MH/NX9YejMr4Mu7ooi5dK1YF
R9qludK75CNK5yijyxXWbhbYZucriGuPtYzqiBne5MQ1txUl09NnXQGrHTZXxKu7iVqi/buApSHa
Oiowb+cDkFjdEz37xaOsj4eo8dHisr+4GWDlzkY/ZlSPA5ZWXEnHicsjpxYOTH1YQaacK7re2t4P
ZQ2IRHD9c21aDBKw55zPihWOGJQRiFDn8EzMXdRronJF8P7OKQxvglCV5jyUZ9IvrPKGmbjWiddv
D5nraxt1aeqak81tnSWuBKI/D0RMC9gd9QkdB50SPINpsOgd2OI3EC0kocdzIJPSAh+3CNYXXc2N
z+ECjzdr1c877IMpP9xKZQcWyMsRYvL680w9Gok2UUtux/NO8fiNbldYgnEqF8LtaTl3ta6uRykC
9ZDeVCDWNs+TrEy+vHfOAUfIeeKEFzilhApVie19UvRSAhDSvYbdakOhqv5e2o6xlx9VQvXo9NB4
r82p/ZEABlWl+MlYRe1J4LVVbto3Z7EIYXAh55Au+JgtQRy3wVdS20w45e4jZCOpgELIGNFpiGiX
g8bCgzd/VUpcJOfvWDwcPfeY1++4ny5f7y+bU9B0nnbqzkyZGa9HXYkOx6VROhcj7lBBQLPoT0x0
jtctrjFXUaV0ttsifh1wHCq1Br/YAPZhgB1sUNsL2QJjmue/JunFKmCQuQUHXsOQ5OLxoblyS1lK
gLpSfWZJbUqwTNVc9Y/WIY5FBXk0hQHMORt0HiCyUGzX7gsw+szKf3us9zcAIanqQ6UNxCiAQiqo
vwFm83pxC/yRoUAQGDWyeQMUeyWRwZx9+gmsyzGDWJC3n+Duc5840vnVBIOmRpfvEAQzYtnE6Ece
ArIYbMzJlM3uJM3Ma4XoE+wYieb5CEw9KfuJjbavwO1uRP0CVbz/OHMrn7KHNLA8rD77U+KB+qAR
Tn3sunS3ZLsM+KJKNgBq3dbUPGRoZkQhdCIRxIJUoqjbbp51yLo7bBXotgrkZH4y1MhGsCo3NbYC
K0a2JWn1eDkARVMpFbY3WeiGkrBOuAcLIr7n0aSweieSK9uGT+R/m8A8ST+OtrV0PmBinoiYWp3C
3B5ltDWEzMk+xdL5B+xNQ0Lu8pKInixpPGYUkgjSt2ZbjSOVEGUPN9cEiwPE0klwWVZblS1mmsbp
z/gsPY5hUGxqHp7TRctHUsIO3KOrqVAi0ztrZMpGFumPHzz273vVh8vFrZmtGCY7Y87ejElX4L12
G3mPVZ6hzgWkhz4c5v1zrvNK6rNBmQgtNjDuBWjeKo1qrHXIXHICrKR2HIlvgB4j1OdBk1aTyH6g
Q6cTjFbvF9hwIVeVweGclGg52LWTEAct8HUzvhFqiZ0s6zP0Kmd+a3HV6j3L/mAJ8yVGx55zneyU
NOHDlig0rCtxNVI0CV2bSlxEg+knCdwiMtsy0BalMLeFdTmYKQiiiaNaCSQnjPYaBotP2mnEVsxP
SvQLTLbe45S0ywJxdj8CE2gpzRKOpx2ssgA6ic8Jvv0A61zwaBts8eG85QB/rGtm3Ct9ej1kxi9v
nDWaDqopaXa+6PIXuTQDncOnJMdSAwDkPtSmUN86tUUecwDhkK9sA3GRsYOonYFFb7qTpA1Z+yPN
LPesM1NcBJKiI41DFqwPby8jCPQBxdhX3RFWLnBH79y8grlbpHA4qXweJ+ryPaohFCNbD7HsMgLl
2Mcr9vfc1JDAUWNmh/211WcDGEHNlN7oAouLuhWPWNGusR74AZDww11ptcvF6AnRwcWzmWiQ/Ult
KUfQrvw6JM1jrzH/sElmPGCfNGzsQgAVkKtk4Ksp8gswFwDZByqdR61aAP2ZxbS7MKZvex50cnIC
6rdGQWJR2AugKzfBNcWr4PIptsV3DEpdFwhPTvmBgcd88CjClUjxzi9ifNCnQfL54d0d9i1KqW/H
oYB3mfStCRAgdjfJAQbW4IBi/8FfBgsXwT9nZB1AqI7xoGsdd05CAfRG3B0eqwkir9K5ZDLVNSJw
6c1oUMTCZOmVRY/KrAErZrsMTRasjk7SCpQF7H17TUz9+9h6QZb70UxX3zyeywTh9FrI6XZGgkB5
n9W2yoSAbWLMxTLER1PeYR2vNOAX8fSIg2SwGU0MdRriT0sO6CtHHCzSn8X1rWL34AYYMYWHddbM
MNH5VpBJ8D738D9amEyXnAUgZhcxo/ZnkYsNqDtNWeX0+FR0lPeW06p0s7FBtYIeaTPLZStLLV/1
5qBo/cg4/M6Gl0HuxkmhP64s4bjc7+4EIPPuf29kJW0aTGTrx97axV8IS0PaxVsFzempjAcvQzLY
2qO+Bm6pZFZAGxSRuwDUoTTEzSVZIFtOFJ8FQlpVkJbsidUg1kFXSuMeyu0Jd9Axlb7bnW+uIYH2
2yTqM1aaZwuaRuUZMJKGRjIxr6cVKHmP29MfPIk39VZ2GzaJrvuZoHRq6SLROegGsl3myNUrM6lk
xHRxSo4k6ko9GuuBqOIaNEyMYPv1IhyoCEBFLMrnI7JHDbxN14mfaZcP2fRjLwLm3LSEDdXAWZSI
fvJUCxCPv91i0vKpEX39uWUwOgN8JluAtBfESCNigER11fMe6urPJkvYpbV7Olq0TakIgcH4TGur
9lCDSA7z1NsieuGRwZ1S4F3RTizpSIKwhDFMrGRPGMqRSL4z1ZKtK75uFWJ+yAcreze5uCJvMcPT
7e3PYiKaRwGw/UffCctV1SxGDONZXT5m8k6SslfPN+YdlCwly2fHn8QQ8BVv9ydKR1rX2LF/1XR1
mXDVH1EXt+j49h0muKFREOyxwAoo/UcXnCEzU6oK3hs2AHh4/BDWkxFRLI22LCxlCZJ45rrfoyy4
rx8gHZmZqqWz4HQ2xbFOhL86H/6DVf96rzuVLllrrSOSAXDVS+7H9Den7UVoLwfww4yHbVQ6FsNh
cGp9xmoGr/er6jfxrKJJWsRbyTFLzG2pqOh/SJBX9lSAwmIj6sW/z+FFd0DVcy2Ypo20zVExDUeP
HJrV1gFA7GcKQDdjl5QIrDddGnGMQLIT3ZnVOYVfG+ixumfUKtYL0WGV41qSj/yRSYnCTX76sdn3
tKUUtUpb6EHgodRQLXiiT6xIdoMwWQIDgkqxW1Xz4n53KvO4U54HWGjsaHZPqf4rxPlIVCRg1Wve
gHn2PKE40Y/7ID1VnH/qQmK1gyNcczRyTZzIhbbYUavErZrhiwRY340fai9Ipwy1CBKJeP/Sb27k
KdHHAQ9NIhYopnQ5JpVqgMc+uaOPOF2PPh7KmiWD8gaDVW5PdeOxPwWaDpxdqMKRDcReuoUs7JUZ
h2Vro7hofV9BJnZQiJl/ixb4L/5xVUYJE8YfKdvUuKRL2u8lNx4QPsH/tPmBM7i64OqNTSQhdxo/
q4QvOyGA5T8GEi+NqKb17yr2+/baF7WPvd3G/Z2PsvPXMP81LUTjTFeGib/bNw2jociFNkleaOvr
sCND6DwRW4Pl4wHRK5GICCqcN+lBf+r690SLzAqbITuseR8rLE3Wc7RolVueEGtC9pwgJPKoYxYh
gnl2Iigm7vRADnGn2krbwPhDvKcXyiDstJP9abIf+lANMLkpAbFs36i+rnS/OFqUpUW1uO3To35A
tFIVSVKvTX4Gac4pnJqsWbZtRcyo5XZ4xK7ZYTkZseo9wRvrXlaeBvTgY/17QuQUJoYYXFmMqB3u
jIRjB4U2e+Q3UQxQgCk7n1EdnYs4EA657w7QEFMgbaKmIPhdaVAnNV+EyQaZBqWPVcfhDX6F29PD
Ogvw8md749gC0qiHiN7yDfsAgsA7tjDAJ8/g5TZ+wEMpthUroQ5eBmoNzcm0XhY6DSKTWH+fuJRF
eHpcbS7YzuxMQFHasdJUTE3tcItr0RRzz4XBlZIwkwwX+gvk9xCBLBTjrSzyLPYe4/C0BWwmZccp
XUYdLPVgbfMF0OmoV8pRsIhBV/CZT/qX9jYT3ihzmz/v/zh6Cl3uUBt2NaUb3CVzwoJNyTbzb+qB
588My4BJoqXgb3l48XToyE2GT1/JTYCva0ws2nJmcLl72dfFxOho5iZLokV7EzN/FUDyuqBhxh5C
g1xUxuCWU4wFo2Y5sZnPOxNsYwRN+6/PM+2ImMG4mBlIA/ZoIadj5q2+0ONH4SF3ZQvIaKTo1Ia7
2JR4Fun68BI1OWc4BZfuFyZ8rQ5eajzNFa0P06A+m7nm5H+W9pw7Uelhcjd/2veXHIVn5h3vyXfj
6QUyWdHCnO73z/ZrqzHlc2BcEZzu4J5u3oOjDjYQYOLiKG82vuduCpX4DnIJHHdIniGh2eVzhogp
LzFd2A8t7ER7tUuseSPA1fqQszGN9qPSFoH52M5Dsd2qRBhQ76DtXqIgYPphNc5NW8EpPT1qDWBa
fwXgkAJB+a49LbtwdXwux3A9sUX2BiBmrPrSN2PLjB6mE1NGZPPFZxGXOc2TKTf6MZ1Qb/Uj4phN
rxILUmc0I0OXN6TPUdLxWB228Xwx/lZvavrv2vfGacs4gtxGwGxErw1Fsglk6JktiDsASMlUpTMQ
1Bw+tA3+/GdkaZ0Ek+ZAkzoEmwtW8pvFNBRxv+RMSv2caklzErq2/YkNc7IYJy477qSmd+uTwE+J
xbk0WFGpZWLpYzL4YYawEnPwpZtthD7ske5Yk+pZuir/gLjQ/UiO20qPhdduds7n6Xj9p1XKp9O0
kUcE72wVhovWZux2iHdSR63IVC91PLsqmqjR70YW5tQHDUjDnfNzTBO2k0/PiWftHP9Fa9oWjKgL
ILGCfpsfte94C3AhO62fN/QWBNoJCAOmEAK6gm7n1D37Vmy5AvFO2re/EGvURtrLCTicY+/7HvA6
1BF+CL+jXIgupsrch62IRUhPzWJ5BAFVLyDrHcOLfQQ5btzy/18HqoLefyM/8njhMFMRH/l2mpSN
TgjOQT7oeI0NKGWfT8CVee6oSEdwEMl76OtnMYRuXwrSarrzi3RAEGnnn+CsSBP9BYdsdIHAOvTW
OQ1vLURsVKKnfbWeB9TionYpEXlGBdUglaby4u2bPL6zsXF8F3MdPcp14oTjqHv8Eq00llhwm766
tLY3ABnYlypXZZWnF+I7xiFl9Dk+lHxx1L1+eUNmPrtmkJZhS9U965D6xcdkIxlmukuMNxxfZKee
N8hIv3QQPwapmILswrccLGhkrME6fimJZDS07IYzv12ywag2yI2WNSuWJ/GPUBpzqW+3lHx2c9nD
WR3VRxXs4cuzSNoH4U2mHCS8EHK/3OdyBG8k1npjiiw0wPPfZyY/QycNrOQu7lo5j9nHLNsE945k
JTL5YxlhJqFlkHqmKfZG+1oNW2z1s8pb15WtWh34JM++MbMFw5j188+aIDoyF3Cnsyk4ymaR6Pak
l8qsRs9amF6Ls6ngAkGg3XkLhO0dwZ5Qhst4A+dL6bVvTcS/IAhuCzSdJARMWosbQdPStlE8t3gl
z5q2BqwsvvLxec0iVHoZ5xK4WGIEimEaZkgKJ5I6anhSzgtg2Qi1ykXv7WqT8k6unx+1kPRzq6qB
Ddph4JfMR9D0oTGqTUC/jzDnO8+Kd3aSeG7KVgYrjuOaCckS7LOSJa2OjNrlWG8aF37AFNGMUdfk
h46Wv8N9ehKrnk3eR7c5fUPaIelIIJ0xyInVAgT5wa1Vo7H36YaXSCDRiDiCFcFCjRAw+MS9XtAq
gu0hgGxgNyFEiv1ZrCNZ0jtQ74DHOSsyMeOnk+9WgNbJbKztnnJ5odRWm/s39kfA5Si4kRDe9EIH
e+pog8Gl1lc0TOccBazZLkdLo2RaC5sdkVF3tnR0BNybRT96mq0C1Kr0GnjxeQbDQF0hhD8Hi/HL
J5AuqryegbCuqQa/UpK+nEqloj+F09pJfSVepn46HJHHyD8QFyPhMx+0JLHZxREwAQVxUD2cVK0Y
zSNUztsUqoRTDEE61ys6N1jbGaVef3ATjr1VnzaoIP0Lq5oi4E9lUyPJibP30AmBRSzXr9pvkVVg
NUcyjIuJZQftc1XVNxOEiKUh5Tq9Llu3PxJ2sWSCL6t9Dflo8bI2nT83M5qlSACHvE5BinvTue/F
ej3TZoQEbR7lfmf/wQEfPlPNw6HwFNDygiDTe0bp4pdkAHy2tOzVGboRXPwzY8eRMq6x5uCjyuF5
Bho3sRNHFvrjvzP33fRo4HCesGMQd6xMrOowTRQl+d9jAghjINa2wKhPiyUQspXwZOVKmT29deOb
soZnqq5aBZ0vgqgLNRlUZMxWlqIj+l/6g6eaE3/chrdU4GewboUxyBpoz/9ywmjPTS/WbQ6iCGTV
3zqeCQAw9JbxgmjbVhnbop2T98sDbpvKROocZtA1V2Nsc2qy33iZXXOygDkZnqahwssy+HcW8Urt
EvFn4mMNijgY4nKL0VHTjztngjMQl7fF4+wq4wmZlly+89zuFl4Jjf20GzuGY+A7aASwTVhFz6J+
dn/F+UpE4p74eBcY0851brlwer1ol2K0pJQLDv/YVyKaYDtN2WOf8/32GvCCYCOR6ln1nEljZEno
JIVtCElH7THT10GnHAfEMKaingDn8CPx6cf8tGQFqiZTCNZ4NfCturCjxY1QvNClRYw4+k2Gkhrd
77FDzNue/nHF4bYXz+GtJuEv2vYNu4c+Wtrdcuw6BSIbY1tUthl1Eb4qR1OgwrAKF5FHVRnXLagx
G3bcE0dVtcW93DYnlNNf/4lv0DWsBIJI3hN1laObMN8WdpQHLX0Fjq8Iy3QqEwYFGO/YzIZ1JI5b
Q1EbPiBsxCPqc4tTU2XNtbQ9nyNx5/TKoBgav7nCH7fHjiyOmueL4HALwVIbm4isvMut8H4KfkL5
MAi40PPzZTxkkPnKfWKtODnIq7c3wlrgcumypbKLaeuAjib3ujYUOFUu0yZk9GKf+9PHdCQUe+wd
FAJMX4V1NQr8c9Etjwj64psA6eg6bxtbtKoPy7ztDKmEEoi4Fow19MFwdojrkIARn/5PdJD6fuqE
Fz1GAv7J1YssHXqG8mOeJlhy+z9CbM3MuPjs1VJm333a5g/5xPYD91NAuHuPkw7FD25m5p0xmnHH
jZYEf8GWHYkBZYV/0C+soH8WL4ZZmB72LTuKaNTnIB5UEBuUr05MrjDlYFCVA89pVz58DTTFh1Ig
W6Mbw1bhNpLFKMqUY3MOs0yQ5/mAIfis4cFGSP8BfFYBBAQl1NvxlggHWNqHmCHJeHpY2yjR28DG
GYD2lkBc/VRpVn4jOUwG54Xwa/iOGPHGOymsdulbGnmel/sJtX82aACg+OFaDDd4RCyyXYht7Wo2
paDZFugJknWMN24/YynkMMBbqXWOLvTtp2yo6dZLkC5JpfLIRA7TPz4HDtmFsGuyvlIVIGfz/6uT
5gD7MLAQyTTknuZ8BLjM+O1rzc04HJHt2Uirce5CF1d2kiViyBu+W03sCoT/nWUXsmovnUNdM9vU
1n35fHArA98gxrAU0XiqcyVntt3Fbp0JelfNW3tzHwe8Z8I+VlmoPU5T3eHEULVE8U0jobvnt3j9
UgxNyFP6+9HTIw38NvUvZ/HzspmqRJbI327SWnNxF1ROCtHWbJ8frmoQhUvvv+j7+il2s4zOaA9a
UWQHGXrqO+Qi8d7AOdNr0IhQirbwQnR8Mnm4rw7gwF2n8bzOS59/0yPmlKToaXLvDbuetzXqjOBs
B631d7Tiut8MOxl6j1mYB0o6QiaBZvSGF0Qc9WMJmBuGKj7wm1Clf2NQi9wniBA0CwhSHkqOq2V0
7lpOeGAelYTHoGSWLuI8kQGP0VAJwYEdXM11f9usIHDmzMOvDh/7SnLMRgLejnxhqdqEWkQe/Tj6
zmBlCWlk1vhfdXSApPTXUiPLHuhratMEFRjrGib8cUib2LBN4L2Ik0jNFaCy6JJLUuOV0WYGROAs
tQpHmSGjcfu+9uwELdVXwyiGyj/Xbol93pGq1YIBUrmWOGw7FjR+LbK9BHMxGqQ+xRYjZz/V7suA
zWeX+hD00jR3bWn+0C2t2oKuRp2PA6zJ2aUedbxnZmAz/wbMI8d/fSC86gSqcS2R84fkR6ixb8v3
lIhUSeMIPLvVeAeZlD3Dy+oeypFXkHjNGjo2Jskm6nzR0mFREcJdPeLsw4+XuhWGIpvPdNTFxcmA
kKb1sNk7zqEbtMesRFLMmYr0QHg3VTC0+Zj+D0pcl2Gb9+jlMPLsKgyhUziJNGtqBWZP42MUkQFg
75UmWV/FKOsXZt7eLXkntVIDWlnLbAuOWtMzfINdXo5O5VkCjUWZsLN2DJz7IEdUE44F9OuW5CEd
B88XKOvGPHqTFYpSnilvSKiqa4ODZOesi+We6+jXj3irfst9HdigGoMpyhtxVJTbzPEN5bzwm2kl
S4xGmSqdEVMdLu9s6lrEzlhC/E5CJheTQ6L3cgg8biC3THXDdKog3DdFli9t+9FG+toFdoWr0XyW
NjAkL5uZIE0QDlhv/zmKWMIeo9WsRzF+smtOxFWaDFqkat7VAc5w8Pn7nOGNI0acE7IN7MuZvtAf
PgqLEcPqlNWUP/byTvyBWJpCl9GWhpgkaee9P1yQ3eUlvE+eld6Sg1I6ZSIcyEUqOyJUyk7v+sYi
s1akuFOXlxF43YqRI5syy25+vNi35jRzIs/13veZGIJmIfvP5TpxON8pFEdJgGe//IzAOQNKw6jg
OxWpEAfWP4RhwcevT92jAKDzurA7GpYNraKxgONO/0s+1btdqvvyjsWG1gjyjstl48nRvHK6B3Tz
NDkWoDQm9UHUrBKzbqkqkojIc1cRM3SsVF2EJ37vhn4XspyRg6CmzSw41EFq995XSDx/l8Y3Q2Gd
S0bFlDC+MEcE+64EE85SW3rnPKBj5e6Iq9G0hP/5ohclnhVSw2hH90syEQi5kl1AFQudZJaseUGJ
27DXZQd0xCb+0/jpcUU4xTolse6lFR1tktbqpqEfOMkJ4S846ZRHKGd5TkVJqWtgpE2U5o7WDg3S
xFz8dB1SrBSwKyv0s+IV6HFXgUQtzIWY96tCbpHqZvymiNUoXEUtmMYcXS6pE7lOPuwabUt81DPh
2BLbis4KCmvtHu+j0dbiKwxv+lTSykB3kl/wnGZEKSaZUKutMyiG6E/DYGk3kRTcnUrHuiLbSBdd
cJs43iKv9hHiPDQw/zbavudIQ95HktEX7fdJ5ZgnOYOBCoPjHmDIAMJndQICpd6fBol7Dv3qOnWf
5SOGSSciugUmh9Q7+jEnfpqUm6Gkxtk7bMqDRp3PIg6vKyZlPK1dI+tNoaq8ZbXkmX3lEaHbveeG
jlDJfS4+zgpqWXo4vOtYGh323d2e+A4CvtzfDHJ4QK4qEMbh4Rt7GUuuRm6EuwSdTxYdobxNJI/4
+HXX+cZq8D17wseUfo6ABjOegaomefVTEFwCzlIDy9XQb3/jOvrKCDnxw80d3M33LAyncQDX3wDD
CpVpFyXFhMcvD8u3crtC3JZdqS2aMhePVhIRWBeD7lCDJWL2goYaTMRh8BV71o+JImVcRwO+/0x2
JOyyZ1eDz3Z/xBlCoBdg1q+2a4qXti5yFAqE0ciOWlSzIhqkgAsclo6Lc3fH5MlhsVaHs+19SRmu
cfx/WRlW6vLTF9hTAneLjHQEG5picp9kP7mW966Un7BlemlF3PWKkydXqZe6fbxBqzG5g3C07AiV
4Lo2NTgWFKg+qis2HXNpLd6xxtf+1xNpLuVtgPPBeXkOUCTKAs9Yr618r5ew/vP9NyVb3B3I+iD4
qvbPm5nOWv4X4N39rwIIH9hIsAkmu0sU0wQ2p/R8d0as04xC1zWG1a9NzkaMPGZQUGLAONTv/vER
UDuORCco2zRD394jkZvu68rMQemOV7GvPB9+IAaOlXdg0tRSwzDBtEzCIINck2ughGzRcJ9MqF+Y
522mAcy/GtESLuM3uBM+4sqVzmHsTULs3Ijphu+ocdZTnbShL8L36p32+XtLWHKqd92qg56v8rUD
jOmnKUe/1d7XSe+MRECXWRtTNFgSkid8iteWr5VVGjrwRs+Z81iEZzdwdDD6c/bYFXo9EKJcNmlg
1Zf79m0xEE5KbAXk4pRQns0xipLAMIEv3Kpu0/irwPL5FRNWqgbpCXB0osG/ap/zX4G8UEWJnnDX
OJWyXk8DdSO9fyTcrM+Y0E7H3khAUV4drdTtLgxPxs33A17P5VSbyw2uO95ugBHauvD/aTGDNYLu
iNS+Q4SlntCIizjAVbUb6w3hFJ37aOjf2iSpG5x9gmXRRc2tKHYFj/6ujYK9rddUyIrMxw8kvb07
qUthglG0H5vXDK4Hhpuq5VYst6/CiJgZpLg8MPpdDMggsy3kidFhMVPGVPcvubWNY9hNrfCAeCHH
CbbkyAzprwiNiCH8gR30/vVCj3H8yh1SPUKUI6dw9EqHh6N/GtLQcwt/SlmcfkIT79MmRR1iRpu4
xFqcuht0KLBDYTLuQqt/SpeG/a9zKhBcJ4q1Et1u13zzq9CAAPDM8npgAEtQpXX4u6RwAtIhMepk
2ouw5BpXHNcnqEG8x8D7mqAK1bwQTHR1DKofOQK6r+0Av8/DIvS4g7+eOPBSAEO8kXxRarwLwLYj
X6HmIMaTRQ4R1Jin2xZ0ll+MZQusYKloucOgSXDOXUCSWVz6WlibwcCbbUYT4ihZXTX6EyfAcW1g
w+0eqlDkGItqPyUpiKi2dpOgjbknDlyvBo06f2g9D+5Dmy/YEmVCGLe0wFZ2v8i33ZQ91Db7dQZW
jeV3D0MG8DeX63bfZmuesdJhmt92Dk/twcQRmb2VNJe6SaGdGH5vMIrVhQRQ/SC7i+e9itP4ouTF
X/Pb3M443GDwHXxD04ZAFf0UgnnZbTLdt+aQulyma0VAnM0bl3nbxUCHjAzN18ihInCNo7dgR9MH
eL3yvAdHimyfE0asVfkJ1CLlvnsk2TqFlnwZv17CPxUjaX05+cUXQOM5yoGwRlFjXFdzFOvPVPRc
2jd4mNpN/i3s6BBFfXcdV/+jS/rKLGVeSj1353/Q5r2FSuxcuPgNNrz32bhTvlLqBiNGfnKtzygV
KwvA/dKG8r3Hoz2nPZrufOzPKOJX9EYL3TnGi1UL1FLmOCpR8DMPXRI4cSU/ykrxHVq7aSLFRks0
kboz9KEVVyUM6N6Z8t8YdyaIuyMRvRZ/L1SY/y0/U7+p/rZZYNJ6ZvZgV0dQzWogbK0el+KdFoKb
fh/N/tIKBQTwbmMMpLrvpmODDaxuQZkkxXtvALe1aM+5d84x0djpbuwuN6l/KNRrRR1EdDIhhlZf
CKPWpd1S0MkHtL2CtdPgBaQNevX6urgsaZg2KZZlLJXCAbNVmsrFE148g2DO4/ItEi/D+Ibf7rSm
nwk/IxhRgQFcQBw/pYAU5CoL/zQ0ZeE7cYJjzZ4NphcMfha3/3mtQ9TljMXY9d7vxm9O2jM03gTP
YYf7L60lQD2lC01qMOEyPgd1IGUJMzmK+EOZB3YdDNm6dvbqCCVeC7em6NSefLBkLcqAhyxGGu0f
wFfQsv15vdzTsUPGS5PtLShZgp0tdfbOiBTf/lyl87kV+Xow7rSh5/sILHjmuIEkWfo7xOey6xLZ
l1+1QjTuQtkvU/3KsL+EpCQ+SawAVncFYS4c7xDuxWI1KFFMq97zFh6nnrv7hiYbvxY/Kw90dKBJ
peL1YiDc6Eth0XoUwbXIkUAgrxF3yKxjMVaRc+2/CUeCWmqE8l6OgYoBRLKHvsa8IkMetpVlYuJ1
8RDHCgxAvJ3ErT5R4oL73hYnf04gKStbcDgxALikvqBBGZQDfYEViyPl85s76t0iPC5LIix72XJQ
Eqo7AebU9l7B6Yny17xFlnYoKs0eF13EGirghnx6GmEnXm7fW8LCHjwamNEu3MtECd7eDu8uE7Cr
7dM4t5DMec0tuvq+KQnsqtt/seqxnhjm40cttUzg80zkjF5EN8n+nfMlUiaQvqcPXfQiwkjSODqR
+Z7EEdez05MfTLj6wlyA+xizqie0jf9/YoXv4Jqzmgd7164AxmmpHGTw8WCIo2cvlD5mOhkY+VdK
szRV6JoaFvB68LI6EruMIMMFOLVhiqepwclyVBJuHk5BZrjRhDcAtnqwaB9OVhL7aH2IO21fgp1Y
LbNbh5xnQ/nGfteLBkLsP98Aot/3ppck/suLlUTWfMcLTVERJgvyYUfpr/fl03lUrC2+cEsQSVST
r9vPcgCA5FNPEWKhYH74HYXZ4Ktq6EuWwD3N4C375PG3oOso6XoQVskco/TzJaVqLJJj4VZtbsCL
tZjELS9C/AD7pq6K1m7gtSn2DsGghJ0I0VEOHYTn8IFvRGxf8ebzuoBxo0OvjZVBnHTPW2vaNJNL
jnP8VxDB+zhDKmCzknVUAi3MmS60H+UnngLDV67G6qkAL78erUhV8jNH0qoQbq3yJOqk2OLCRfu9
nqs1r07K8gX4BSS2K1e/Ky0eUUFo7UtK5b8xKpk7RSp+WO//2gMNG0JI+zYO9fbzpgn0vrRFMK0G
x09UyZ9ZxVE4NTx58v6TMUjC4906OvdEPFlNI4eX+5G2+Wrppy7tWB8gDFsXSyPt3OOSPn4A4OQy
qp/GTSrh+cqXoHyqZCiETOPrTuDMr8N0HROla4E3wQ80k4AKqqONtxXQfjLSVX245QMMB/SKnla2
wCd6VQLfUnSllNAL+PflhiK8fSICTIXZJl5ndYDosWR4qxnZ0Tbo8oFhLhl+EEmrcEh5qgOxHhXo
xgQoktxnWaunps78KTHWS5TPNocHZ9fdZqdUIA/saecpTY9FoPothasrGFtkUHMRejZ4WJiJYyYq
7owgUtqMREZBTDEI1E2Ev34iad21+HMRYuB5HGI15kKa1ty2+BvFbi8vj933mB9prF24E8C3oFdI
rjL0LMZ0U/QCaov5vMt5xZ3gmr94Cbf7pmpEVp/jPHrWy3mdHROx2h6DMpXinaLg+Hzm5M47/e7x
VM+Vz0eHNeOsHC9El9rl6ayv1gyhjI4phiotOPspTrJ+l3N9wln45zZyOvT/Rs7+BYVpYJijT+AH
EVDRpZ8dXsAMhOp89ILXsGE9C8rOlVMB/kFzAAIQoCGW2bUIRdvcZvjZ5hObrbW3ao2z6clVSI2B
DFKKs+7+M0QSuKdfMl4BsWX5wu+WjKTcIhZwN0hTCJHGlXZ2Y+xyyd5FNwoP1sRsUb00zmUgfJKX
DicYRYGXIvnA4qSlM6IC8ku7T5dtMfeJiHE6sZWeiVBqBja86iV5A8eSOgae9reKR7X1lpo5TJNr
PgJopaz3QGMk7SEUFEAqyW6+/qze3QkLAzHx4SrO58veVARGRHBoFty136hIZjaCaT0ED/MFjwkG
A7PAv0S6j6eAZ3X8pqZrrI6i8A3NNAX28FrE4hJCdXWGpJsDZoVjlGoyPYNlSIL4ik/yO7n1cZkn
2WPRSJjmKzQIchZKkThVXIqPMJivTD1+bnyGPNT4PTM6QM0ulmxjOaPaAGJXLzV1aJQ2bdPm6O5u
z+UUyGQXMUthQ7w9lg6jptdovdFsOj1FWA0cU4zjrUz6326It4NBIJoSuQFnBR7E6ETRAqXgIkYL
sT6iQ4np5AmiTmkHy2pbzxxWGT8nhCgUHsypcVAkF6yJ2E2LNecXn+xd6u+YIa6MaRqT5aQxLSGj
jl9Xc3PDrcbZvya0SkFbHHqYfXIqkAWA1xbkBJjLJ9c/DIKQMEmGKrYxCRFAoPEKfsLBV5aE3Xiq
4wQPDshS2ovdYxvHm7kMRWaUOhgAVNqm4fypXdjQ9ITUeQ70nEKlhhJj/jhsqDWt5nNUfDeIzcNM
FBLv0xAZzwYAUpukJXThMQ2lHGS7XlENcO/9Uu+FQd2FbDiRcAuG5L/XJkpzIc1DQKuEMc601jhr
Np/t2lix57nHFh4RFT5+OYeSk1puL05M735rbzPOkNHhiePIFzaEDybNe9d9UzDiYSBVlORxmYYi
4HWHNLAVEyXfEMJH5xFxKTdhhw3N3lZsMCGsZPsJTXZgEJZ3SOkq09Hekao+suMkwdFOCuumEiAx
adpVhsrDRg4Zsw/eya95iuOUGTmI1N0+IdTu9BW0cuuU3OmeM2hfICkrfmO7/1ezsYO98PHeiVru
btLfPsHScL53nDSB9L7fVnX/usOGnIIj73gueXfkibYUsvRuC3cUiXSPOrWSMKkRCwBjJjhrmz8M
luAZdZkaJ992X8G6d3YzjOq0kCqwDebi2CQy6Tn2EP0ngmSweQ0oWvFyjLd4OI3dKfxRhKFX+Dlt
5emNl80r98I78NJ5IGLc/yj+QirYUNJbhfHWkW+aEcvZLYFi4kwO19KSS2KgwyWV/dHBUrv2zPEX
ysKmNvsdcnMLlUCyIwvaEUUfET4iKcu05YkmFZn3QKhjFyK1ZYyWuBKE3l/+bf+stlkqKzHroB3u
YJMARGHqci8Kw+o1kJLJYaLy/1TehLl6BXufpJ8qZLYgxoT7ebsDCbHWtB31D2JMCTjw1ZNl0egc
HYFx1ewPNay+9swIUFK7EoJW2g==
`pragma protect end_protected
