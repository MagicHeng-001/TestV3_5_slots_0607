��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��CN�M��rY���k�d��%�����]1�d	a?���u�P�e�q{�;&nĲR�OL�D��M��:O!����߸���:�6���R���{=I�9`�DW��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�I��U��RT�k�ҡ�ˊ�\ׇ]`��:�VF�'ު�ƿ�-���%&`�����Sz��g̟@
7��=�>���Ɣ���P��U1�ȯ�b��/;d��?�`���:@[��2)<�R��E��/"g�[3�\�Hp��Ml�~>�,�j�c�u�'T�0�M${�*hQ���KZɿ`F�l�7�jX�|Z�m�9��N�����9�pYKRD�5�]ĭ���g>�0� ���(b�űt�X�uƎ����c�Uҏ� �Hv7V�KZ	�|��4��q��S��[(���Ͷ�t�&�3س�����\��
#�J���:��4sſhd��2y��	܉
��p�d�a���*�~��9���Ms�*�b��A����3���R��B��i`S��sQv:<c����Ƥ���7	^���]��/&Bp+f�m5VŃ�⤼�,�ќ9=���/�=� 8ڷ=>q�1�'r��\Z7�U�c�[~��Yy�i�H�]����n��]~�O`:��u�e�co1��؂��ɮ��Ԥ�#Cro���y�d��".���n�<�t!��wȺ�C<5@xo�����S�E-�<I��9�c[�&�`73�L�p�I���T9��:$�TtL%0.z1S��P��%Me\�ϩ1S�^E.q�<>K�a�Ұl��A8�?�DD��+����s�o{h���WuXՂ$�|
��K[���Jx�%޸��A�S�ꦃ5h	���� ���� q�����UK �C�S�ǌ<|�V�)DU*f�ݖ/}�Y�����d��*_�c��{6�0��;�@/�8Cʝ��?���?���B1�M���6N�ֺ����y}nB�K-��H�js@�'�F<p ��(n�vw���Du�#�{K=ͻ+	8H��㈈��`j�]QZn�A\@/���Fe���f��Պ&��o!9��CJku���Y��Y62�J�`d?�@�0d ��?��(��l��.��aW�RTw&1�D=�m��N�����zơ����;8Fs �)� �@4�)�>�b�tz��h��M�f��W�v7�z�8�#�H~�k�S��E�y�JKoح3A���쎽��H/����L�\n��T!]-�^v�	OcT�I�T�U%�l���r�#w�����p���tϒ��p�ڃ&%~$MM#bw��|,z�Sn�/.Z.8�*��m\�m>׼�8F�s��W�{̓c8��o�?JL��5�(I#��)9��d}�1u>�ܧu��N�a�=�Zý���6����V��4�T�f`�"���p������n:h�����9��4�HVq}T��T�������V���)FbLg\-8aǛr�6��{Ad8���jP�Ꮭ`W��W7=���7�\�{W��f�'Z�;�y����J�!y,�U	���1��Mx���s�����\>p��Dx�Т��R��<���:힞��Ƚ������@U�[���߶[+�!u���Q�币����\<�h_mZV�g�����vYC(u�1�H�W��z�dy5��Sm`)�(���6�p�6�^��Ħ��:"ԬW����Ej�*�n�EA&#��?��Smpo��mc�f)�5�Y�W8����h��JD����i��'+��f�V_F6�s���cQ�}�6��	0c��-�]I+���tI�����r�jȝpNU�(�g�l����{���r�P�����}-�+g �ɡ���I*uӛF�{�D���������,�=�2�-��H��i&��5o�זH'��8��	�E
����$%�`(�xz����D��C��F�S���ů��L��K������
ηo�����SE���%����>#IwV��M>��b˵t�i^�ͷs¸AM���K/��չQ{CZ�m'l_�٦a��Z��}�9b٤�Ȭ�w�f�΀��3鱇tAv�0
���~��7�i���_��Q�_��V4#؞��i�AC���qR��ކ�������I>��!�G�S�Ա_R���OK�\o$��E:���V�~M��W}�0䙆�(GQ�}3�]*T�:�k���o.������dS��Je��g���3 �	�P����6d�%n�+���!U�/���I��Z<>y����ZEܓ����L#���J�����FR{��,�����8Eޢ� ���|:u��G�Fy��ZT{�^1�K�v�lKp�b��'Ijˊ�&��$1�
�hg\��oN����;>L@)V�%��D�3�y~A��2>��{?%:jE#�97��Иv�!G��
��`�$֋�,�X�w�\С�[;�Õ��m��/O"Z�.jB��3rh5�>����[��g�$)��j�����7���e�lKg�/���2O�6~�Zi%o^�:���2��`�%�aY���k$!P��kR�}E�l<��Π��R8h��u!��%�&���,��В�\X#�����nϕ����;�3Im�K�t
�z�df�L1�L!�'zd�Ol4����^F����Unw����h�k���o��B��-�0�ʅ�]�ɧ��ܙR�#
:�Ev�Leh��H�:�����7X*N7�P޻�\�om{a�������Ǆ��"��t�p����������0�9YN]���C����ܗ'}c�W�0�Ê�x�CB�Q��*05�<�����<f��*�2�9�<�e|�>���l���G��S�1�5��#��u�49 �e��!�����E�I��ď�����i��v.�w%P��\��t���Mp@���gv�7b=��|���RC�=	ar�Au 
ubN.�����i#酖_�"�hCo�E�'��ZV�=���tr#�����M6S-F~D����^5z3��b�6)1��Č��&)�i��x)
j�O�(�o��z}��|�[��Oh�v�j�J�hS���X'��:}�{�Q�����W��rX�3��+�c�l���?SxIR������hԔR�Z����U�xֳ=�$P+}�����_O���#�В&�˺�2����)���s@k�l~Z��5&'���c��z��F�X�Ŗ��q��˭�>����"�T��0͍P뷷˦K�v��D{G���w����b��Y��=�se�>4�@( m,d]gv��M/1�o�a����<S�DvB���<��P�@a�ɱ�B��>3�ҡD�8���%��}�G�Z�a��G*FD�k�Т�����~#�n���>KiND���*�o��|W��# 2YH-�2��^B����9E/U�����H�Wm���O@Q�%v:G/P�EC7�vW�+�LŬ$d'[���[�/	����4'�}$B讬���@8��߳���M����Qw�֔-������6��i#E<3.J@ɤ�-]�ҤjIɢWzM�ׂ�������01��U��V�y>��3��{ۖ�����n=�!CU��DM��s�8��D��6��o�:w_���'����p3{���5�4.��-@f�%ߴ�`u�@��������k����X��>匽�
Ǵ�w���{���J��T���S��PZ:�� G�FYu�>�yc��4R��{Bɨ1��A����l[ޛyC5F �[��i�袖�Ի��jY������UJ�Qʃ��+⯼�����J]k]:ɾC��7��A�k��F�B�[���:������@bcG����0k���
m����<Ѝ�YՐ/�7�)��ASr}�E��i�Z�;��^(�zmzeW>�z0�)-bzT�����\Qɍ��LN ��	����l�8'I�f���;���""(����mM��ڸ_����a����*�y�d���!y��Jq?)j��$i�J
Y��`m�4��{�����i^�j��i�z�7I���vm*��Dg3jO,�p]�U�	����4��d��-E <����a����(G)��	��Bqg�^߻T�|��#XAi{gJF�@.��Q,dP������)mR%9`� �@qwL���D�c9 ��
��"&��P�[��8.�?/	?��ap+��+6�Ĉ�a�Θ��(+j;��O�W�Bά�=_Z��,."��4!��#�S�u��|�o��h	�E���4��]g�az���o!7��Ԑ�y{A~���*� ?:�����s���U	�i�H*�.��
7��G�S��K�+��!=��ib�䅦L��8�Z�wL�(>R� T��C���B��--��WX�
��P	��?I1��v��ԏ�EG$Vh݋��]�VxR���d���y�
��bI�q Z�ڄ߽^$L�_��s*��$�,��خ�����G�|��/�����֕
��m[Y3 ��^|�tD�.���Q���TO�>*�Ճ�RF�ջ�Pz�Q"���`��	(�A3+հ�_#HYS�z����FXU-v��9G.�%��WU��	��r��~�}eT/T�ViP��40�q�j`�yP����@7{��hJ<�X���pb}�<���ǿ����O�
V	�{��ܰL�DP�>�G���]���6��=5��<(��0��3~�o	U$����ug�!U!���	��)��y�P<�Rmi���\�0ޗ)��76_�**� Q��=a���Dɭl��(� �s~��W��f��9���|Ujݔ߽of���ǉ�������{4MK"�S�C����G��*����n�L݈��G��~}$��Ԗ8�/�����"#u�6�^�܁�;ZD�2����X �����oA!�ys�Q ����Hq�4b-�_M:i�y�߬4�DNt=�P�E7^��\������*Η�n���vy˝d��r�#Ð?sX��P¨8�5����� w�}��/՝�������0���V�d�鶇f��&5����#�\�X�����=��f�κ��<�i���{Pa�X�ھ61K��sqY��ި�#(�XNM��-�Js\�Vߌ�^ 5|9��L���`W�fOھ�
ЪʹI�h�QGv�G�m���\�L5�G�����܉M�"���y��Qц�>>gu3Hs�-7��+��~�5�Ň�1�'6듰��(��^!$�K	K��m�QH�n��G_e�L�74X�=@U�vN?*:�G�ƽ�Ɣ3���J�q.���F�����-�2u�,ڕM��:���s
j�a����5ȿ��h���{�\;[3�笃h�~��}�Y����HN7�A�?�u�A��W4r$^���=��A����W�Gڞ3h}iT,ѭ��^#�;)�m�6R�y���Pf���v�r���Q	��2�/u�IrB;Uo2�gNTо|�j"^Sn\o�). ���`g�.����7�Y?f�\7�=�&H\Q,I���ȧ������@����D̢)���9�ts�xt���G���^Kb��`�ʷĿ�A��Aa� �񓡪1���˷�{�pY��yj�X0!(S��#��F��aug ��d�X]���毈�q���2WFa�%���$��{��F��9�V�s&+zב�}�WB��R�Շ��֚6{1�ĤQ,�tSr��'�cן"wŔ	7b��wF��M%�W��h�-�F��zc�'oTX#���Ɖ��f�&�T��v�o�#:��{��q������$x���ۜ�\���+��o�b�q�W�M�Z��+i*u��~$�1�S)7+�������.�M�ہ�����8�C~Y�~���!��s�͗��|����ߒ��W����t*�A�X�bpٓ]?T��ZԔ��3OQ�	�&�'�
�0�����?Si1a��D��C\&&���j�-�^�glD�0�B��(҂���8����xV)�(��{ 5���#E����G��ҏ�z;	�:��]�D�p}%Y���"��*j���#�T:8�x��,P;��钉�'����"�R�����6╹4�BW�zO�f�)��� �^1<	F�S�׬�Q`
R֯�K�q�P�osfd��r/�T��`?��U�|�(S�삅5P�mVo�7��57բ��rI5@��n_�"�XGɀ䤻e��^�&���)��굻�c�W;%!�dT�U��
��r:<�]ɰ/�x��Ƀ�j�1q���I�.�ܿ6#�);kC�J�d�fPL��rc���ǟ��H�`u�I�8"o����b��gz�y.�R��ڙқ� ]�n�u�YD_'���P6�F�m��jwG{4�鐢>3��dVӝ�0
H�~��F�cIo�}�}�,��\\Gɮ��/�>�-�i���lL����o�uʛS����pu������x^��\�>�pIk]��15XW����qXp�O]�Kh�SQ��(������B��D�Q��V'��~ʄ�b�l]��1!$��0��"�E!�/ HPk�K�(���r��ɪ|�@ �{'Gbg2�cT�9 .V��	^-�V��������懋R�JB�6uMYE���nI����M���T����;��3��*�6_9��^���riK8�l�t� <f�՟{��{B�k���7ͪ��e�~��c��R����(��>ٖ���?�m�>=�dÉvrXj�)��I�wU���bø�]�ӀpH���O)ߴ�K�����	tP)�ۤ2�B�ɪ)l.�����%8��_@r�. ��y�{�`L�����v|�]hT����$v���S��^�z1�X>�F��j�������0)�"��r�*᱋�NL �ړ�:IXY��Sq�g=}2�ɪ~�iS�D�9@4:��CLnȪ$GD��^����Е�V���I'�o�O
��������V��y��5��yC�[
t#x���D�5���=ųdu��*�	��Ҝ�g~4VZ)�K�er�R]�A;(����� �_�n6A	pqj釥�bW���
��"�ߥ��	)`Q��%��L
�(48��������hIe%�V��T�c1cY��!���MU[�0>�K���6��0��)B�gK �D{��$���`aƿ��#��+b��5��5�F��(̟�:	�DG}ʣ��[�V��~qlr3����]�`{>!¡d����Em�'������W����=#�ڲ}��'���oJeNO�C�L�g��W"��|V��m�uN�iäk��GbT��aA�Q�h������ |�!���yG��M�gb�T�^�v�C��F�u����&�K\gEU���'����LtL�Z��L��\�s�"wC�|�;fl�b(D!a��:�Aik ������)�cz���Z����Q�mQ=f�\���%M��J��[�y4�䖼u?mfƁk��>X��(��,�ዑ����R���`�Y3Jr�c�04|O�䴃��Ȏ�@���������ec��F-\*� �u�����sd��l��s����8�R�=�1�3KNMV}�7x��)֊�}24W0����'�k�SM�v&Y@� hY44x#�Ȟ�O��&�����ƚ��B��D��Do�XZ"��UT��fD{҅�٬$*�-yÉ����M���|���CY�Ɇ���͈�؉L����ࠉe�)�du�'Z��kD�ƺ݆gKB,�@kq�ek��M�u��'J��8y��%���p?�-vH��)��{Ss� $�K��M�,x��IcA]-�at"|,�`�w�{��Au̧�y���,\�W��+���>�N�?�n��U�շu��0ﻉ h#'%��L�b� ���Ot#\�'d�ʴ��j0#d|k�%'B�+P�R��
��6ם^p� ���.V�8���z2��~�/��6�>blǦ���D{W{���d�6��%�SS8f����	��DG��L(��'5��ʭ�+�I�c�Y)�E�e�ɒR�5�"Rxė�w#�WJ���B�� O��E�� ��
ī2���}��HS[�ߢ��֩��p���2��.}�`��a������-� 
��x��d���}�G=D ҈Z��At���g-��_r��Y1r�-�9a�|��,�\�¿���~�Qe�8�̰jz��N��b��{*���[CY���[���Ii�pAbH\IH�3���D��b�7K��v�W6k��_�g�y��4n5�H��x��f�+�����<�G���ۃ�_���.�dh$a�솯��Ii����^�+=��G���8|:�ƛ���++�(�i���Z�k����cEN�����2�4�u-n�ƕ�6��n��Z�������oVJ0��fk���!�۠t~~S���������E�$
`;Y8y]E��G�z�l1tU/�����S����`*�h@yJ��.?y�s�=jlv︮7���}.E��D���:V�����Oo���1��R���^��ӿI�������o�X~Emr*]Y�fP<��D�j%ߘ�V�ةh�,=ݝP�ÿ���9&�8/�K�k6(�"�»ұ�*���p�M}޽�]0�N��Es�]�U���D�BOe4d5�`��|g�$Y:��Ws�)�& ��5��ڳ���Y_�\_���X�T�h_y��Q2��dSE��XY?����B}�*��r�?	�ݏ�Q�N\nR��!�Cm9ôT�ȇ/b����$�ڡ Jk-\�(<)�R@O"������U��ܲ.���� M�r/z�'�ޔ�, ,Li��k��MLsP��P���A9�����M�vm <`��C2R]V@_`��Q1�H�l�4=E�{,��<ZA�{�<#z榯t��'T�wi�I���*�h�wb@���`�n)*d�۵�Ω}��6x�j���9sh.fD�E�nN������q�r���0��+���C&�k��}E�Ӄu�Uc%V�����S�/q�W((�Z0յ�]=n����J�����ꔔ\[�
Ҷ�t�L}�t�~m����O�3ᙞ�9��f2j��O���U�'�6;�`E��.��-��;����Q�yǽq��Y��O���&C��`�:W��(��+�=��(�N��p�:�*ޡl�eb���$��>i?���hm�����j���i˭	u~`}����j5�&���թ�<t��c ד�P����|zS��p��Ȁ����Ut���KM�N�s�̔����iZ���紦���n�X��ێ�C�S�%\r\y7�!�<lf%���N<�I���iSd
�0tIrl�LR����U���`Җ�S�ԝ�1�9\�ÖF�#~��ЩYC����$�+p`��@�&��]bS��U�$����.��B�؃x��vɄ<�V�aDE	���hk-������0�k�sΓ�❚�z����6���&�����[%j�����;��'��ˍbx)K��hr83{��5*��mc;���)j���XY;ҧ������!S*`�_3�QeEW��F�ۦ�꫉:�w�.n9��:O�H� ���UvĘ`7gl>�O'1Ľ����= ��Mm�	&F�������O��'����թ���TPn���T�oO�V�����R���l�?������_�u��¤�҂6ʘU7{�T�'Q������N2^����NN/��������B��a�.�7�c�'��1B�0��"f�^Z�Γ ���[�?y0�4�i#�'Df�Z����9�+w`���/���=E�}�@�������G�Q9ߪ.�J�zs�̃���!�0G?@�p!�x�^d����tk��g��hc�����a�?�(T��.����t�֑3�&u/�s
�v�$;�W���d3�(����Rm��.��{ⲇ1~�0��	��Es� a+*�� $��<���������v p�q�̃�l�$"�y��}�6���O5|�(ߙ�h��x��vFaP����s*w*�zvH��&|5]�HC�5-�+A�TG�ӥ��gF}�^����oo�Rd�(d˂u�^�ع��aX�	�� �= `�KK7Q��xj�_"Ս�B��(�j�����킶����a�K#�b[�8�Q-��
8�C��lx굙��+g(T<͸�ԗٝ0��5XGz�Q@�@J�Tbȡ.C��}����A�Ѽ�A�r�(+l~y�Ti�"�p��������:�k���o��Pj/�&%��h$�o�/�}���˱�����6���j��PZo�=�#�r��fQ���=IB��L�W	�;���{����L�e���"K��\ޭX�H��KJ�EU���G��xN��.)G�? �sC�쑇bOΏ'�*�Ɓ��^t�g@MG���ݨ�������T�l26U)�+R�td�E��?5j�}ŏT(���v�q�ډ�D@�GM��al��"���m��G�\C�좨=��~��epq� �	�H/L7O*"'_T�	:E�@�:f�L�ba� ,�Zݦh6V�I7GMk�M@fZ?�3*[*�Z���k�!�3Eě`>����?8��*��G*El�;t�����v='�'[ur���茠�/u�;c6߿�<0�[���`��@�{�A4!��󰞷��@���ui*���s�,��(͖��mV!SX�(yl��<T�%�c�̬�sgoɑ$���K� p)�w�x8�6�x��l���/N{�@�Q�eU�[�"Uc�g�������9F��X	N1������p/�b����� nVD��\��:�|�R�6ޔ�	͓��t	�cfv Uyb"��:�vw�{�g��?����ѱ�a��v�(Ox��o.���¨�ab�D�p�s\��]�\�y�) MW�����������,u��/�
P�p�f�7_iN:��R9H��W�>C�6�=�PR�a�Q�$�!�J�d�nz�~��ݵ�?�,���[%tM���$�M�)v�u�3=e���g\�������: a�Z;�p�,+ҍޙɄ�1�dA]J��q[-ͮ��k8{)���;e@-%��X�2� �v���i�MTz�DW������Bķ!	xF���/���'nQk@�K����=�5�h{�X<)�LS������5�+o�"Sc�����������WK��w�F9�c�%�w52GoY��v��UI,"�x2�V���-�Lj�&8�m�&�@f�� =+�?%!��!�h��X���0$«񢻅�h���NJZ���A�o��2W�ay;�$�(�=�/}Ĵ�pߙ����K��l匚,���E8���2�����-��&�H1x�E�D&�_�6����\;\����Yr[��gR�#�9gEj���ZU7��1Ѹ{�k'f0�b��=�!�Ӳfx�^YX�M"�-��N(L��,|��ṵ=ƗLS�Z�>p���4�R��4��N����1�{Q��f
��̢�r�e7
�jU��PX�w5��W�oe��*6-�dH������B�y֋ɯ+�W3�ZPv�m��[<M,I��@^I���n��#B��J����q3���`�A��y��j7n�*�$�4 b��jY�O��0;�}�)À�bU��I�����8؄�-b���l�ˊR�� qlw���kH�ky�v��H��)Y�W	q�Bҽ]��
�eD�NAFS�2r��.�ũN�����<z\���p#�m3��j�բ5�Z�x�\���?�{�Y�T��z�3	�X~�9�a�#�[���S:�S�Yb6��'��꿃N�'Х��UX⹖bhA���n��=������dK�ꓻbRf�a�ʓ:����7(�ײ%���3�v<�c`ÈG׾w�d�xq�^"P�@QX���:�W(%��������3J��57��� �R>4�6\ź�IрA�ު%��}�Q�ڂf��?O���n��;�ʾ`K�0%e������(';9���CDg�( B �W����#��}+)��϶y�"wjQ���_��BN��P��f�E%��������V����Ff	_�~FR>������ו���"M���EO��(h��2��Q_���ڴ� �s�AzM�)�TX�:�۴��Z<e�X�@W:�M�O1�#�]��3E9�AeX��rM�rT����S~O�ͳ�d���x��
�C���$�8�#eyl�#���LDh�����-%q�H��/��iz���Y����a>Y��*�.��I�i^���J�K���U��T��R��Rt
hQ����C����v<UUB�Si���#^��n���Wɱ�mʖ�59�S�Qk"qr��V�\RY�z��.��!˟vI?�xx�ԗ�*2�)Ѯ� �"߿�A�+�_�3R��Lgf����iyG��\~���9q)7�
{��<���jJ�ےsݨ���>I��pkc��ٗj� ��l�Mgs�.8��O�E�l�s��7U!��({�iO'{N�f��(a�m��"�o��Y~I=r��4
;�&ͥ.�v��������l��įg���$?��E���I�/2��$a��B�RL��

\�]^ ��e�i{[~���sblV���oe�Q��6�� ��u���?�ФIh���0�s��[��-���&�Y��/s|VU���MFt![�+���]՘/%Zk%�p>6a�5�3�O,}���t�.QQ��*J����M�t4;NC}�U��8R?����(��r��	����P���l����_�Gf~!.��ɝ�Y��OA�����;y��3��s`�"�0⣛�}��J�;B��)���X�1!޷"1Sp�j�O��	:7�����Ui�٦�e�X���ϬKF݆�x+%V��_[�L!�%d���g�'e�u{����O#>^=ec�\���;Src�5�d�J���d�-��	Sy� 4e��a�C��I?�rWc͝� 5�����"����εPF��*�ȇ��v������ciQ(�p�����:$����z':�hJ`���F��s��w��i�O�	, 5�b�9>���W��b;������?��Z�5q���,1����Q0H��?�){�K�bJ˭[;����I��&�d:�(0MM�"�����j>�}����p�%�[��9�E��+q��V�ᙏ3i6��,������_��a^�"�e���s�Y����x������-���x-����ٞH*��drj�n�����(�Y���D=�H�kEpc��ɛ�t�|����~HUSm��=���(�N��t�g�7Z=!��SǨ��a,D��g7������N�ZG�n"�I�ϴ�NBP��(�Y�&�=�?����3��y��z���ܘ���&�Ŷ ����`j5 C�y�J�x�nW��e�9%}�� �xhfg�Ɔ�@;��nZ��G�+��K7¬O��b���FJ�21I`�'�~�m�K|��좑0w�4�N[��b6��(�7��-����8u���/�g��y�E9p��P���i74���q�dC���o�3.PoAT�������Kg %���(0$:���?��h�`V��c�ެ,ff3{"��|$>%����Gc���}@���ͅ
��
�8��ּ,>�0R���h�w3�5v�# �Ys�4��W��3�T2bŏzr�Y��3��h}�^���7��\�*$bdsw�^�}���#�����lJ���ª�.�-W%�=֨?�i�bNb�}���i��Q=[�F}��P;�<���8�7JBRn��/�+��1M���y~���5[�f��������$�3�~=4���c�#�F��78�U���w�^[�޺�c^P�leM�j����R����~:3��=u9��,���K���8HxLLqL����Ę����J�a�
1����c�q�����Ƌ��>�?���=��%9�sw�YR�)C~R���$v�El|݄{Z���������(���)���f�%2V�hT��ʖ�4T�B�%ޫ��cz��&�X=���WW����N��;�лo����}LYt���ϹNhR��t6�g�e�b�����a V�xO�6�>j����YT�zW۫��$��@T��ٰ]�򺦳��I_��A�<{���V�`��Hx+�s5A���>#k\>���m�r��Pމش���1���JL
�ak/�#��ǘ����&i> ����y >tA,�h��X�=$q/���6�ى�Ё���x~Vg��9���H����7�����O�)`&V�)�{�\��[I��y�ͅ�n0eӂ���\�m�5��~�UK��}j�f-���C7CsFy�0�'_��	�Ŋ/���|Q�8@�!�Z�IF)̃y��`)>sۢ�q'��Z|�������`��(󃻮5>fZ=����X�`�s��-��{6 KB���ky�;����oN�?�����sɋ�B�c쒣�N8�P�F)�S]��O����jr5���=�W�o������f;a��|�Y��N��԰UIf"�Ak}ۅ\[B��Z�q���?��=�R���µ���4χ�k��#f���`�_r����I�8k��oO��u���O��-�&^�xx��6�	�B�d�Дo��:��0��4�!M����Y���K����P�p:x��?�4��ʁ�z9O��y�4�Ѫ(�?� f��;|l����dƗ���F,S��
�-�	���r �#x�ԧ �g����G_� ������c���*s�@q"���� v���M9�%
��c�Y�?��̖*�G!�mj���˜�e$3���Z�L:u���_BW� �k���ɯ��a/��׭LoF�J��9�:4 �ֈ���!�S�]T�TbV�P$R%;ߢ�O^��}��@�d�S���]�_��p;�������>�\ �<�AS]�N��g�<B�_R�@����e����N��N�&�6�Bob��0]B����ynY���,t�[�Z�\`A�ڊ�b�g�}�B~"״��p��1A�ڈ&'�?�i�'�j4:�����*`�� <��7p$ ��P0C�?J1K��S�S=]��<���,�n�=�d��>�1���o�)t��=��]j]4U���e��^nC�U<V}�υ���ym��d�7ʦ�`�'l��'���B�/%����qd����I�D��E�'27��~�e%H�r�k��?bDi�ǈ>_�'e;�(yM�҇�T�ؤ�`Ħ�R[֒�R0.>{��M��s3a1i����� ��-1ę7rs)��qP��	G��+��6&P�7NlX��[�$���|����Z��E�-��I�J�Ҹ;�����En	�؇�9i����p$�JsP.� ¤K�5	�"�§���A,�H�A�C	��S��94�r��#�9N�T�"f$t�d��z��f��Fv�}�ٰRG�]��~n�Y�t3��DL �6�����v��昀��|l�L�*Ca*���?�v��?��+v��x �[�{q�(�D��pO~���tI�h`x��t��c��/.���-��.��a������
�ܚ�Zr
.l6Za�wi����y����_D�.�򎔔�ڪu�|0��*%Do��ݓ��y;"�������;!%o�2W�]��I�LV
>g&En��g���Ј����
x�Հ��x;�UФ� ����=�����PB�r���)%�"��܏��j��I��E;���� R�n���И�*��Y���!U"������7~[q����{���3ݬr/b� �t����($j�F���`׌��nqyT�@ ���%���P�$�%WS���IO�-n c��^��e�Jئh���L$W��߹����� �Im��"@V� ��>���=<It�{��/sB(��ǬO�U�`�"-�a?Cſ��44�R\x��<]��t��B��ݳL������e�5Pm9U�?���[<K7�l�A�D���
	��xTued�#�$�P{I�����K�)�a�й�zU�ژ��]z���_�<:�c2�t+�!&㗵���<��̊������p7+�vw$��b��9tR��h�Y\�ë���!���@�V�m�2��% ��}݇�B�PM���0�)�S�YU���T�ܤ\CJ�k��S�)��z
{���k4(��8�����Ú��y[����/�������G1𤤀����z t@;Ѣj{��e.���f�A�ǟ8�zs18�������v3� ���C���c����`�MR"Pi�K�f!��U3��&�\�/�;��0�1�'kufPa���D[EA"�~���~����&�+�~�U���H�*����n�9!�8���K��Q��di �E�����'�OQ���g v0=��f�?cK8�&���8~��+�A�}��l�*.*n���W�Rk�-t�O�K}ՠ����p���;��I���e���O�jj����D��VK·���-"�ظU�H+zH�8����n�I�q(*��W��~%;�� �
�Q&�S2�!{X'*�y3��0�s�Ε��cAL��P`&N�0���q2��e��'��ʆ3v�ؠ����BR��� ���oƫ�	��Z�U`;����N�w��#�D��-�[����H�J����G�g2���C1�#&7뙡��!>o9��Sզng,��su�p�Q[�R)b��+��3~G̪�}��8ǝ�3]^K���S�Rsao�񖝬*W��sC�\_Rg��er�vh\�W�Jz/$�te�?�"��M���sC�<M~�$��l�3�)$`07�]P>�R���䌌V59����"�̓
�kx6U��Q"���&j�E�/��3�5�h�˕Pt�oJ��x]~���6�p�<�ծˉ������~4Z*U��(=5v����Ǜ�t��Y2MۃD���U��k�mN��@mTV�̔R�ͥ5O'��𚷟�D��PλU����FC�	�M��1�F.d�֠��048��)"%w����M��4�b)��z�!,�"E�ҽ���vh�Ҭ8����p�,�\	�J�t�
�B�y�����8�&F�`F_�xE�R��5��I{�/����TYJ� p��;�_��PB�A��bd89���(Z��k�7���4v*�&ZݖP��#��MzL��Ҿ�����Q*m8)�U���ĈL=}��S�5%m��a��c
�4л�{�.>���1C��!J���A'���}%� 	��`�#���}��5�0�9��0W���Z4OpjB�ۍ@G�2P2f�c>�|�v�q�����<4�fv��٣�aiۗ-��4�c%Qv��~Z�� ���S�9���3]XNT����Sqi�`MVp��7��tñ�}Y��ڣ�س��F^D� ��y���i^b�^�°�^�O%�Pc���׼��|A�D�Ts��uYqN��B�FrSɅ�A��hR���>��tzİ�ac�����(�a�GD�������Y���S�]�b��R�5R���9rc��)�Bo�U(@iǓ��3�dG� �DWn��Y��)��a��x��"�pA���u�9(,Ik���E���3���0{#���id�'e��E���0���1�?�F5��^�S��];�~+3���o,�h���	l[c���9�o�D�kۇ�\�A޾e�fF��3���tyM� GmՃ�w��4�Ur=�:^�<)�X��M}�2�൘�`�`-�Y�V����e3�M�l��nmv*}�+�f儔*���W��EJ�a����W5�"FN�Z6&�`Ԗ�w�����]��@o��,� ���	�e���\]W��5�l������n�՛���{�Jy���h��W:�6r��� ��zs�-��F(������1U�l��}8 �..G*���&���~�:��N�}MǬ9R�IV�^tp(��ō��r��P��a�=��ӵ=4����$��H��(��J ���n���H��i�ޓ������5�MǦ�ܫ�=^T��(%K�ك0�T��R뾚o�~u�g�N`�l<uc]��S۔����=��%hg@q� ��n;0�L�X3@lH�.�����6{��qC�r�~����9|�g�c�M]ByUg[窹U��������yvs!U�G9�dٸsg��cPP�����>��F� ��s�����A[�_,'SU��I�^$��l���LS�6��|ʊ�Ű���MV`�ǵퟸ[U_I�[w��ȷH�t��Tc�W�H���WD����ߺ"���(�QzD�-K}`^��⋅������"c�-��)�鱨�W��~��b-ë=.H�^u� �r����Ȇj�	�k����F�0tj��n�J��{K
y�)�= �c���Oc���e-k���[
��m%d��u9��"�
q�k��� I����"W�	��e�)�떚~"��Mُ���u�W��p�z�b�S��f���fͮ���p��NdH�'N������q�t_0�*�:��k$�GZ��Q8K��	Ę�x7�� �b�;��V����,�oMz�V��ep��!��Ƚa��y��2v9�ڍ�(I��e�܈�ݙĝ����P!*谛A�yƚɛ�X8>�t�!�:u�s�ZP�0WQjT���T�۽b{���
H$�ct_�;�ӤYz�z�j�OL3m]@��L�[��Č�{T�E�[U�ɖ3/e�;7����X���p"�
�$���y����M��xUk�7\Ӱj�U�x`�Y_B*z��KxX�$"d
��F�d/fÀ�a|����"�5�W(�fVS���^-�e02z��z���k��65G{�f5g������G
���"W�X��1D8��9m�X��X����g�W�T�m���!�NJ�����IM���4�ؑ���0���v>ܰ;gyDw⌆��Vi��`������>Y���k��.+�O�r^�J���X�ιR�)�̼7��%�|+��}���
�&گu��.Hܢ�E$G崖����M&j�J��jd�����85�U��c��$P���+�h/'�>_�/��g� ��mu����u@��n��Z�(b�ȹ���""�6�nj2@��4�tW�	�A״��� ��9��'�Ħbu��+ԝ�ig�7��(�+dt�p�}2�y�S��\$���z�K��� Sl�B88F<m�	�X�F�`8�)FE:� U�ߞ�\��e[���}�|�j�Eݩ*`�㏂ɶ�>�gB}���kO�~�N��*h���S�ЪFCeZ��4P����2\�@l=�ݭ�꒹�,'������ZE6����ߚ!
&��5_����������y)EL��'��,o���t��٨�͵�������Ճ����˕��o�.T��N������T{�Ez�E�U� ��:�&���S�b�{�~�kz�b!C*�C�)Un�]|��J?"n���K������6N����Γ�W)($H3�p��d�׋߀��$L�Й�����u�<l1�5(�����U�,�c#t�����ĸ�qJ��Tp��J�]z`�R%ub>�Ĺϐy8Ӕ1C�U��zk�)c�PJ�ʾ�u�I~ ��	���1�aS��l�9�f��Њ�M�̠G�X�?�N���	��Q$xxj��ǘ���H ��S
� ��>C���3!^j�?3w���V��(CI7��Ş2��%A��T�D�pz��9�.4Cӣ�r*O�����fܙa���rrZ����������D6�w�cdF�&�Ć��iEc׊{F\�����;�dD�oI�F��=s^�<���[n;"S�w�ɐ-���.��&��'N��g7�7fV���l�W��*�9�G{�*��c��[�r�s�X�#� }��k�)�ݖ}Q�%$Y'q�dW1B�W��T�-R�J4�0��?� ����R��z��SS���E!���cJ��fd��r�B�{;�s�r�v��Mܬ/,��`	�*��(�|C��ӗ0a���HB`�f��H��~����	q^+95t�I��:VE5��@���wK�"�0��q9\��9������`9hl#�;ג�P|��0z���NsvXM+��C��(b�ͬT�i�|A,kq�P!}Q���Dk��V*�ߡ�`�W��ĩ�p�S!}U�dgЂɭ�QS{�Zh郺ݞ;��05�Oњ��[�ا��N&O3�v�\��DT7-��1�o.o"���&5+!�� g<�|�,PV���tS]ſ���<5�Bm����O�ы=h]��+.��
0�g���	�����p�Ҫ��`�s�O���ֽq�F�G0�9x*�P�.;9�A[_"�8w(��W���9t���LxH���}��yW�IM����'UY�|�ƠE3�|���n
���m��R5��Z"Ti!�hY���D�����6\X%��N�����=w�P����k�yR؍������b�p,d���,�ݩR�vq�qp�es}I��1�m�	Vg��=�Fo�w;�WQW�n�9�!E#9L)1mb��I�q�;*�+�e�Yc�%���3�,�P�f��װJ#���'��>����J��e��u�c?#�*&�q���� �^����`j��X����^�������w-��
O2B�1Ԍ���/�Cj��\�SCn����+��.���W��!i��yO�b?m�I�SK�V�c�&/�$w=]��8ʩ"�H��n{}�T#m��w��Q��uN�"{I������A��	]�r�;:�;zԴҰc�\�UJ�C�d:Rif��8��f��:Ť��@�TC�<t����5����<1�<�T����d� j6�g�os�"^[�>�6�:��y^�SV�t�t��� ѡ��@��N��7��i��Y�"�ي��&"�z�������ت��"��u_�&&�¢Gj����X'�d[���<������;�U�R���3�U��o�糺^�a�GEr�q;R$�f���E�2��+L$AVbr�^~#�9{Q�����_��N��;KnW�Z��e���{����}���i�X�;�q�4a^� ߺ�|\�}��/�n�����4������zy`�*���dI)Qt��\3Jܬ��o;ㆩxf}���7��4CfZ�V��Aps�m���'����*�3�[��hѰ�$�L�L��IK�I���s6���@#|��1�Fo!�p���;���oS����{���q^F.y�uR`|��5�3�#ٝ�ܗdz+�d8fSŁK8�����So�*�A!��HԴ�h��X�N�nrZ-�̵4*a��,�k�8��%�/�'�	9߁���� ���פ~��K��q����]�v��(��˺��AQ!�}5��W������������󤺼�Q?m����򿲍Vu��E��.u���B7"<�ٮ2h��9*l<��X�7G�~���D{�͖�{о\�5i8�A�%D���.UR�Fn��[��͟y-��u�$�8F � �M�a����.�|��n��{m�U�8$%�,C�^�1�-Ѥ	�f�	}�-�"A��JĸC�q	�m��<��x @غ�aUp�Tڞzh�A�Y-�׽��o�;Zw�-n����-�ř\����4��WO[����Ԑ_����3�{���U��~|�j<c�@�bЉ{$q�\�>/pRY� @i;LVV���_j9��H�ow�4u�����`rw�ö�x�1��E�����)B�y"ћRt�#��7N"�\�J��*�g��>r'��c�vp�:��r�9��g7��C�Z��+�E�\Ø��|�'�m_��@��H��h��$�+q�I ��!���M����j�V���u1x]��E�� ~4b��Jr����=|���;߆+캾Y�OS�"˶��t����?���9����syPl򮫲�k�LN���@����e�b��J�&#��OL�5����K6�RR��>����	*�����g՘��I�.�j"�wJ���.��QAGi5"�N���W�cg��X$����D�}���ō�$ϓ��-�B�*�`����n:h��E�i�ɼ�~c�/]l�ߡg'�q�lJa���# �$#Caf���8�X��)�&�^C�X��ÒT��q�ɑ�.+����ukr�"~��=�si����j���p��=�����P]1�v8��a'g:�jͯ�ԝK6�#ɠ���A��e��/V�9*��L�9�"�z�]k&�2nA��@�e:]��c�P��gv����n�!��G�E������+�x{�G��� S�J�+����5�������S<�/�~c�H�-�X:��V\	��eқ�R��ƍ~���
��6���[�n�o>b�]���
�KW���9"?;Z�o�}H�>oo�F?�ŋ�'��K��۹.�%��5���N>����m�X��^��EY(�� Ҋ��z����pv��.��\�>ڃ�����zU��Z���M4����!�9\�*d�|�H�D��3�F ہJ,ִ���nx��ehg�A��"�-�Ҁ=w��r���'�l�'9�^��T���Ǣ$_`vJ!.�z��F��������>
~WnN�Л�;�v�t ��Cq�^\A�9�gZ,�w���_��O2솜�3f��(k��+�^�tV���Yq7��V�^P*^U��5���V���1�.e5�e�$���/�f+�Q]g�B/��wB�У�R�^�%	
���^���B�g�>�Gl��������{qX�40|V
���!�cθ-�m�]2|}��l�go�vc�E.�I�ré����?�JԞk��%.��ޔ�Y�#��bm����pO�����3�eК~���=o�������~��WL��%��!4[ �{��C�ɤ���B��Q���~�`Ҵ�IVpnȊA�j������h��6�17�A�j�Z�� ϻ��M�(|�/V7��%�HH�׾w�wW^���"����.Q�lӻ�/��C���8?[I{�&��j���z���m<�z����g	�K�J�������
.{��� T��-�r�dvm�@� ���j<���?�^�I���D[��C0�'���=�ԶP���j�8�Om����D�<|�������	�:�6D����A��2|ā�:��Y���=�Q1�4�����=nx��倧6	p"9'�B�(�h�������[�k�E�"�u�j���ni'�-�E�Cr�EQJ�'��:�m�||�mMjv�-�o>�NmՁ53�� �t5���a��M��UEnwq�4r�ِ<�G����Ӗ�s6F`0ǁˁ;_�R ������R�zJ
!����_&�N9R���(�R�B0��������Tj6��g�%ey�!�7����~�2[>�-�XLtȻ2���6�D�����>����r�և>_�I��Lj,�E�s`l�-���2M��v&b�qE����AQ�ؘVѐ��ӋQV�5�و���r��;�;F&w�}d��bc����	�� ���E^SW�A��sn~�9�n�����Ը044!xy9փ��T=�h��ء(��.]��g�>�n�s��i�>��~�� ��q�;�i�Q���a��M���,3�[�΂��b��,{�-����T%��h*��>��~ok!�%����l�}]�G�]��w�� hQS�2+}�K2�w�3P
M+ZTq*�z��z�/׬^)���>̥u�6��R �)3���*����-t�Y���g��r��I���|���(�%�h$�8V ��"z,1�M���#!�+g�T��zӒ+²0ո�^�S�$���|Sn�N�VP��EX2�l��c(]�f�� ۅf����H��HKp�a(��(�ki�r�݉>B�Ni	�p�ݲME�D���n����P���@a��M�QE����琀/#�1�y-��C&joUc�)Owƣ���5I!��׿�@ʉ�B�w:b��-��*:h{w�L���x�fO!iȹ���d��H8�,��*P��6�� ��p^��a0�<Z�JP��y����|�ï�'}_e�,��!����?��vn�B��l�-ͧ��O���D�4��t�x�Ԙ&��P��g�	�b0}]e��";����l#sS�y�T�ټ��&�J'C!7oOǋ��b�2B?�D�m�+�%�k�6u�)�oq��k��֊�����a!�<�	�W����;ei
N]��i{�"m��T�Z�����"�.z�t����҆]�O]>Z[�` Ai����6c���1Aάdu~R�~V�� �G���!�����õ�1�����i��������0m��,�JPVAD˃!,��������Q�10<�m�����¨����"�hf��gt�4�I�;�c�nA@�!�z�A[��h��$�� >�5�NVn��a���S�9��24����3,�h5���rQ�pq'�s�	��8�A�t�����Gʾ�E#|^[��Nl)�(~�r�&Z[g�3l6��5�o��헄���@3��]5i���Lſ�F�2�y�|�*�q�`� �����2�չ��*�Q��|�즥�Eq�G>�L}��yKo��R���&�ɭ��k7�!�='��1W|<g��>�,��z&��JË�"�%��:������U?6��x_�95�ցR�S�8��2a��>�E h�_�Q�P����sS��͠���v����-�N��{�Kz��%h���@����c +¦
8T[^V��(�yՖ�9��psXC6�}�G;�]>*��`�r��b-${��m�N��<`R����X4�Q&�[nn��0d�'6��i� Uol��&�f�M�N"���N�Q6�EP���ϼ��n����|؍���hơC��X�}rW�.�If�z�����BDv���w����!��rǌ`LĘe, �S��-�!��ɯL�����`�T(��q���4���������`����Y�/ -1q��=���Q�LF��5� \���gݲ#)�����;�����������J/c^�*�i�E�8$�u�6���݋.�<G�d0T����V��7����Z�ǫ��6��,�2ƃh⒨N���.����z��Yt���pf}ڰn8�$����)�ma�"8`��7�KX��������%w(�?�^x4ka@p��W2�n��Ͷ��Z?8n�ŞKnzu��SP�D5�+��7�
�5O� )4�h����0r��e�|������*���w˳7`�~C�9wn��ʗ�g��^��}".��6Q�Ej�9]�6����6(c���}�'I�aS!��kvV��'�x[�
n����(��~���:%l3υ��m�J0j�B]�&��%��� (k����eA�P�i���:Ķ�@�&lX"��D&wmÊ#���Nq{���e=�u�=��y=AږB'���$��@�SnV�|ȍ��; �zd�Oo��w�X�\�f'�{{*��Y?�H�E?X�=ϔm{Lk�ɸ���{X[��C�KWq��]���!T���Q_N���>�P�$(��[#��㺧�3���3�a�Q�E�2���S�b�VdU&�'~U�q�\�w��6������;�!3X�����O�5���.���K.�*IM��5��;b%����NB�*j'/�>'ru�P#:?�0x����t:�N��j�7Q���	1R�4#c/8���9( ����a��YR�KD��E;�!�Gw�X�h����'���������I��z�Y�_\��ʖi��ބ�2��UJS��c�`�:���q���}g� o�������q."�Y	���B���K��zѶ��AOw�;)}���'�݃��ߦx��'�.�m�?��&@�
�!%[U�?Ђ��,.7^��曋4^��p5�jw��4�UĂ��� �X^DY�*��2�5�C�!S���������C��a� � �2��g��Z}��0.��g��չ�f�Er"��d�=�y:��#bc���}���?�n��9�����p�b����U9�4�I��f���́,�	��D�#v5b �-萗 8���\L�����lʻ���_�T��U�)v����	:!b�?��4��ܖ,jd�8஭��&	�()��`U0�?����h�I|�I9PDI��ϫ	�3�:��S):ń3ـC|w/�q�zD�,al�[u9�G5�ｿ��Ө������x_oݞ\��9)�F�3A?��^DI���K��2E��@H�������~���[�ٻ��.�Ѓ[��T�,x���U,M< b����%�H0�d�1���귬��G�I����Za;_;�����)�Hi�����V �%��L��띊p�����T���5�����zm\�F��"e���t�a*�5��n��+�+����;�m@�ꭻ7iI�Aj�# t>���ZČ3-��;.?�q&0�Zzj^B��L�y��x��۰��*Ȅ����r�7�0b��\���&�ަ��}"�/v�ϵ�?�w7�Bb�J�8ӗ=o?[5L	�Y��͉�M�"R���[︒��gY��.�k�p'�¼�7��q�,j�mC�I��x��R
e:�Z�~��%u߫��+qz�%6��6`h�T����^���K�(�� zBl��z�
�ez�kA�㡪H���h��n&��k��NsB�2?lk��$��MQaa���aM!�� WN������E����/�����猀P|��Q������~W|��C����0!�!�K����ލ��U�|�(,���ީ�:)8P���g���̉���*�D�"�q�?m�5��� �Cʴ�=�uI�%R��'�NZ)�<�h�Gp	7�g<H��8c#�@`w/�T����ǐ�WE�2��s��J��ۀ��2������J�|�r�,z�CJ���k��|��Q-�`ՀG~aa�̡�n�n��l�҇��XZ=Q�J4�R��Q�(���(c?%V�ov�`.Ǒ���*q2�H��]U//9d'OF�n������bN&�M��xf�I&��%���w�/��힀(=��"M�d�D`���!��
�Et������분1wqb����חn<�C7;aJ�~<�:��(�d=�	�J��:�#�OJ�0Ζ��׻]2C�h�C�B{�ܬ�*���N���&��%��9�2'w�5��I7�"3��_�f`���'~����t���/��Z)5�G1T�5�V{�0�[^7`'KI�����B�7;��?�D�	[���eHୌ�DaŜ&U�1�H[�_����7V���.�I6]wv��#�B�0nr��&(yG��de��d=R�~�F9qQ�ْ�R;x�>�MCU��KBV逷6q���Dq[�d8ᧆa�����i=�W�,"I�8x[��>�w�C/R��-4�bP� ���?Q�a�83m)e/�_����J"l�Qh�����|�c����k��`  �xa\Ћ�� @�|��1�����E,iN������ʸ��,���YTp2Y�
90��k��Z�/�D�mB��*�]������Þ~Z{�* ��r�@K�N����[���[/��?nVh���������J��t=0�lrXzk���;��h�Frq������U	N(3�	i�NbCޢ��s}<ؿ�oR��-�)��JhR-��f�� fC	��M�֍@��؄'��Z�T�ӟס���a9D<�O'n'u�j�W@ro�Ys8}/hn��w���T2��^���D�,d���ʹ�����J~�X�2�P0ǂ����_�~e�
��Ȅ̚���C�;��o�����*F��w�P����b	�u{[[<�M�L�(��/-?�2��zه�Qd�����ҍ��0s�1r�/b��?K='S������jy+��s�,��/�l2F�� ��5��Lz���5��Dk�Ҫ�2j�Mn�u`�?�U'�F����^G���ww@����5��X�����ʐw����Յ��8���Q���s�u�Ψu�z��O%G���d�V�����/K�y��"��Rb�r�?�X��S���n1B��u��8������g)p�S��z_���M�D�����ɐ#X=���8p�V e�c ��h�q�i�U7���՚���r�]D�R��Q7��^���K����h�����+pes���~
hn�F}Ȫ�
��U�2oY���(8��,��B���+i�B�!�B3�4��X��8zT,	5�QX��wm	���X<C��������i/�T�EB�Z����nh���4)�=��u�ܪ-��bZQRT��.0yaz��y�y_�)`g��0=���:h�����Y7���G���f���gUt�Kp)s&'mgb���S5/����pːa3 �G!5I �5���Ӗ��SW�Y1���|�Z\��Q��p��ǋ5�7$����~��")�lh���A�������c�7؃�0�)���H���	�ƛS�a��oz����1H@ ��2૟+o���
z�ݮu"+���#MC:�a*�JH�%r?R57+���/��1�^,@�İ��FS�Z��\�m/��f^�
>o$K��hnO,�9P]�g����UH��F����d�_R�M����(��#W*xr� �	�M1=n�&w{�oP"HiWP��i׀���ߏ5��ލ�Y�J�V���l���=k�p�HS�
)%w��+L�bS��c%�.�e��B�����l���<!�G�
��#���14-��ȼ�� � ������-��&:X-f'O�+TG�1�h���d�P|΃�U?ZZht�,e��k{�W3cțx1� ���Nz�J#�{�@�Q7#�ۂʯ�o��`�~���΁�^ޙ�W]���֪��9_��B�������P*�ɢ���pn�fʩ�oJ/��#XV��^u��[��@u��"�q��1�U��N�ʌ�8��BnTn�շ�y���mq��+�QL�T˰i��8�	����"�.���o�;�cf:�F�!Jv�F�W(C� ��h�駮����<��p�G�Xewm��15�3���\ez��L��C�ku�	 ����Hz�ج�J�'v��tQE��zwQ���|��ؓqh9W_�d��,������.�`��j�nؗov��D�B#��S��=ȋ��_;z�@�I�1c������j4�2G=��.d6<=�;X�2;.h�����v�E�G��f`�CĆ��DI#R��J�QFv�@MI���y�q�0Jߓ4�~����z)Ѿ�'O��:�侮����/�ތ�{O�L՚��\%�4�h���$vu�����]�Hڧ��#��ؼ�px@X`Nw%��N�ܪv^�wb \H~�!slVqr�it�J�I����Z�V��?$`�pC���i��	�ձ�P˖�� O'ٹi��"T3�Аs0���Ҷ:� g��]�P>|�!Q8I�Fء]��O����L�ƥ��83�o��̲;�0���z@P9�z�Ў�Y�BI�R��s��q�4+�3�����zCE�d�"\�])����q�'Qװ�M/Oؔy -l�z�� A���A!߰!+�$ۀOQ�!��?�s�hY�cٱ���a���tӐ�E������̚C�j��O���i�70-ׇ�bf��VR�t{�\�ha`61rmAu%�0b�gS�����7!�������I$�TpX����}�T�k7���_�Fǫ6*��e��zH��o�M��&��w����l��[?���'��'!v?���|�'L��C��;5<N��y��b�ɋ��]>un��A�����B�u����?�6U*��;%Ei@�����,6�a�2Gy��7%��t��g@be��֝3��P�۫!�+�@A�f܊sR����Iry���p�7���SCC9��Y��b�U
!��E3��ۙ�^�?zY�<����*dǥV]$K6֪��'���b���#A��hL籙���5���I���8��1 �P�ح��soR�������@q[�) gz��[-�[����[4r�;y=�����a@:�2!"Gʤ�[�R�w�˃B@'Ӈ��`g(�Κ�E��1��̃�
D�r������fv���o�n n/�(�w��zY �n�tH�h��S1�ċ�qc�������Ǉ��d���Y۞q7r����1��Xrp�H�C�@ =�F[8��pAJ��v=Ǚ�w���C����r�7ՑKq��[H���� q��+9^�Y7�!l����z��&�=Q
e�묰�Z4�Z|Mv��O��.?*�2d�F���{7ۻl�T ��:��d�?<gA��{u��'��7���/�n�q�]%��v����x��n@\/��z��|�6����崓��OeO��b�'Aa��D�"ۘes�/�u��$��Cj��k�Dnn��Ys�|��f_+��__@�}�E��\�,�{t3,lOAI��L��=�Aၙ�\r����&AW/��]y�H����6 9�[�uEu������[�����:�O������Z+�}2X����\�h��p�Wa�?��"�9l�\ *v~�@�#O���2�z*�;�%ŭ�2qÀ�d?�Ӿ�z�9�+�43�&=-�dmc,��]��͎$��tݍ��lq�HA���;4)��n�QmT+��XW�>���0������S݈B������
U��a\O"E.�W�!&$�����JKK���wS�x�8����[�� �Kb�rZ�7R�Ѭ;%�*��@	�ǫ))�� ���@�6�%��E&�p��~�qPw����RYr��,�A�8�Ǣ��%i������)�a
��۳z�\@wW���:t�n���y3�d�r`.�����]��n�"������
	��q�P(���k�_��J�>��ڠ�r@�< v
e���w}� x��h��O	���L^�Ɗ#��G"hbg%SV�$x��,m '������M{�u�}/R��	�
?{q�����D�촘5��dˎE*��JUo��W|����)r��CVI=S�%3�;�b���m^��uݔOjj,����J��5	)�b�\��D	
o�,0�IV=F>q�!�����mE~�f�O7Y��z�DIƳ��*�dzv�%:[J��%���O���P?a��m^���vL�D�	�s�b�e�Z-6�D���48]+����M����5ABȍO�%�e���gr��O�L
Ǿ\�ԟ	ƟT� �!ߟ�T���
'�M�O}ʩϕS�sNzLЩ�S($�	���I��:�p��htz%	����n��P����04"%̜ֈHr��v��p:��0�>F?mR���7�W��wA�>/~�#�NG25KX�`�7�'��#�^<����\��s�3Z�kjOr��.���r�����#\�28J����K�����!h���7��
ߺ��U^16��3�(�u���������ݰح�b���f'��h|�-��8��D���VU@�C�"�Չ��KO�~^�~'�e���F&�'����Y>ot(����*�rQ�N={�A�וuboh�QL�g�U ��y�'�V�s ƥ\�����J�}Դ��8삌8�o�U"�\�f��H]&�$��ftٰ��J"���$��V��d��:�+��5N�@Ă�6bw���эb�2��g��ysr�U�������wǜ��~Y��u�$�-Boҫ'��&� �r��4�:��!z3�E@npʇ�h��x�7�(]zpm����t�����,�L:�V�4��>����h�O�9�ș>�	�YUG�dw��ᵦ<��y���j����i2P�_d���ZR$�N�)��!�̗c�Іs)���a��K45ff�z?�0Y�d2'�P�6�?�ٻO��S���6̬�:kA��m�����e��!�Ȼ�����{k�������u,B��ӝf��������Msޟv�؀KH��D�P���,	.�ag��1q��i�`K�ϮR*�ǥdJ�Xm���l���RV�c�g��liO��l�j[�y{U�E1ŧ��=�%!-�p�ĺ���*!~��-�s�6L��L��l�3���FA7Rڣ'�Tc�������������-���a���M �B)�jba��\߽�g�?�9P-���_��aZNlk�ǈ�,C&��(����эT;��C� �L��<ʡ��Š�I�����_u-p��혈���|SeEfD�6���Q��#{ k憜��"��G���[hh�q47��3�y��nP�van*��p9��R�aF�.�*z,E�5�����U��S�	�B>{LS�!A�[�qN�';�HF�&�w�w��FJ����*Z-:�H�_�8����3o�)�m���2�����?s�P��#�� �z8��Y�M�L�;U7(ކ��X���whH��`���tx��xiA�����a���QH��i�8�Y�G&�	���N��L�Q?���)�Pl|�k��U'����\���,c@���B����et&(���k5�C-X��[��0�l2ǐ�p|������//,�z�ŉ����"�4��H��}�h1_�V��*��r\k�"B�d�������Z]�'��=�//��O$��p��)��/e���