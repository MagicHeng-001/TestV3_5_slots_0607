// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:10 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LoMAY8uM9Kb1kNzaZbR9xS5ZSRNiElNwtJK+9qqfsk/iCwyqgVWpN5H3+KwtkVs4
b0fiN02dslD9QZOYOV7p3T6xoBu3rMqQtyCxWouQJRsoXVDn+jaJ2nmnP821NX/3
mn580FdpuJLD+s/jEMLUBeptGbydXs1WXRgFmhmz1nw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 103552)
0Kg1VHjkbBFiyIytrN3BBV08MRex6UYJinaggSUU5LIfjUCOWZvYjZYqd8uavGPC
u0+piY+tT998AN3uxIIcf04LxBUIzF7XaoWR0B/wKvgtZLwVCYNXu6/BPR1H7XmM
9IFTsxKZU0t3fmkxx4CinVO8q7JQZCHixJZ7OF2WSYswpH8/q5CopXAGuVbCmRQD
dc/joCEBlvkxsGC061NywIYO5AOeW325eV7XyDmH479zDq0wbvisrpG+CiUrdO1c
YhePPtXx6c9PXuxGoLfPwcZz+dLoAL+KG2n6SiCR5N3JFuyjgKqzNu6Cydy9NE9e
KrAmWcgR9xbhnJ8NsVzIiRyxm5y7EafatInkVhYagDMagD5fZK9GoDIlnlAOPMUl
du2uVBpYsZPrGXi58Ua8A35Kh3V1FjZYeid48Cwd3JdE2fZYHH+4FGJnGq94Qc1Q
yzKBHB4rqsy8HNckbRfycFdT7ToD12zZEL+kAaTaSeQEzbr6hXXcMhVBzaoKVLfm
jsbNUg1IwXRX2L96uOY1njO5j5qJiAghgAa+0AS6BYoH5pFkXIzr625NAnqkWLYr
Dk397UKiFfG7G2PIHYgwR9FfbNcZrR2f/mpFdNgi/RPf0ksftsYcbrtfpNHo5eil
v4uCbsBNKGpnMadStVf/nTnlIaw7kmEPSFA5hsZyHtqs9aoaHerBmaVzA82SoiCz
92MH6Ku7LtctWwQD6eD6/x27xbcyXHe+68HT7kSPt3eCF1klJ/EfBEAvDAhl/V4x
/7tVXSrxdLKXAmsA5e0QRiPl43yAZxB9UV2tTT65YzO6Yu3n/vsyy75MtDCAMtpL
6zpzyhG+e2R9R+/WY8VG8U65PDAdXTxp/mw8qlAV7VYYEUrPflv7xk8mF3BfwwuQ
ZTF7li9wU2UCOGrA63mkeEkW4nw0spgKAlvGavvp7m1eCJb1ciAjcLP4TEU79vJ8
NnpSAu4P6CA+Erbs8SvUetXNcZ8GVYOJBCMzd1FT4ETIrtRgNxecpg8Z2orR286Q
VMmLtdknfQkbruyF1L0rKfbIx2A9mcayBMFFKBqpWjUh2Cx7Apar50G/pb6t5Gbz
oGXDY5aGvgsbkE+HVXx8zrZIGZ4rUK0QeiWWJnGcMmUKDduZq5YBrEna6NUPlCHo
Jn5vWQaf+w3Jm8dCTlfWADyNGsMVW7LM7cfTEA0ly2afWNxPqX8LvXbyZPvXhOwu
iTi3NF8FE1cwtsbyY8gli+z7rvyY18aT+R0TQ87HEAyzj/5iegnIVGfLnGnAGqu9
vzxOG8Qn+DAJnN5fGsCNZkCw0hB25hBVGe93041bd1xlhF+cubjsGmgzSuw9A99U
iVZCNYC8SahMihLOTmInnXdjN/D0gHr94i2BiV/qcCom/YNRJgJcVxEQ6SQBMbQP
Iczp/dEe+wZvdkFlKtU1q4Jx699P+ttEU1XPkywo0JJ5h6zLU1h9TR9JkX0ITSQl
DHzCmL0ZY/QhsvjhnyUZhRTL6WoNh8pqyAGyFXetTvTa/SpHp7z6LEUzYvLBUODy
4V7vHvciJ09bGiu4OUqv28fI/QR1bKw/lYe48Ru0CHZpIOMt57cQXaGmmGLaiUHz
s6t0+1R+i5eJb+72Agf5jEewWgt6mOUBKpK9weJKanaif0evxzTn2XyFOKrjiBq3
tDeT3agunvdeaeLgy1MRwH++Oy5R/hkj7V14JowYU8CNGpGFL3QTy+XIMyo5xYFS
WIflg36Fq1D1E8q4Cz3+0xjiHciTIxTDXcsW/KECRfGrwGAyVbMDEFz8NQwEGRoo
+0ABqKzmb5M/iwEkDhIDDni/n2NzjQOA4PjeoMrJEzA38IlM2Bbv05fVHLQZq5QR
LNRLVjxabw+xPw8gwqwIWDizj1WKGgtQPQ0Rdm8ryU4FWNWByZN02Rp6VBUhMhhX
t18WTcatFQNQmQDE0Ybfa1dI2MExRmNXW0u13m2F5aPfbzCpAbJZRIChUB8Fo+eA
eYVooOse98RrsGGhb+Xq4NZvryDI4YmmmSFxksJoRLJk5DS8BTlqbDCUvuOnOVIq
BSpKI/6/RHvpbR5NpuaDTPwqJ1H3jIRyL+cxV2WqpZFi+YdHb0uWJD3WFhpFWvWE
l2fatVt06DDPoOl7BClhpd54MCPh53a6c5vaVG35bbdtpIsLOwjX22zzH1E+IuuP
YWuMcxbX7FpSptW8eRMy/wuuer+EvcVkKepm3UTGEFPsUDChs1gM6+mPA2TxT2Ag
OFCgrc4L4VU2YpDiuMIIvlQe43Pw+xZsENYMY+cngcm4CJGbMQKRKoC4gddi+sl0
k0mhA9yZMM4X6TkYkdufAV+CzpM1qR4dJ2Q7z36xHGefZs2zNV1Sk7lF83NXsnvs
cbs/YWwNDUTedrzN3wTKQEPHQQ9Hx2XCABGmib6lUy/sc5UdTCKM2oNnr2fykDVY
YAf+zxemzwA0bLJ0LSU+XbMZfhTl4bU76itwz7P9IkkQf1UyhZFa8JeDZA6DUgXQ
em6qEeMLa98C2tQCmFn6UgqSPJn6wnfNmfdRpo/SORAZhT/YgDeTTcrfGNz8zNa4
ABOmO2Hu2hE3wEc+BGjcRFlhjJ1pELcqawX98nIr6qXDqjXBgxz+ZBF73JwqkmVP
qjD0NBQB/qAnGDFljgLsBOdQZQAp9agRlXV7WKPSndnpDfDINNwU9z30Dk1gqOA3
TS6aMZB+VaeLvSpOvvtPCyTNsjY8QL5BNM4u6C6zPdzNzpORfm2Pvn0wWjNByAv3
LkyOCu+WOxIK3IJHDhaeI/JOH+uIi9PqGwd3H0itrJLxvGOySyQaO0S7rVQHbvPS
m9lL1p9bM3tI/7dvFKAAtBkrV2A1XBXHVMnYeq6+KXX9LvOeHP1NiUrW76gS+P0X
PioxtGx/BypJD3RPLzjzuz8faLvQOcczN6OWvI0HMS6f51Ci6dLnVtF3t9vkX2YC
SL+ozzX7YtYFgrhSaRoxAKfCl70yLW5ZHpH58lQg9Hmva0476mfV0lxKfyHdHCpa
5w54WE1LIHQ16ttksOA+rMxfzTjKRhrhO78yUqtPlYmyqbjCoa+gp0cK00ee6hoH
x5NECN/UuZ0LTrW9glAaRXNfTRbEpMUndcq5FjpQsBgPatPYBo8KsEYRxHcCjPLS
Ixw1X7bam9/ZT6O5xrCDRGGrfg4j1ELTEtWfmfDW7zDLPu5/+4aNUUZgrOmnUTkc
vKzypq3EzfPbXLU08XWbtgyyMooQwd7ORMIwEehqGfufLGW8fwG92z8M+GUVcnEi
Cq24+YUpyE2I9QeR8jhH5QTn3j8/kL+WZOFNzCc9sekbScv2h0QpJzwkIshD+C7N
OAoHXugX8M8btwOcW5g4Mf3XcOjAzmNyJPWTOvAwxL6BU2b7dv5wbAkR6CiZ3yvs
+nFqEhFzrdYMBdrIKBaVXYVQv1cTcdJe/5SnGCQ/ArJdBTTJoICb6JRVd++2MKbD
9YqWs2Lj8+HSFX4wj7UCKS+AoJD6Ubr6o0SMJJRCygl3gHwmGMUpRvwJeuWR27dj
C73NhMhmTtG6Quj/+JgSfhjXA4Li4ClEC4pWL5jmccp8kppLOpB9ajHerHG2Shin
gwgr35x4s+DFCKQNVTOU5OXij3DoklLLKdtuLuVhHCPSbU8ymRXZ0WTSxDpIPhXl
3dgSQCjE+sGs9OXCffMwBDXggVhNmwhM8GnRg71yfwbhhRrEVBtsn998/htcV+Y/
Vc1pdVMqHd/19ufoV/aukjXK/XSXkfxtqgOkjFpUrU0NQj15b+xNNdIimt9JeIJy
XhVNgVUQ88oWwstW2o3Tjq3n3hKixhItg1GusDB3BXg9s/gkRonNPy2P4I11fil1
oAZuMLDnkirX1CxLbwvt0A23MGX+9DN4DiCAk4C6/pN8YckUyGdqKOtQaAnVS71+
Rb1OuB2zg6O4tliDcE8k1p2YqXuEODtH/gFwfEOOBCvVTvQwBkXo8IIOn1WbF0ae
7bDLX03ttx99ZHSQcB8bWHP4hbu4rqKwvYSaP7wj57EavmzmIo/OrvPkj9Ef65nM
0JSAv2hqL1S9EQz8q/qZ+Cno8WHyiJgiHIFfNHmA893kEaQiaIUoFmb4bmLTaQzo
zmN5SCpeGdhNgeCh6v0e9k5yEuRO+dhp5Nn3f9I756oEsdX+xPYA/KqBiDKxYInW
PmS8XIVvpgPqeTJxnfLu8TbVGqfLNsE5emv0gElqOij/7AUbz+AUL0rOBQQljxAi
q1HYA57R2BQtXJ79ahn5BuOJ50P7GkkKTZ7uxq1ZSlqUgEiitU8rKvI4jr+cAd5k
8B1w2333OQnGmJSM/WO6isE2pJC4gnMrdTxvv0/z2EFxUiZ5+wWbYTGcFECWXH5L
HO+84KNtSy9JWuzbgGznR3lT2NvQrrMc3VgMqWQfMLWXtVz9U1+Vx0s10gCD4pdI
BB05Q8u0vxvjv6goxhVyQxuaUqsEh/EJr9ZKzeXxK4ZengZ2UyFPIzpt9lYyA3jg
xsdTu8OguCaj3o0ygUEhKz++brmol2dDVYgkPhFLkpRWyggQK5koh4h9UMqtzke+
pX1A7dKDcZXE2RmEd1eXjsdri624MbWBHDPuhgWrDld9QykyONYn7IAL/uyOfd/6
1cDi+OkV7Hc0Blhhw9QvOajgNljQfvERwQiKhfUm7oCVvui+GgOGPX7Onr5k7kKg
43dkBwLM8QKc/aXJM6clQ9jL2zaLgi949PPr+MYjWrNaoaAAS8KwqEKiqAB4DfN6
6Uo1YEcHtSB8/MkJBV2aTha8QHkaegAJj7mNQnM50+z9/I4roKf5BGGve59mJ8e0
E8dWeh5Ar/0uOtBmp4sX9joE/vyADHj0comoJRhJz3jaad9Y9D/RIjT0r+WgaaSh
VzcYIkXTA9H02eRT8yQDGOywZlrtsz7eApyi+GdiQQDWqY7Kbq4K4/KGDq530Sy4
/SGYa/zWE6+TxFvv++I0z2DJVgzJSM0uCyJPXOSn94BXIB/uw5Yv01BNbioxRxqG
fEydwk9+/d4fHbkmStFFWflo8r3Vr364hmbUzcmNpf02sYoIsW6P84pjE/LNmGPS
AgoKQeFTjn1+LmHP2RwYh/HX5wcfq/letkQwoxpnJCEbgOxjctgtkT3lZoUGxVkR
lRvz7mN/XDj26T2XhL/Kc62qCJudLbS4DHXeoJGNP7R8CNkh/XrKXL+wvgBZIUv4
fMW+UyoT5uIEl5liI9JitGjshKpTYo7cGzMDqgtDo+9HsMMNPlLwaJ/lQpyFnQhU
x8LUq6g5J0v0UCrLsg1KkX7I8PJbx3n+kmk+GNJ8CzvzQaNBCAok+47rexB3Uk+G
Z8tLPG9xrBGqT+L0v1xnuzCqJW6dTK1Sa2Fa/01Bwrz0KoE41CXIbE11y1+0zpzp
0KiterBdfFQ07OvMWNq8P3rE/rtSlBb42IiqlhHSEKDVYytQNeKu7Rlx/AHfyg1X
6mZQRcDeo+zvx9lnxCkN+SDPpuR3jUgxWk7MShvjkNs5zy9mEyQDhHag0m+/hfER
iVYSCne0e62tMEqtxbNV9efXjNSWIlaL57TlGMSoiKym2sq8TWm0aJnspKKXeKh1
c2aGFXtHgNkrD8iDnQ6IVPsqAyDDUKCHoEcUVcOaL/sh5caW52s9sRsyGYkeRo8p
MxmCR9kqJA6miKQDweIVRu6ahpD4DlcKlJREu0DfjEjPOyTwp9rch+9xQCBhjcd6
ls4Fik/MFrjYygiia5TNjAN2Bq/sUM3Ixgp9hb/IzgBpZkBDcayVBtJmjYQorV6I
NggKsfF/nsL7kd4R8bhX4VDTb8tIm9md8Om/rQz4jkXj8XgoH3YwnuFHfzaHe8HC
/clqDMG2xSJSp0RH0K+X8qBapbuHfsv27Be/TsnOkEMewtUnfRXhM9ksIOOONv/I
6DiLJy1lzlJ0e91VOaM0/JZFN4xXRX4z0ia6qDPfBF+eGCiNbsObih4KmTbN9uT7
bV+wtQiYOVSiNUDz2aGKrwEYoZZ8BKbDKQCZI77Nqi1dPQb2GdLoA/urFeMDUwQe
JLaAWBw2QpgIBxEdxlb6BxxkiYPOyOm/vr/Z/JnMBpWd/2CqRTGuB0CY9vOhcaYT
AAbNJTBSOqJnRxmTR5OP3jxqkOLCbDyQ6emi060ZDs4S+KXlsjD2jDyP5cdsR1lU
O65nlOaZtrxGfwOnQ0kG7JBKdEGaFV9OJuei/lUc4ncP08VaordAvrOtTI9cCbox
gj/DBYgvtAQ37MJ+GxWUEjo7NLWui3gOiULT1wLT6+VWL0dE0DwG3hnp0oEIplc1
/Vj4IrBT3klhPNUiHCjwInZ6lTbFyrFJTGluSGrevKB60QIHEtJl9jr/85dkZBOZ
xxWhtK6F5wbfjsfz+XCgvI2qZWxeMbbA2V7MRg1KtdSkXpu2AjFtF/AqSl0Cn+9Y
OBoAVngKNo7bJoNUa0O42lJWRASuOIB9eWY3zxEyNizHewmqZE211+j4IgxeHgo4
Xxho2GgOZxAZVjhrMdkyZSmH8tKylFGSskJDofygylsGg5/WEd9xVCPi7hFbIgxG
RKvrvDu910+imYvdzyqTTOlB3L7tzJdtStCOAIXL8xkX+kpDbC1SdAUYoqw9LDBg
AdCf2vq7SN0aELFyEg6LiivENuIr95gKLRAJyp1hv1/qnBUxwP1goWPPuN42drYn
97m7OEsxek4Nz8ESC+Q+pT28fI8WXjIePxfYFWyz1KiqjeMPXOhl8LZDTaTLxzNR
gTzMs1u0j5pfkMXr4Erx6DWW4bB+8ciQVYFVnxWdv8aWhsk4UVCZjpFMwO8WufAf
dEODmTunHloBm9byTHfaJRkXXE9t6cwmiMobDumaFj31NIDMhjExUvXlX8UG6qkO
VNIeSd+ELpTUqJBLCLMQYndAmyACmOmlLXgnyb11INPv7yL9YdfLSVEYAtWr4uAx
b+25rG30wB7aNE+znzT9I66ZGxXkhbUlDtIvVkde5K0zs+AERXeboo/DwjJzVqYS
1jCVE6FbkX2kv+qipG1wKFA7Zy0CjCGUh2oz76hCOUx1Z2vUIxPoBgiD3ytF5mav
qc32lMouCXY8DRINHmclte4EmKXfvjsT0t4zcpZxYxF1XiqEVebg5l+J2FkRKSMB
I+940JPJeNK5FPhmWGPgdeJa0GlrKUfb6Dfo9utT7Jt7a2NJjMm5rAlZOa10EgX8
0zEcLmM6QHIurRnVmvvHQW746+6oWH5RQGHwwrPjC52X/yAd4BE95OVIJ1hUjIVG
FDMTcpf041shmNk8yFp6KNzFxMXDvjJXm/Nbj/0DRTyljkqpz8vUpO/P+xQBR1R5
th/IlmKXanB5wrt/PBcEag8UKpHcftekO+QkxVs9/PBrHVfXzjoisCu32v0E81pu
A6YdZnsCvT/P/sSxFVcpPJRM4tdTvaW+LpNNrWDKgmXo5bDXX0atthU59GrYjIfe
eU7fdf8n3c9yaqE7QyeXuqN8W6RBsWq07i23ePwJ8+AmJTCqN+1j1UPaxsAMGCzF
ftcSC3kCGMJAa9KYuDDWNm2CdonaNCsxO6L6u/SSnjUe4eAYvL4p5HGp0gxLJ5dF
itzMQqx6cXehFIeXq18NqfuKXlg2yVf0ncATlS+g3N7KzyrPNZuwsCf3yL7yXjti
x7+o29rnod7v+H3Iit79axNxAlI1TN5cycI3XtUIa8k6DiI9ERE0jW7BT1+kq942
uBmtcUNLKXo1d0GfWzbNtw3s2IjOhDvb3tydNrGNKTQeP9VCCyEdafU3xhxBREaX
6rst1Pp7PnrfkcXFAKgn3wJne0qG0KUYhOrQvDxJpcFsF2CeITF7VKd7Qrpm5i95
U5fqlesMANme3NWdKtaqGJha3ofG0vZcOa11ZALBxo37ziksmGcMfmFNE2H6DXHV
+3ZKMl4qPpQc0CVvv+xHi+jJ4siaBrTCXVPH2HeG32vsyLklP7ppyNImVO4s+Kzt
X+bibVfRUa5pRt745pcOJM16tIxkBYqYdcBeImgeG574C+x5f85tKJQKUQ4XtRvQ
Cjqm12XWlAcrYlSD3Q2Ev4HG2EU9309cUc4FaqyugQG+1HU57PeqAQl4ZPW9k1cb
LFil9fM8/vlFNbD7tEgGQH2Ou2IwunUI7l9TA/ER/HUfsiD5ID0jpj3luiFRdalk
Xt8syDTe5f/EjS6eRwwZIskhHOdnDJOPGKrT6+tvZTEIm9oEhaHCN4xiZaI+XMeK
OZ3mdqHz2IX/NbnmGkPqAe6EYxQhI2MpR8KNspAK392czuOESL5v4fzMk3YM0IC8
VChPTKrmD4q+Gi9VvVyOZvcJ23MZlV/Ng32+S7xZ8+OfIvp3aD37X4lTLOexz7KR
vZy63RkiPedBr1K8fzevrrT2/80/alTWKsiQtQ6Pp3aPVChfSEFmJ8liEgk75Ecj
aVAOBWrYRnWv28hNnoKNVakqOvW6unqFw+pUCGQ7OXGYSvlVp6tUv+zGT0JnlcoT
9ffQ61mozY+9D5rDi9yqivE4Sp2umUZSt85CrbKkpHRZn4idzy3PXYtPg/2P4bqt
THNCS+CQZdwokhf2yMKRhrh5GnpRr5NDu8J0gAn7xCd6FISDCRH7TOBvvqmOoz2h
Th2hM3YoVx0Sbfd3lLMR1/fYyCDfI+ALTHJmdwPdFSsZ0lBL8mwCdiGal7yAmV40
3w9ZmFpIAwuIKL4YRyc3d6a6Opn8MwbECeYdwkh5yyz1WMD2qZbnO1MPXe8Pncur
NK0QnwGG4MpSh4XUK+VDQ8oM/wl5e1BOgyEcueVRst6IlxMle10AMOWhpryw0vQh
U+pihVQx6tcP/nw7wLJPNgjHP9yAvRocPIyoapYP0cPROtGqq8n57V/G/5CMMjAk
zWvyQiOUr/IkD+KNQqizvvd9rlIngB4MITtjrWrQu4ckRo4HAD95TZtM1OhGKNQ7
xroCdULvctHJmmNQ/YBDo/sL227Oju4G4Y1sSesEZvYNo/mPgY5TiVmvsyGjxflG
KjSrWWIqLfwqbwd0x0yXxq841eDJc8L7cf/o3nK7BPCxDhKuguflvdf8ZnmWZFgR
xxweum0Dk9ZAHvRDFwdDd4R25d31y+TrgheKrwzRcLTjoguIQW3FCVwYBFgbRGGm
5UjgLkSojFRKSezFAnKQIl/AkICX7xzeQc7gei0fyDxILvcuXmbGF6mKgAjBRody
5cSVAeRMOHuwW2pWaonEKRUkDlZwO0OsK6ykRpoQ6MyqRbEzxpGyzctSeY+W7XVP
8ADx0rHtYbKppuTvwOYZQ07NZQvi9aevxTQYuNg/EvpWbDRUnAhomM6KYgVVie68
DvdMiUt5DX2KCKhas2zWmtL6pqnezuSp81EtT4eBQmQzk0U0DzztURPJ1GiokZZf
RSxrI9s2fRwsW8q+C43N6cR30MR+n0uPIT/8uOgf8MClUpKPA5//1sE/zyIBnc1i
ElRw+/7F4lWEtCp++93KM7GvTOgMo2b8qjsOwXTuWMexPTrg4aD5OuA3PpM3mogS
cK9TNWyOspK5kCYU8XAJCP9dboGQbeN8OMyh0tGY8GpdeSBX35/Qj1fI88HHClsZ
9oilI0bV10d/QBWMiAq8pN8mrCEa/exTUpKeSBL6F0uHH5x8G6SFbIRG6eg0yWlm
PJJh/ZoIiB6KD+dd5Aed8A+RRWOYcEYnDHwXHMJohsV8TuBlUK+MU+Uyzgoj/bgK
Ngt3uFLgsfxgHhU2myf0saoMo91I0f25FLlLWm0PT4hHb3N+YM5Vc4ltjf1Tg/w6
R6Z5ghDw2aKjqCbiHYUzX3RGVHt2VWxMqOPVx9Fu+OSgdvBJre3APnxEOlz1jyO8
KuLd1JFkFWVXmspsEBAL+Fz6Rdpb0VEWCipoES9A8h7Byx8HpdBhWbOLvf6tipMA
zaXIeOW1hXPnlq239fPU26ScH6pcAe/2+HwcqlBdPHefNKqeiXN/3UINXiCdCoWV
j7/pPYgKICopQADELIqVaqDkjaIgUG2Ls7gWFB8HHEtYsZfR+WOPQJQ9UqVXisyG
5XsgZJ6nIOhrv5+v7DVSKPH9cHCbwizq2nRoVXIk3Lu8AFaYxq1R3uoVr3PG/0i3
NNtPfZ6SZqHyEDDPgIVBJ1FR02SKUDyn7Hok7Wsc8ajLN/0PHcc5PrFsY+LF95Ke
hbva2uDjfshncCeMtQFgnlRva12DyFZcwEncJc9MlfVkKDbaKb4OizMtNZ/5IzwO
mzcNyoRcLwOpVjAUrncxA7BpmpXMlS+AUrdPHxPpZ10FyZjEd8jzyySKro87vkfB
6T5+SNfhLim4d/sW+VylkdSTwwC/BqaBVzhsds8iRP+ZUy06czvygEJiDLspuqzD
5ZKURSDMkuh5uSvCB2AyBcLkb19tNfr+KWfEJpVyWj0foL08NVC4an4OZNFuqa1q
CUKpmG/XYX+g6GoBWSms2Ke78w20BcWommt/navoFaFXNpl7gMYXs/mZ3QwnTEwz
D00GplKhwsiKS8x0zVXYEhLStiJlt+o9HAMhAgkOofcH27Lu0tfF8k4r2alODPyU
Wa77o1geYA5q+0fWXnhwAxa+qRCOkAtQa1SDYeBey6jobu9y9GMbxEysiC9xhpvS
SFxoGRrxqW3jSlmWQMOIyGdBYg5Pf1QGZIs/Je7A3zqIAbJxK0vq2irTf5J4RTeG
Ifp7zGKyCf4ci30RFrdRWaR+eP0oJGR2UzVTYJ+8l3H4LQ5HlhFFJMhyksVemUGb
c1IP8nDkGWSCvw/MtbUH4z36B9EPxRA7qePVovMloKg7hLe++WyI4Z8s6MjAiZej
hcL/Abnl2MfXnCWda5ydgc/T4brDXq1e4GNPfsD+EnjJ9SxxUYYKxc0zNVTbFaWq
OBagC5+fP4qBGVjfM5FT/XX4DCdrbpyubbeCrg58AwHjXzElIekLw4mL+m2pxYs+
MvJ5WuBW2OJg0l5sJNxvx0Io6kMjJxcIzdU/9ZCvw62sM0GJHO3iEq+1QrUl5dTI
4CmlQYSffnz0RtqCMXl18OTwQdXOPgUS2DLLai6c5AihdwSErwPgJ8TSTithAIfJ
uyU+rkSFtH5BH9E2jDjlHzR7+K9V/EDTcwLUKI9znelNQn31eIu5VbR8NmQPi1p/
FnZQQ5qy70+LbJSeXid1AjrIrkUdLaaeP0gQfWEbua3ow3q85Mc/58HdN06ZztqQ
4NmR938ghkrFr2n3SZ02oTxcJgHvYwASgwImAcOuSN4j8Lin60TjSVUq3BUmc9xt
2SH1SmjulC60idQEMfhCxjOfE6IBFf46RXw2INMB6FlM4DlOHWrtBPEK2hqDdc27
90tQ0OKXkD5dIwh1TkKd8iQTjID9Cy41CDIT8x5LyjhmtOnLMwhkL3T6zV2l8DhW
L/GTg7+OZVgsdY3fv9FXuXjcLJQU6trSBK2wfEtnByBBWSE1yJsGsQT8JSBKihFv
KOWrdRVcMvC7LTRSXgh9YCeIQOkN1Fy8gjPZXxKzAv7GSs2hX9N5hWfmjaW34A1J
hk3W26I0MvCo0miv1CrGNX2HgWyZCF+tVRXj+LawS+zZL6Og3fdP00E0syupvxa/
6XdNxpK9N8A6CBfdCsayY/Bx8zPjHsRcwVrmgIXyeZL3DhX3jyGn67QKRQezAPq0
gXfYrCv15wZDv0CmpJ4uXhUOYxHaQ7LJwtnzuWfRhrXhsofZuGHb+z9lFnel+Np+
T5KSVKIZMjrD96yMupuAMDId3zdAa75UpX9wYLnd78hrvSeQcX3FxFu4cqoX5CcJ
crGblVYkJWk0y64JpNoMqRzI5M2evQYO9YUAyllKVpwfBFUym1EWNUWXrdo8HJnm
Q8CIn+lZDSGvApKK9Il5aRF5kt0iD6JVB5TQLXOtnn7sI2tJR0Gx1JJ3YSQigvXI
aMmkTCwML6HO9Fsxt/DFmVO6a7sa0M8QB5ahA4DBwnvWlHoR22rRBF7S6wX0ruea
G9NqYikn1OamZkxADGM8lRluR6EDN4KbcC7GbdU+xdYjdQ9Ud8I2hEbCnUJfDTSN
VJEv4U9EEJN2v9KQFIAc1LjdfhC1a/600dG5suq8cousr6hvr8fJOn5eVumr8ZnI
89Pkairv7jCEaYrhkZgheimDBLr5h9FPNQRwv+3DOac5GPwPTm+1oOEk7/mQHwap
Xm14XBcJXT1/fF+B2CEb2hcUHyNicb3LoSwQGt3lkszCLj2vMXKuuGCi9UiGBbfa
eQtCfEUQCnLRX4A1nxHEfSpZzrp9/UBJcPjotkC9TyUs9tAg1ZYp3zB9Xy2OxXng
tHl1NVqsNhKZskDJbtnCaowIGz+5+i28U2Ja6E7Q42p6sKHBZ8DXkPotnJat5h8t
87cd5euFfVvAG+13ZVcfBuPjtwBXMb9bjzsuROp7WDL7/6fM0/53gtIGYh9shg4V
WiFXwN9xMS3SnWvFwyqYSrD0FxfBaXjoihLgyATx8+N6Wrc7winz58gv9PbZdQNu
XCb3/qaD6OU9rA7pflqvdPhtBRWCVD71MQOS7QylmhUsINGVJteBKRzSrvAQPHLf
BBXAczSw8AFmlRhlHvp1Mvl1wo2iIK1rkIOtuCc+RdMz6/DBQ9UXGLb7r0SyFtMV
+oII1mFIvtTyanVhy3Mzou3IkNgBuYwiP+Mc2VZtz3uWx+YtFIZJGYPsjRBDg1ZF
A6201qKT8GLyYXgscWvQhxrimPRMSpw/EKFOrYz/KwEIVT7PHKPSVhwvaW4+RYk9
SkkxgBR1i2AdgfKf2iZEJMZj5p+YbKL3lAynBlnrsbemxF9RDVIln/xbePoZxZ23
HXh9/ct0XrmdvMlp78FuoW9T1wKmAs1ihGwFGgqZJatsDefEzUCJLSXN1Djl6G2u
XJesPAr8pA2MvmhylXeOS1dotVdqqbZ6w0upqVV0P5SEc3Tkp7FGkSemj1EJnPuN
ClOWQRxUOEeNS6uj4KFD8yUmFyUgqtYhBPXym4n41nnXXzUZTy8ZoHpnFt/5czLc
u/eh1VfuEisj9zGKDEmBlunAB+rTgNvPe1M17TVUkDXdWQYsRs6rQM8S1v8lCgPe
13sABLkkbb1qjOtbDm+hWypqK77nznGmW0mS/2qrx90VlZjksODwING9f5XLROjV
S/vCC2lyk+oeSFsFxKjnrydHxRTnXd03emP634t2DhZPhLDU3G/QtN8Mjb8ogPHy
w8OX+2TZnnTenWLXcJgRMrgWdUE3g0MWyAAUVRZT1211jF+fHvF3Ae0JXqQnHGmX
c/vdNZrZ+K/dY5sGl62cs95c/dfqwVHdj/WFSH9ZyLChyyUBtpsIH1qC2xmKi9kd
mRHZfi6YRFUftfsYRgPglNd2TKK8FTwDfsX7zGxJ61jUwXfLbFg84LA6a1Nq9cll
etYQaZ9CBlcSY3A5BC/ui84avzdTtJqgqZUzLHm+1cEzWogxPuYZXa5JNCnT0NoW
BtBACno/V3Ka6+tq6PSd2IC45PjN5dkZWjLeDzezfpTLiRMo3Fx6CxAmWlSGOMYE
fxXPpbZ6kiuTZyX93fyeK65I+HdXmn0sUHa+2Kp0e7sh1g6h9eQ1ed1t0Gn+f06+
V0mhWIUPh8Td05aacyeDrS6doE6QEMdpN5VdQWUcAR3sazLeK6wr3/icI236ro2y
A957hItOzIWFQShLYJfbvAUrjMQinbdcCItJoQBsT1Ii/O1Dne/5SkMA3+QkUnN+
YE8kAcfx9OeZr6ioCwlUntPhcmqzvtRCbm/NhM1pgIiao+dZmmm1jeMAotPkddxr
scVP7sXA8lrDuswa/yubu4NI6BPRq2bzKZ4eR+zXS++1DbHj2C8sddh+zoZeG5mJ
WDCWNdXkmx7aXV9w4hGP4ythR2CinaeyT8ZSfzi1wSXfSyHc6kZdLPnXL2p/4bi7
8jf7fow1yZlRBQOOnqXsnbf6oqSIFTpCB/OpjpWxJRGZAL/c9PxQ60yDWkY8o21x
IiKzhoECdHX5W1/RcxhlL0wj+nX7GsZTAu9oNhzsQFiSQxLoNBTl7PudkIb5ZrCn
bGAoJcSNd6MDb3akpyhICgjpWqqCzC97heP7R4liQulStdfOyfwMpoX7wkzbGuln
OBOetKwJfKrfAYWkwLKfeR40U4VYV1p+OkNjyjlQxdeSXPygHVxDo2ogeWrvyOaT
daFbjxMj6SVPH8xfxUGCDZLKl7LHhfTLX7b+yvhnSij/P6aVNcJ6d7AqycbrZQHA
zznSt6L8vXvXHI7DFL2OOvwTromvTQHzkHUDsh4Rnx8WCAbwkG59Ubc3YNR+2Y2q
nJI+E3T5io4ByMQrSJ40Z/iUXH1iv+03E9rzZH39hGLZtzTgUPwbarOBdXpJvZxT
on3oJCsIYwoWYaIrfhKiyeQ0REaqj5HMFeDOnx2nqfbxrYStTU1IxTWIKI68JmWT
xI/ydILu9l2yBSmQqt9Kt0fURCPZ42dRyvNWUC/PJGivUbpBmZeTgWg0E6+4DN85
T7AjHEEzg+LIPoE2MBAWcwGcu+kPYyBCt78OTXzzBsaZLZKDCGgEVUyozyQvMoMY
hN7afjA2Wy5YzhCqm2IvMEEm2XM4CPPiGGdv5hztBMJ8Mv6ja7oqCkEkOxthLQwi
iAV9yel8idF83x1lUfQSrJRW61DIslRXjUif8uob+yZkkeox/wUXRQqT2v7eca4h
bmkA0DZIWKRG89J90mAyWpKrpwl2rQP2TltnO4r0GSPpsyVtbP5Kbk2KhVV/vAB7
S0BDykT+UIHpyUvtiTT7V+h/CmGgxlyoxAdL9Sy1fpzG7Imk0mxb5cCDrFKrH3W9
VPP+8MDBhhS4stKyxjmPV2PdolTR0Op3OgafO63KzspzidKHf+bsi26kwsig/TCZ
E/iT8/w6fV2vpaVRrPX929jbXfPB0H9dJKQD3S3+74sW8qBOdfcEjKh/iOlUtbtz
Xu4IxKJDae/qV7XUwmWLmOSZOYY95W9SX7SMjUJUzPvGHU3aDr1ADtHcWQr9rxx6
Cf1M+EE8W6DkDFgXaiqXX2wBAHS0JMM1kZ2Yzxvtm886mkpPHRlgT4A8gaoTatWg
8Arhec3QnWTtoTm8qzQWCuV3BkmYAVsLBIbO6cLkkTf0ZeVCfNWvdL2E03t11s9M
cpqqPZrrBkCKj9zGVy034JT73F1kcFYkIdtqPcdMr4hOpTDLRPX4whORU+/5u/Qr
YzwqY2BlOeH5sZi6MQlYL2R3mC/f8sZj6aku5Dfg9IXVNal0+QXo7EvZozO8pxqt
/26c0JYsHMLDOyQC4X91CWzOV1mbRDAaghBQ4RIKMTn7G3GqTKJ7hQvIKj28/ak7
obBdkxoy3PBtTXCSnrUo7apMjFLd65JL4eL4iS+sLRL9QRG7hPRrluPckjKlVfxf
BUipehVZI5qhd70DO91X0Q8o+Wirn90N7OtUExMSTXQsv00vwsFdOSbaEC9LNY0K
JAoxaonglmCun5v7J5pLM22XOUIDUWjgsyJNfOkMlLXcjasVa1//M/uOBZJCS3v3
L+mTEc7ukqyet46FZf1jlXBv3oz0YlsdLkW5MjDxKPT23yKc5BbxJYd2CpY1ZT2J
Fhtoy6FggQHL03euQZfaJ/rdeFCBqMFd1RdeElVqv4oMwXNOuKoDuX3Oa6+0JB6M
zMCVe5xO37Gp2DmRoT9UnsnZRY10YryNNnIy4pWGEVtU0YPyn50ZSfm98Zgsjv1J
142+7XM38Qw+VwtZ/jWbUJRdZVPQNIn0LxH9ep49/nGlhIJdOl1ZxTz/VABsEaVy
z7e0YPJ9/GJhGme24yXlvi5wfSK1dzSHsfqplI+dBO6c6TXyuhI4+rCWjEAj1a1p
kmK4hdPvoD68qtrxadA6PB4YuV+AX8En3qN/dyXEUZUnlxGSZ369Yp5lNLRnNAGy
2spVAdMbhC6oSOFYTrZ3W+MjsmAbmTTWtzvWAzCzvl97W7kJNW0jmFl7feNDqX8/
sxBRr7QYRboyQiUWIrQPArK2zQ1IskaX78QoYyPSnZMoBR6f6JtbfeObMpiwd00M
RA76GEuTUeUVrl10BH6Jzuj4ZOIf2Oni0ybH4dqPQ0sbXmJGiV1bUEfDYAhTD6NU
rdF0d/88/yDT3CxqpP0mkgpPguKdX76CXyaTZoPJ9uz1mecV58reMOsS2yUFeXO4
R9EuFOCxV03Zsba/sQEJmKUkIr6nlFsSLnlka+l98xRkriNrfsUbby39C5gNtZWK
tnT0a5vu5hhOEmEjtUKMhL79LI/Ecis3kKMRW1/dHW/HY+fFOSEx2rxVZf3RFq/d
ddMKczv64DSgUAR2amvxubl8HNEoeHg0FbD8YCJeM6PInojkb6xXX+rSDTmjEWI7
3E+Pf0NxYt06tErFiMdJG0a3KdhdoIPH3Y9aoZia7JEfUj/3bAgDl7I5WnR6Q/+r
SYdZoD++2PHA96uslASUdL/kGr7i4fswBiF/EwQEfSAo9nZ0l+E/cIy9Ei7hjqL3
XwXx9q8v1DVMDcX2VUGfuYp/nVQTncHl8y7abm8LpkvSUbv2OB0IeTX9HkGlbe/Z
93H10I7ys98kzTHLfeJALQh4oZXQ2v/XZA3/ezP9zOmPE62VB1Mh7kswtRC+rnd0
dqDEDJayLoocX3dKxs2hVDieiRDcjznQpyltu7U54qXV/0TN0NTGZhdJArusgQHK
8oejs9itsiynXD9I6wjzkcpVPZXYsVdmT35TZJ/US6pz3wHPwMuEYaUTgZNWqiXL
VQg72zxXNEZVOPoDci++wBezbdwCkNGQaKQDTPJUSWvOL+4CfMYFmwsxx8Ro8/eD
XP4/Zw21bUOOUXw+6iRJBrgQNrh4hV4c1WLkm3K0Hc9EQ8seDEjoV2TP81rGxLiR
9obHIko05DgjRbS3GIysEBVfsn8zFS3cBrh8TPhfAPfS4Jh54pf/1xMVACZWnNXO
P1B40blB6Ec6hbYaTlcTJPf0C6TyWON5p8HTxo2eVqtpo9dyxGiIySdpS7Ei8OnN
fJKcgAorCARgodjtpXk5f6FlJzvDZRfAh+kQXIl2lVM9V6rttS4BFHs+ro6teVi/
yh/dP79OkwPMw1JOBGicBNFbLOFt5FZLkMN7jA0zVtB+YM3JJovs3eyL6biasfGy
oHry1prDnZu+LjX6NqSR0vTZTU+u0kA/9H5/2q9Yu1DS5IRaQTFuiNFSn7JXPBv4
iRuTNvb7LucjMzQYua8+tnxqaY5ajMGBWnUZkRFZTHRNljZ945Q/3+UjsHL1bUKJ
JTOKyAOi2562vjUjP/UtUpnFN3Lk1VQKKn7MZxmRgoInrfpJaGnddpvcLcXbbFkq
BmnhQJzv5H13O7hdLV6M1bve8UfsPCT7P2QjmroRnQ3AhIuBprbNrgGdZQBY2Ug5
tc2qxdrZbMwAwLx2i7/fD/w1WExDJwlX3jv4bzHnSIZUpP/92mE+haGwWSVGMHHW
rLTqtemARamZ5U6NtZRJKHS1KLv+wM6wiwAql71V0fyOwwktEES+/VaTWhaOcg60
QiG4pwCiC1MJ08HsqOa5RHGEuQQIPhm7ZCXydzDXshi0nh4xzQxr8uvQGlM0hNSF
0/B5jUvn1YI+e5vbfWpTwNRQ2XxMtvWD5xtzG3XfSq0o4bkEdx+gbXgNHt59GXMP
RHqE3i6wYHOEOtTnHBtvC9WpJEbetvEBMSyzjMzZc85ox1tTwiWEDFPhfFtngRUQ
aKBGnLNEXeEdQEEi5CXZPB+jrnhMZbUbRtiJMrJq66GmKAH9k/Nlceo69BlgNet0
8iT2heUUXSZO3fDzLCwOoRRqGp7M5kOw1+V3Tz/O1YD9/A3E7MOE7jJjv3WsiK0C
VMkbgQd2xPBarwfgVIYvb6MpoJpCJYks0p3TVao8NGvDZ/3VpxxoZWyeG/n0E8UT
u6K5RWfJk4R6X+VM2k2hZb8u5B0VWZJ1BMF0qmvhXRH0CixioqHh/0MzD5qHM/R7
F8LfKe5KG1+0unaSCtyG5Vq20y00XTOb1eBWhhpUiGuvA3y0aOwNFKFQd0QA8WGG
5Nhu697GVVHpz/u424NbaLzXY7KGXmL6r5pMnwK0jFT1Q+v3DnQ+PtFJtjJ4aXYO
pC5cVcdxDfBSQ5+y9hQtkGFrjBOsxNZ/rQbcNmHUhDaQfUr12CyceX4vQbYMZxIp
Ck1hZGDfnffC5GMJw5BIg4M+ku8AVdc07c/E/Vk/NpOE+tvGPoWhzH3MXaDZyFkC
72JDHuQypEsdTJYopwtEdfRPpXjl4bV7/RM4Uo0D29kNK4e4A+H+T4OHBOiswfcG
+j2QVuA9hQJoNbaAPoiXB47/F9mlcJVU9hLUTH479HtLHQp6f/t/R7ktm+Bo2X7X
UIYKxpzzFhkrWbIXGXFstnqae8AFnK7TaeIXO6A7ggcerUX8Dwa/X3DlJEvMg6By
mZM/+uzUhnPKNi4P9aH9KsOOOKGbkEUuaMnVCYoToMEpUJVlaGbui3M3tSqsMH5o
4oE+fqXE4C3Ysb4t1jhC9Sbbn0eb1sI966f3WpZ08sbeHvN3z8aljn3vqF1pfnuh
qaHbgql01VQ2BCcYvNHFIhr34NfPsmDlUpRYhG8Iv0RJWG7mmOnsQ42ZQDoa1LHY
7HUA+ek/tTLmwTSOf4ZzK1jZkw1A+V5sPLaWlQ8h1a3c9QqRMyG8jjS+1L0J7RYi
rWcV7LYtRiW1mN/Cuw5nTRCg1M2iLWe3/V+k3geLyfi/RO/1LunzbcOrTI0FzW3e
ZRvELGk3/fG/do6lRszed5ieuNtB604maq2riypmkl2UDIXpdAblOdImXGo1TC9x
u9MLPkrE//TeZsJob01Bhym0CwgURe0Xk6RL+MxxWB5p3RRMxAFXKDtXlqlHr8H3
tg8omVXdcUAzqQSvKvI52I6N5z0HsoLEQ1jes1p3nuQaFL6n+DS9JZO8MukOPm2A
2Jl+7XpQ5gXlXaqnY6ZFon39Oft4oPIHhZ4Sk/Uvdu/jJNl9AnSEk46TTTKrTH+9
NcUL24gzb++3FmV07cRRRNSfReLfGZfZ7S9Fv5k0UlQEYUeQMNpxuo/qLUpfFcJ1
NBzB4juoPM3E3pWnJqthlu1YegeBH/MCsT466dkho13wwteMnm9Olwti44AcapAy
+GuMPHuQ6P/Daq1q7Dk/ywAEqhzs7pG1NKejvZVWosR4AdEm8qh34MgO48qcK7BZ
Z+xzF53CPMpYt6mRKX27//kYTOWDE4zEf9sbt7x1Ee/Q1RoGILBi6DCSt55ENWlS
3x2HKIwA+GkMr9w8sPZr7eDXFe0NxPpENhVEXcuZWTg1Yrl3GC0QSppGwEHvbU53
TU4Lez96h/wKaQoG2kGChkZ2BStY99O2uLFeDQticbg0XhBJJ4VcuCXavSF949jD
4yrHu3gsV6au+FbTt0ee7svbrQfRZpLrJnEdO3Fsgjiqr01PjjwTL5R+m0kKXthl
wiAcWWYg5RUgF3IFOSERR5kwsAj+2QhXrKKl4LIZgivFX2S8UJNAt8vi/3KKhTSc
YX0fcQxw0+lXki38OTSftXzNFSf8X+ZDJ+qChV1rjvH9MJG48NYVYPGGWMEZYANb
JmYWuXUnHphCDYykjLi74Q2gGdQTV4B2TR1TUnuHq91SAgydE/j6fQW3JCKvDzFy
bWhr/Wwh89H4uNfgeuFzEXDevoB7t9eXXnteGdsFrc8P/9qI+Mflreh6v4kPQvz7
VbZD/y9rdPjf19dS+lGROz6EjFfkPZWDKYPKY1xNASf9TmDhyAXRYKb1OxlQnbPQ
FPW1JoXw5MB7QpxMjX2fYQslHLoR7KY3/tPadncOEbhqQ2FTEq/Bv76Phz3XuvSj
RpChBdIIcAi25dVv4DvWFLT5b8K+4W4BjX014gvqcP+kg+ThRU+lHieY0AjliYIi
fswcLY5wXjFxhK5T5NAKaK2afGgzQsWrNiaoBVHiWSvA4oxI0GB09hTuGY73NZpU
X5IJANnY9HT7BbFZQyHzuMMIxiE//bteMgLFNtSt7kiMnfpszIBlsDmjFsHBEPk+
rhILiKCV9OUyMJVyQrv/nOM+zy5MeY7cBPNX4vWoOUdgEgjn9+WJAjAptMRuWAY9
2RH0EStvjJiuFCB7ADQv0HNQon4QXq6tSofVQ0fEvuNkXTDzhjkGd2eHy35c4GCJ
FwZi+A8UcEdNq9f0Gpt3rs8a0lrMXg3okaq0sZ//4Kox1jWvkMXejRRzUAmXN26g
yeUg8lqQXSZI9b1q5bxFUXvhWLtbivMKT0fYSFAyR8CCKJeSa+tAf2EuguMSEEDa
G8iO2K/xccMdsbbfwin/sbjxx+fzAslBrkXsjP/OT5R0Y4qkiKZSzOAnl/Zjhtdj
08CWb0qYAev/+nD57HJG5jimsEBk2Loc+KeF5NK3U2aakJliEmtY3rxcSe82IOa5
v5Xkb+faQZUc8p5DGXeby8I+FJSgw0oeLBErsq4WIRKz7xYlhfQWuQLh6Iw+lEgR
IEkPb/NxjnSsmrg1GZXJnvKfVc1AIRQmKngGJaO0rsrcDmpA0rRu67oq6d+yqF7e
+y3RpQoxg1VeUrEwoU9I4XoSYG8Dd8V/zUCqoFWNhd9RHyICCJyHHbQuL80wpj7m
l86jT3Sa1SbBELn9u2Gw6zFDCoWrPGERv6YwIKaQXrlife5m2kT9tdb3kQuyhS3G
VMiUyXphlVVdzZJyEEeqsxgs6+7WcWQEfB9GfXyfCEnUPhJxNy8U87xCK4wTCj+8
nNG1c4nN2wv/FTM9BCE1IKAcRZZI2JEUv6PrOc4KYQ0vqeayx5u3mn7AkOP20R5e
4dJbJEyhC7535cUdJh/LiHwQy4bRZSyYR9eZAIhTZQ2DYFC3XU+LCxLTsRNf+Fxw
fOY/95u9scgslJHGT+KQQANvacOYBU4+Dj2NILnm+74E0yr8Qmo0S/9nzruc523J
Q0Q8gr2SpQYtYr5huzCw1Z9YIoWVHWPYeF0AWG2v29VOW0/VYE8+tRUywuevpHdA
yQ+zIl+SHDJIARABLppAdG6It3tRcnliDE8WRKOPBC60SRX/0aW3R/ZYJYOmB2TM
9nbEfuZj9Pi0fTdU3fAzUeBtBE7J9ksW2LvqGAHWhlmtOORCO5dZOFC3+UvIcmoj
rjBA3C7GD89MT/NbYOASmdrRG7l2H0bkOMVByC7OoTyI5mlzSX55CB4AUBo+Qxs9
Czmpb+H/5ilKCqtY5w7T/oU5JX82kX+Y+dgj6iQlTZK6zuW/6bNDnWj1ECbI/5/Z
g0oo1OKELZ2i/RdC39Zfg6fR/mQ5xVWNPjTFXDj3vj8Zb2dnSoibAyjkK+iXZkDK
2m+BHN+Szcrlz76B+gKBbKsCqLJDVmjNewEU9Tsxep4kBJS4XmJ4yt0uROKw3FcX
/9oTNu2XuYbO1AsSxnzpGOsUCNnIUH2fxzJADROml9AJZW+M8pXvzXBtOIpWUhBG
mNZnGcPS5tlxK+klqX0ua4m9ETdFqg1H+CVprS1jeJAuB6NsjlRFXxk4LjjThkgD
a/57wQMnytxnNkw7IGrywb2No24B0SqrYzv/FxrGeYTbFTf0q/C2tn3c8nL9eEbn
C72Fn0nQY7JrdI4JoWpWgmUkRfdj0Gqxf6B+urD8/WgcQW+Ayf3gj1Smw6hDC16q
PtTbkMugqD5rjTCIYwxD26tmr+E/Zy3kkHsg2PXk+bTtaOyvGQW7iLB+JlX9aD9u
OrccOSanUbf/zTrxNFTTK9n+YJHo86QfHmzXtcI1CMBoelVzOsCYh9KNhUU9FUQ5
si40bvyQ+er/O+3LZvqn+0t02AeenhUuvfc2X0Ufep6AQAp0Gw/x0VJ2GPNY9Cw7
fVHMI6Wn1tOFJjyR68R4CaOIn4g8Jv6Z6yQLxvDFlo+3ZrWAlcBn6ixVSggV03k7
k2IuEzdVkCL3mCTLAK1ClldiuRA9+5/gFA677uSQSSTgUA5LkhbHdB3790WEj7cD
CV4eRXKJp+fm5BxNi3vFVDPb3RFZ3uhuTxB/ipg+BUz7OGCw1N3/ISDzZTPeGSRD
c2shrty9zFWUPoDnebWnDQP6exE0mgbzIgsaENRqDdXgj03LX7Z35/64tMQAtMXM
v7NyGuuxG+6K2O6gyU4d9Oz6DQ+M399Mktd56aMX7F3uZYgeTOxpBMtO7aDHPtOJ
+eUDa5eDT1erXkPqZtGjgqFfZ5k4QwxahizaO+PKL6Tnsa4wVuIi1LYud3YqVNuL
OBrampgTgg9cFDaS3xqKDjYeLqBwC36uj4AotVc4t+X7/eisPORe09MMTtIVzAHp
DQpyQQ3Jn+ACh4WhYOzEdJf9w/uUdLg4YF0XMsIRgdKukHmAgCM40iYFIbo3JLCn
zSsfWWc+5ANC0WlDACc1UhPdG9NHxIdRG88R4p++vjrFgtqoKJGcKvjO27BRSnlA
6dKxvfJxPmYCQE9/C4C81rgrI1tF1XGoTwzs7MTwRTwmuS1Nusc296gcUi8LNnSw
p6uItLYgRKxvoQiqdbFD8Z3hM9NO8HwnzMT3mwiP6RxmlEDiUao+dnkvyQPhShYS
U5GtBgeZPtK/mZEKaFybM7izTcsVzPZX3/vfCs6Yf0gVRGsoTsPxuvzqVrX87tvK
PRrCz8gqBh9hcTd2ihZ7yiIwgamf10fGNMqXDYwasW5+9i/6/ZtNAYB9+ewaPT49
eYIPWdLjPfcawc9BxqFg33pfwGgkvvHZ8s9N7XLuI8J7UDE8UWH4bfPKNLhsHcH6
FQJz8KDNOcAr61VMF+S3CYzzBXeb+EzrLI1AN+fZoWhI/rCPyFiyyK2DqGHmdBnH
4BTVKWbRJ8Au1aOeL1iW+P+It9ipXp9dQlXyTb8wGbk+eb/Lfb8L1O5/bd7bSod1
XA1IEyN3p28UfOpu4hL5lEjbiQtFFAluDvk492FRiyaXGL9ycBB61XQpPF1EidAO
Lk1rDpDQV7rNDTAQYYq9DgopWNotgVbDClN+hQuJtt67IKYfJ8U+SydzUytYzoHp
EEmS24uT7VGSp9i36Peob2mbmy7DliBkv9RKMkXgIFzZNI+M+6CLf6atlZgJLPgV
7X4jA/tN0tpCbtycyYO8jSVZOce9SWgzvKUgJYqW+FQZ0kHtd366afrNqoeOwTE8
F1k4q6imVlyq6hW+RG4oDGPSHuqPg5S7BIgU0FRoQuI2cbRHyLlaMXRQKjFcbrcj
4FG80CG6Q5g09YMBAfimWHZXfWfXlfmQJM0PeWMX2MoOLZH0PdHX9Lo2nr5QOlEh
rg7TDzLagCG5Wuek0uizoXkDzikPvjus0hBLZHcwfidbGnoqE5JCbV4odhOWe/fO
DnwW0CyR0FpEru2fw2dtMUR9NFeC0XaS578gHmX2wl025c7ll4dS6PqOnaGEfz9D
C2IIoTy+xBM3N6RisGx+YbqFY2J0g7VEFg3lchrKndLxtQs+E7jky9LBes8oBhKE
J72FDfpMKXRKO8GCmQ3SZMnV/iEAmlkFvIcf1U02rlzYanUDWF39wQsUZpXyQnGF
6+TeWbOWzBHZXSPQg/fFH48UNrtxVgsR7whdB43KktWKTanYyqAnZ4A4ONawvwZh
NGTFn4YOeIbl7WemL1PC2T36PWGSNuRs0tcRB7927XqtiM1elzfkpl1Rcxo5WJtI
tgin6qXUt0mNlmkQBA+VLxOLHI/WHG328bjPhdhkRKBzmJC4MndZb6ubKhezulFD
yMOB8B2ciJ+xXAy7XKOKet4XlL5lN9Q2ZPZGBZUxTQ4D1R4eISl/KjSkbgQ7ubk8
KHeWQvSDN+yLxhQu+xtWPQArQiZ6D41ibWfa/aRyWCPMaPzQUr0WZB2eKse8nVJv
XA2K18M9J04ThhWVE+G4dZNEILi6hm70J8tu/yrDQEgycN1N6cXaMxZB0GFX7vEe
1gpl0ZvvVv3CHMTpX+BQxdHcmnKWGNNlsWDi8U+jFTwzA5iKMFxry+Hxxdq9E1yZ
27oQZW2dBqrJouT/sAxFcWh6nQ2+S/nCbzbrjZqnA+lsxkFEc3shyXocgNYbn8gp
Q90Ojp5EMrBlGYvfCzP9kiUbLbWJkfeC5dwVhm6uauKk/0cNtQGFpO2UDc4FXMVr
Q+MahFSkJfQEL8ri0/owvgIVx2GLewLgmVRgLssndWYrPqKcaRdqqgwOGH10FQA0
a2nd5UvDPZmW7mMxGBUefwXAAAhTzFteQ/uU3kCLT4RGrMe/9HVW/MRt/2WEhOSE
ZZbFk5kSJRH6Evzg7gHjcOOxPQ1UxYypV5GG9Vu43o85Nw5bCBVhkTv374xJ3A42
rmOueztS+xMLku6NDtQo+qnVoVB6Z5kOj8r+9+MYxhSwyHojQafK6/tRXAQLVLWt
H16MNnITSFM7vk9qUFuxNgLmPftlswJ11g48Z76A5aK4dKilbheu9l75MbjK0GT3
gYl5AeTZ0deZvub40IJEGh8RWIncFd1DyEY8uUKPTK4n6AZc3xrhYDXdVYwDkv0H
Fu9LVSq1GHRiGL32P0tRZyZALUvGNE1lpEm1HZPSlRwMfH2cHNMJYKoFLRzhkklH
kr4wKZnm7SFB4IPFNYi1xMi/cp1u8WO7r0UjBPNnZWENYqTSQJxLcz3H0TdJtPO+
bUZ0Tu3Wv4K8dJR3enHxAgZrp+XyCT6HYRBc/n2Doba8GW2io9/IGjM9f+nrWGrH
7Rp1smxucsI9J2CzlHzmqmBb1g9y2wsqauZ2PEq9nMp/Ll/NL7bbghqvdes7xxs6
J7fVlZA7dRvjeElv4XrNZoridwpwcbBugrTcuLg+A3vwDlzMlbmR5M+KZDbNDjnG
nobSD9SIkGBZ85mxCYQz7Umap1Fd6XXwupevDgF1eVgvo2PmiBi2iAqm+J9ig0hb
wE3eReykriWfDkFnpS0CBwH8u3KvgVbyLRY63JSl2UnXItIolonfY6fq7invRziA
ZN9q+WvqfjNPkmS0qBhYJWH50LI5kwWAHbrGIHX7NCYTINoanVu6sDykdFCjMIJa
dmcLlJ7xNhME/Sz5A7o5WDEbb/ipzLCGIR/kYwzNdbQvdI61VTEnHy/5hYHvXI+V
CCu/Fl/T/vbJ7uS7Y1RgX8qx6e8iaKwEcvbf2smA0RVdEbRSRzhSjav23gWgOKPQ
Ew0lkTXRAv6zxhZEGcShmQksIF2w/SvN11m4rakHTP0vGf+TJGCLfhzfGL3me8l3
6b0nHk89lhpjf4ForBeg9Pk6PlxnI6H43EIvSMRLDDud9KwPlfR1Iytwsq0xj4G4
R4iUNVt/11QyOr7quBLfXgNN1OGAbd9EHNSYwcJg/RKljC/MNcxXCnEz6kj1UB9q
DWy9SKrAFa3qU+hQhYe6nR80G1SgbWNeem/9UQrF/QvTY1C8+bGrDzwYsVgEyDZC
eMnkzxf3GuSzh8GOEPTGGTFqhKBzvSN1ZqxtSHB/PhImhhfpKTHJDK0XMuJ1Lg/I
nj8e2PobLsS5/G6w1tB+4IgBmxdYmHlcpE6Cy9aCblQSw9b013Tu3K5LQpwfABNg
6JWgeVlyPExqnLkZgHyW3dOWtP6notbhxk0zjVfWeFlRfb5jUDNPVVytNO7wFdP0
YhZNVLX1rARBX2CZWFvjf5fSIU32i4OqP1pdt7cRmsUF+ml26WCa8G8F/nKnuuac
ecE8opRJ7bwybpI8z9Q9V9mA93ZMRI5lp1wbwCTnRH3C7B4atEEanJdkN60i8nlK
JdIhNECS8jLaXfsdzIr+VUg7tG4Ky3P6AMsw8m/5xgqhCP1H95eBMXc3nomaPPnI
v+F+VZgHa567+7ZuK+NrH3AZYPR7NFv+JbQOZYQlLHKdnrOdqFAONlWD/IjSLBHq
R8beJSaW038EA2oohidIU7X6w+yMC0p+MmaKBtx9bqCPPWFj30biHqPpmXlgZyGQ
VqZ9Ked29GG9LLMTHP44EjTJIR3C3mL7YPYts5nf/Q5qsT/jtvfCnoIyaGMIOShm
UQIZuD1Uajz4ZiG9S4QPZQtcZESCRKZ6HAhx6Nr8VBEXE8vBvpzlxqdECA3X3d7O
vJbsBOvaPRlXh1Gt9Gq9XcvMqG8BKs9+//SkXj8smFls5uDQw735loHUKpiNbCRM
86Xnh/x8+EFrc/YXuAIRlpwN/FXHWFExVUM9lVwosvnBriK2r22v9cETnbZhq5/i
yTWFAqpq72XRWsa72w3RxUAjvnCRgwOnc27NII/bLUCFBcWN8eY2/dxTjK7MPUvk
tMw6fgI0MQe/ChC6gHAwtQVPqa2Uhq7wpJKFCpPyhMFE/Qe0dptIp8YI8sdvy0t1
PZ4lxbzXjg+YefiKIKZkCmxBhk3PYzT/u+J9i2Dy6JN60nUPuq3GvqI/iWVXK27Q
FndvgGxf9BhoRO6dhxVK+pu/JQrHNr7rihWluQsUJxbPlp7uONCk1Q795YV7R350
DYWg0F4MZoXg3hCL/5/11pl57wdq3Xtk+ayrUqvFGDDHKG5jVG+SdtC+LEiUyPQP
n4k6xOPuCCTcaF7H/LtOLuPsNoYbYidb8OxzEKn0OO1zCEBCqJtKGQB+2E9z46O8
ZcmsYv2Y4ire/+Z1OiL1x5ZLAr1YsTPPQh0vT+XgnoI6txUTGa3/F0PLKlKWZtv0
+mRCEEfm0rxvVLMJwO0R4qsA+p41hYb1VIrAp9sFmQfmQNixP6oeEy3Lqs+x80Qy
Wg8Q8G+VvHEj+ySUhfWaU4dX5V/1JmOqRJ9v5AewGXS1Nn5XMXq6nIx/HsJisRiI
4Jikw1YOQQfHDmws9GKKejNC3DBEHRpqXczSqZGGnIQ3yYsYmZ2wzs5WY09Ap4tR
8ooftDlNYl/qcjCy39Iw1yXdSkcdvOl0kZvytC6rChvNq1wkiYV6yhkGEahrXLWC
kONo8UCSG83JBmxdfqtDdaHKsbhB/nXAT2aSUmojajTUqaIMiochPZ4M7oU7f95a
WmM4i+LIp8KSREVoXtuJhXTIcZS/8DfCPglydgDTacW3PmZlJRjMzojSb/GMFqjH
9PF3VnCMu+fMOCVxck4lUloWLHWaqUjhJm2TcAey514UJGL0wujUG4OpX9hJloXQ
eUfOvt+HQgvcyNKumnSMvYJcNWW27vkACKBc5pC5Ku7D9QOTsQ1ikJ9jpQo07dlm
zQ8JmKhE69HjfnXgX2GPk/zGp/oRy4U5LUBWvPvRiApq/+A3sopHrpUmVh//gQoC
FW0YrXPE2xlK6KhGMhR6zDCZ7PcWirz3tXQghsZdveZVwHBXUnIdFRf+j6vQFDMr
+3x6TP9nmdsvLmRMr9Au5YoNQp6ZI5E/Q+hE8yEBCLQmQCYUCLT+mn5WI7NqHEr0
GC2xhiLlSqVsqMT7HvoYiKuYbtd0XLFLJN00InpGl7RA8jQ3uAg8KZYvGvmK6iUV
cLD3dB1TSSMTXnhCHN1cRwzaYokCc2GldHfxnVGVwEmi+IuqEu/NqtDhYv8hl4VR
sDdmlvcX690iArFg02LgGjR/B0Dr2weCxy/9k3aQy5MWk85+TwwsxUBzk186kLXF
CUNo4iTD8me/r/oTUfSOqAlL8hac6WIMA9W08uy8JTQqaO3ERjhrM/4J0dqttkSd
TX4tWtp9uDgh9hTGIa19axI3TstN224GE4/AybW001zErGBo41BvhRdNfOJcm4o8
vSfP5aTEkwm6kGV5SPMAJk60n34zFNAKFmF1oO9iIHF2iu3ywg7TitRbP6igYE7Q
s2NK1vCOOdx2IMCqK5Tfi3YA6k5u7Ko5HU4K6iwPE7g1T6OB0awPxc4H0WrOwjCl
Un/X2fGiZVdc1bIZ5okd8Kjx8KLUcmko6NiF+eyprrp+qDsgxD3UTLpdXKsjm+1W
/E/cfBRbtb3EhBprwpUolAg8vBvEHvHfudVdxib9zNWfzptS/hW6gl5Z4ktFKVED
Dv/Bn+Rgxecua8oDcfnRSLAE/6pivjt2l5B8HKujtFXw9rnyULX3GUOPwrWAU0AZ
wfZGFXFlDxfSdcVzJyz7qnS4p9AhCJyCuX/KUDcXCeQDzTSzQMIwFaKmChehkTGx
JwuT/WmXxrBKcJXaZXWJ+LRJR6t1xMZFAgWWiIUL2Lxq0/UzT8N/wmi1jZonGNgL
KVoh4KxX8uq2g9kGL5Rtu2Gu60vTLrEKgceFj4Ikkedd3BcWC2dnpveuKz+0YEYM
EsBllxXV9cu2SMFhPj/ZXC74yxe2HDLK35+r4/TSoG5adDxtwbrgF9b/yy9n8hlq
jHjDW1+VSaqleR3uEcPrNS6P7zhA6KJdzZX/3zz+PWiOlWY3pxdqz25Zmdu9hBb6
1ujufQ7ITFylgQP+ujTFXpeiFUCWFFG7L4YnA89RVSh3sMGn7zOyyfD6zcyyCb+m
27qwPa3hyN5TOlu59ybtQrNGPfJ9w/YreT0P0koCi2LIKdPlQmL8796297d2Xpgp
LzQJ7gdIxR+e10EV+aoC/j+a9iIiLoAxA6X/Zj/K9xI++XDuEG4k5LInOhAvTozJ
uy8dAQSNqg+cCjOnitFiGrRKPrtDMPSwaaPECDnNRO/fepJdFtCOOxVTT55OZ2ca
xSw9pGAXLftVoBUX4qm1hhMLTasSJrHZ4o3SGlTgzi+NEvQomwgcmNKNj4Oc1lkB
Pbm3DfqT/qcinYIPYV4eYeC216FELdbF2msGezWUpNb84fCZ5hyMAN5KB4n6+CHU
j7JjGMgZ9O9MDvrXYqnvupjrI/UF3KpU1S8yD808xPZb5kUuFxowjr8ZyDBq/Sx3
B1Zuxklk/kJkkmY6o7en/7kOfR4vem5pq8LeJBztK2N0fwsN3w5U+Oke0imriP/C
g6MDqTBavEFfBjpaJwhX2m/P8kIB5g7qDIYwRtcBWE5Ig2MsgC9/6xBC6VVQe8Yr
J1rAlRVwQd+GnOwRSuL7449HW5rzyR4cHMruNVlJRfJ43crCCD5b2ay10yWd6dlY
84FQK8hnPSbSfmQ0zSYKmTZJsVyw6tQo/lb+v5heHBefr76L8PLMNGkF0ZtWbnJN
K2+iGGDQiDwpmPO+2O3/JLlhm8NM0aBnNjzmO/AwVg20S1kveFp5AySjQvShMg49
CFpBvvFdmObWBxGO63OY/ynhvtd2EvPKZzs/Z062UGBglJIpDezFgiFirZBdpbS5
F26/Bvl5rFg1+s01xh9dq8BOQbksytJrWEehee+e+CnotU/EIr0aKo4u2GwZeacs
gkzXDpux8eBkc2J8SnyH+Gg2VFkBpeYkW970nJABt9PIOq3hixUlniTLdH76VVIl
S/g0/+eUOD8wLZCyd0OgiH36rvZ45z3DYZSqn4v2DoOOFYaevLCwtVrXo4XGgpD4
xKte4OSODd/CBW68/koIudwqxRe9Pi6z+I+BxImlAg3+HyMbBP82LumD+N+PboTO
EfJYpIFu/wfKdSmdj3kZs9iMwuEzoqihxQE0So3kTHvR1GUq+gBfoCVLoCSyfX31
TNstvfpy6fAp9Sd3VrFO12lNcZfv4zZKmmdjm5wx1m06MkO4JrgM9qMx8Di1o/uI
yciaD6uOSUBl0gP2KatXsVSnrS8G7kVkQnWuMWsbYkXfw9QjnGMDo/vwhoyHIfBV
DpIYR7QLq1VoFuMGs6chV69ZnaoaWrvxEpiHhGyOkZxO86GR+Evz8qxzJmCJ6v0V
m19nlnUd7bdcufRAsEyQVfo2BY6bE11ceBE64kvySWe3DTYUi9wJHSay39lTe1rY
ylxvt9AjKys9UyMg1N8j4heQ3GPSKmaJqvNYB7CeTIX1Tg3Ec8J9ZjvjLHVJyZyg
LEBLxietLV+yGizt4vBF//laMsBz6vzQe8kAWkMLSjB6EhvblRwhDeeKUBVHRZaC
MbpdumYBnX7zFGHSlYxiHbbEf4djejbOUdocOePGfQPftlsZkrgptokO1VS5oqZt
27TcQj+JDYo/a1mz6XFl9yY6OlJyN67MMETkDVHY3Mi9nmpSOcX5lxwTqlCiWtGD
U5A9VWvzAB546MJWpCvETs31IgkS7iaf3Moyv2OSc7dLtRzSi+T+bZ5xKItjhuTq
Rn0fucZ7/SZmKjCo9pezfVEnRplyLF9EtMkv1nHhd8Hzra1eu/huUnlEiLm56Muf
rzHtwmZIOG4R8upOJ5LJKAYJQovC49awL6IpJP7ZYjutcDe0bCRnh7FMfJGTLZrb
0Y3HA7F0FtS4CtiI89RW/0lnw4iYTLG38CojA2jIMDfXfHXKHdPCsat/eFYcnJYF
/7Lua+CuscgX+v/9NEvqji0GpNDrwM90cMSiKWv4J+Oo1tXYX3h4QWwrX6Z/kSvm
vjIEPOm4IeG98l6lilKJoxtCbt1Ex67dK7dPTFQB43Goo/th0tLdUrSHmmRKJHLK
ybpVqQRwdLt080GrKFyUy6qoA3mpA/aCB9/pCyviI1vyGTJVNOzN+5NzkffPVlAx
THv4gXmEXP3VqEhM0QHFVMuAJ73gHKCnguv1t3mkNVjB866+w6iVim90RKvrqZ0e
a3r1kxu33I1pbmw/RR0tOkg+8PY7g7zNjKdAEvZ0ihyOlrxVjtqETkn/T8jJnvrY
omxx5Cd10n3fMme8K6zJGuIB84tHh8U5MI4PBNGiwlII2qcbpIQoSb5yk4ekR2sq
YZfFY5VC99e7s9pXjy9HPYLk5r/OfPWfMjsZDfcl5t+wcX5sCKgbpmatEIM1OM6j
hQS22vlQ1iWmyW1+zcoUUqHgFq6ks6uk9Zx3FVO77kPxsbIVWfcASKkFyLY/hgdm
S71AdjrDV3C5hQKLj2i+X+RxfajW29+8N72I7TPa5kikRUkX6cVW/1H3KauI0dQa
dnFk7F97+o5/kVdOfre1Nwj4vyCOkhdUY9At6z85XiqLiehYaHoZVzNoxJcNTkIs
lcUY5CIqMKEuvZCi4+Ky+NbOoedahKVF8JK+fPwGDmNeuBFfnXObjgZJ7m1GeEZn
/29/qFGKJCLe6i/6Qi3SdQJEFwVVPemPYhHMEzK89hlNPAo5Xl3wePI+eIeSFBiV
WC0Qb8qHa6RysdDEZ9pLCjca1/53f90Op02AphvdT+IfCMnVn3djhI3FMvjDm02p
dK4JW7DPO5xW9AQ2m1twHBDf3DwYw85XLcpLEJIbf/QNx/PnBBEDtDaVso90BtA1
dQl//XgMLvsmEboP4YYhpiVtsTINXi3p0t7td4WXhUwYWJHKWySoaIUHh8S/oOdm
DhGvwgygbLMvn+WOBkHgC5y8APjg/waaC5PLYLGD5Io2CHXHh+IDC9YcmKwL4KlZ
HuURQmjcbMOj4Dwi+g/Cs+b4y4clqSaqzAHPDGPIwRKm4Pxnnok5drOONEx91dx9
OcSd0mhkOCXIHlkaLbk6arYTj6SmNdjUKP/ODiDQWZqLZ8lJDv8lHIRXKa68abBz
XRCzLXLWg6hB4zVpu/vnQklum2Jz9D9MRyvhZuyL4TXHamjwLTvayJ8s8OS6ZUJn
haPOWzd/3HdPfMuTpCr6st6WEwfHC7L33TbwLTYH1VbslDmWmE0MabFy9mLCweg7
99P87ng6z4YQvlX/hAl8LkMmYfBOGeXsYhvHi+FOyO+evJl/g/BQCX5iGlFq4+FY
dpVpmFj37PjCtji41nw1TrHxtGFTvNXSpX0gR6MFAkvocYxIaRGwUjt1Dq66kJpl
RXCuufjrAqSkbzR3+1v5LTPiEuAGuC39AOuMX7WjfxvmC8WGUiQb190BGxFDU6Py
dI7AICS2bUrq7pwnpDA2Vb5bc6a9wJMKxiXQxkUvjbMKgz0va3DDhcDgEiwjVo1+
La490WuBAVeDHIye6nVqvdpgMTgPe6T3M9WZs+TJrYdWh1gMjP05pAwkDH6emiMB
JkG7zmEGvMf9MQ+u1wog6Qf9XY5sCkRU2YZP4Q9k8le9m80pzJSoAeSsu4V2GxQe
ISdHrRkoCr2bvUP9mKIuqr0E1d3ZxdHTgAXy6FAFkVFKo3R1YQY4SIQ/rRjCs6VH
DrRdxLqusmz1riDcJv08X86FjzLEs6/qV/E4xK+07rtyAA3vwgg+0mopqC2lhtnp
+yvAWpgLZ53IPqGxyvWfPNVCvpoGQe01hsw3w5qiJ4M8mBG+JEe2im6tibwXr5KX
9usUt+WyDZl6Fllnps2UTXB8qrIBzyp+O1DtmhVqe3y83epggO0Rr7la04oQ+0D/
98cYkuX5rN0bkK2jH7PV6XbSIERDdxtwh2Of+yCSTyyoYf9vlEJIp9nQE1PWq1b6
7o9lpOI0dWFmGrLHOlEiLLzh9gcLL5AobhjJLisKc8MXO4BXW+eUNez3N9OJvMVc
A7JP1+fpXiWyjmLkUm3wZn20yPIH2JdJFFwX7f3vLIJvgotCrr4XFhiSGoO20Won
yUELSQd2aqp8fleRf1LdR76z8w+DtbcocnRgQ7iqQLZVv5DJo1v6NboiTrhpJkqH
454bYDfhewxrl2MmQJzW7POEWrdPDIxHA/RrWSveJLiW2O5yw3c3FtHIRZdbYKBP
4QjWWEsw3jvZ/A7R3Fp39UBBkHomd3MI2V6wUcYtFIgu8P/DFr1nAhVsGX3M3+yz
WdALpMWNlyqpN5ZQDFgPlLr1wvlXfZ8HPHe9zeEAmhk5KBa2GjsaEHar+TN/jB1K
Avsr55FMD4n54jj9sWQxIsJAGJA9IzL4vQMFEQSylgrHJxr9lOD45p0kD1qnnz5G
8Oa69pkFURhm8QEbMh8Sc09fvkMWjOHitBINd1F6nvCQoInwZdthD3m/viH3d5RN
/L1J3BPimexJrWZL5nHVljdP0WZ1bpca2E+D6gtse37+QEf4hRlQju7qz5SBcMpv
KaJ5noR775IMee2CHO4or55DfM7rzaXHq0olTSzcPDxcxT3BsN8fHK5MUJMACIge
fDq4FXCc5Qgifnu7ootTvjskkG/lQ/wp8w5D0KnEFrAjjIDtL15ARczqtHtILo5U
zjl7OP6iDTkfVufAw5SAWv5VrEQKcU4pvVv0i4iiHGlXZQIQlHQANmFYGCyuyUVd
WjgCiob8QsmsrTr4OaJATOsBwxxdbp5WW51hJz9kwQeHqNgydxJ00APg7+Sx0DgS
iip/qw5OiGy6Lyjoc2m3cRccowqPzfmcdDELlTiHbJNXWqz265/L9zdLb9dAnEe8
IA6DP5Yi5qRwgmqW3csSMeMLn8t4bCV4WhkNkOrzvFVoMhWnvuAbP1HMCNSCD0ah
vyeLq4axdjnPxVh6x8jbWj1/9R6oG7KNlAAaT3V+EuaJZXlfQsZ0qbqww3pMwSx3
QbZ86HaWeqDsTkeyjCS2nDHCyK1zXz+5o0fJkI0zf8TCOfOcLB7fROzD6c8krrQy
bZ8T5bpL4od6R9MIkide93p3IdcCRBJoUteUQMYbDwlAfFATdv82f8zem1mstmzE
fp5Nt7uliZlL4h1P8EhMEFaMRbL4oRSD+XoxWLoEE97lzLa8S78M1LVnd5M3BUBM
plVXKpbs2FOaiXg9NgcryFJtiHz2d5dLG5vEpRTE7K2beNGVsKEygCMxGzYWI0XW
dbwft2tibhimoJq85NmTN2ho+6Hl9lhf4aRjPvEyg4aDkg+xx4DbBwRl+4z4CACk
WuqOiaDc1yIS6gFkJ29aamGthmmpEtlh2oCbcppEl6ADhWpWBnn2NbI7m3B0t1fJ
wEoSbC2CZqumYUVDt8Z4Kr1ZRAgKlVEGOtpuUCksPVJSH9lmoanmoE5VXlkjIRak
9ZjCHh7yaHI6enbZ/KiysgxYv5jwc2OjsPoS9jr4EhxRqq2y2S7oehSU8cR8RVtw
GMEFUrdbeyiow0RxFc8gaOgIJS3p+K5MrrR6WiMffe4tGCLeTev7RgJ0H3bwugek
AKU4rIZpzwRqeq8IUAZAefKr64Q8bfZJuJjt1cnhIHefc0w/CM/ywVn2LT96tBfT
seAPho91sRYNaqVxB0+p7o/PUjAmxCfUTd1Qg1VGriVGDdQeH+6Oo0Emf2Pq+Wpr
GUNDbOd9AlLY31OvLyiJP6ZGumN0G4OA8TuNeGvRrrjKZNVo6MQSUSo6y9naSQdd
lDePh8L6Pls0mT7LaOguwlmJuxCSTPi4tSkFQiAGbtoU8HAnIWvGfCp7IXsN8b14
+Xyjo/IUE+FtdmqH3Ny8WWGnU6up6HmEKYwgK2Ah/DvWrehhslv3Y8YSYgdjZpcu
6aAtEbI2oL7YVLl2KJJ+V4tYXFmwX4+5/6/izpfPMjW6SG9NZq9rbRwAeJevrMyt
/bYtQEtksrLt6RCTtZ/ho1BgEOUqZXgkqmKRYFbNoeV+ThHlcibCvF/PAyAG9ikE
sBI2+PPOQ91gFMbTCj54GV2lhucNUDMgRjBY+dKh9FelnXbY8WdE588mAq3Zg6LZ
HsIFiGsWoP+UeWFEkCqhYIqrAm9ngeVILsOkFSMWVWiL9er0GHoHzwokPg0Zsisl
XFLkp+lgRD6EXjEYq+H6J/TeFeuDveIJ29/CGzK8ow9l16Z5hjWc8fg2x2JHRsO/
QQUd3Y7N6NMTXnvqVAApanOq7v8RuLwmJK2mp/9kCdEp0PKDbG3XWgbYcxPa+W6T
2vqLA0UB4W8LfWuhcw+KuaLVi1BfupqfwOEoCDZZXo3eBccOhCWJdRy6JFsLREnW
v2YSPuHKYDsvd/SUEAbZ2K3gWD7yxbY8rHJcR2guuTFuwMaXfatU3MivaOPaXZVG
jdK6a/KPeGTUYzU14Nvwt1r5ZtrKjk0reyWukUHMO8wtYWGVNLwP+H+Xb2LnHmuX
s+JHUDUgEt6S/rh4YArp43o4HwHjpmkWWZwm2fE4Qj8+7PrKUeycSdpxNtP/Gm50
cJnlW1JueaVTz9YeMfyrprqThEiVdXlTEsLnUh2WIuIuqtK66HY6hxEGcAxeloYD
RF9O62lquUksY49lYanPmfLWlrC/WCMhMHbTozwUxOyzuBLfwgLizWxKvCmIsQzz
CDpitatKjAa2JWq7GztZXzHRwqeAUoUqYu/0L+qIDNqc8bcXzvibGX3X+jCcbkQ+
EMvFn6CYTarz/BUyfYHAx9GCiS2WeZmQhnGzQUBTJaD+OpCBzaj5QkaaopXXB12s
BmLCv9LibEmqGDoTEzJedHiuwGP4lA5zNlzlxK+t7kxeN7Kb6uJX+8CdnOIfKL7g
PioOy9pQd92vqXCsxLeCbDFyGiiqSe149smcZfdElpKGwxj9MQiTXTk/5Kdjl7Au
u8wbFlLv3nFSv9LNgmHVO/NHyqpcQ1pPvsoQ2pwhihohQbufT4HYPTTWKNaKlH9N
YDG9/LR+nrjANKTVdO19+tHZac7PmqTVG2DSNLIrx39mj34jztA62KPQpYn0nfBz
3nsLsw5k8aQRZ0lNeW9zuGt4XRGzHI/rggthhsgA5+c8zevMX/W8ncKUnKOd103e
EEb99sv+PKN5rnY08wQeH5JeBYBybjP+1bSyqeitYStVt0kTm4rF2tUm0QqRuU7f
ztTWFSDuhiNw/qzz+7tRnEdqQwLRapE5aTSYrvf6WBp/BcKEHkjgYGqC+FeU6Bxh
YQViuFPJxqAGVCk7byrSU5xLLkQwwmHVCl40ngxOX658nubWiPBSEnU/+cgoLTFp
6SHQnQW1O3aq1Hc5kHm2Bbvw94czoR/kINr7t0seajiGC0zD4Qelvo2A618GO8BA
Thk2+Toq6FE0yzNfQSMMZW8zCy+zwsX0WvBpQe0+FUnCL4UwjyrGmKcm8AT5wZdW
snqLPdBwvvJP/DQVITAin6Ku/tKOjKyRJaUbONN7iQH1iXl7nTOrVGhaFGEMwGGH
V+wuZC02jsFqZlnEeoCxNXcOZ0kPSpuIrhU1Y3EvxBEkRcgXp24iI9vLbRR7TuDl
G7LqRssoKSOi0ikPVXwPIglS/bI9Ce1Ryeq2snChmFq94dnytkQDxO6t7/9tEYIH
A0Dw+9FvzczidYRGTJlhE5Tax3eztIneb9Vqr4U87lae+kMo5t1UVXaJB+YWNJE9
Fk6MBPD/uyuQSTzPnINcyzzBo1UzwXr+YnVL+Qq2Z5BqJpUjipo3pJJgcjhF7MTV
SxUW20S+XmDw11sHuo46OyZmpbBc6ScSQskppEMXppD4wOc7HQvtQzpyaSkvtM+C
0753zGpI0TJyGOptiVh3vItN05vjYNoamT+6BtZdQJk92p+sCkApUs2xmDnfMwYn
c8HNoaZzXIMiBe+ucq4mrBr3HW7NF1M1RMkDayEKBsUQDRbk3mDXLyyfirJwFV86
XQUeV6XGUVUzdZQmAr9884+KD62rnfwlvmk7uohGT0DXl5/lBXSuSPvGsAsxJQP9
GGjduFIzWKvxQvLCTkIcFrHMTsjukKccVYdcKmVF+33QfjDaQph9P5kEMCjyX99g
JlOse7maS9Ev0ZUoLYSACF1s1BXvilu+R20/k6EV8m+sTjpBS8tPqyRU2t74dvGf
ykbWjQf7fP0dsWd+MvUZYUsaPnwfXkz1GXeQk2mbBZeVshkLDSxlOWJAjFWOooV6
zjw8r3oKfs3++eqIJGNjT4zWx5n1o+jDbap/xLWYiKgkV4rDEPRvFDjiG/DU17Jw
pAHFpqwYnlKn3VNG/jcmHA8hYQr3EUXkC2lJPM8is/aEMKQSypuEhpbyn0Mu4SHP
BE2xYPkuN/0vFEq+CASwnXuNdkfAY2qr5sj/M8gnnyLvZPOrpNKLT9ksgD2Ejr8Z
uOrwCSOZNw5H206pJLf/m/tYqqSbDj9Yh/kbLVfRdZ/TGjWXEbfpaq6iawwqQHLU
OSuYZ6K2p5YBQmLkLnceWcJq3Odao5Wm3e7JuBgxZL/Evo0ERoVTdyOuxcTrYA9K
tzT+KqRVaty5swD752FMzhnqy+vfQs2lLloBPs7cPnkdHkBVXhdjuDgc+hcKPKCd
4qFOY1pjWAPIRVhyBTxALLBw6A5BlLEtJzTEIRjLzgm32Gg0Ap3Zv4CARhqk+7MW
J3sjuyPgQtsy55PQZLGWqYzmL22WKy86wpeyG17glntvEbn4FjWqC8haJn7a/ZxC
4UivoWWuNdRefihBO5X+iuO98C1aQgc6PkIQ/AUceoVk9u40hEyXwj4d7ECUSI79
eTAOsmazk96fI7Sml+f5CmwccEST5zGxRfi+dnmkD2TQN30r2XubvVcA0d0GdkdH
wMkKam8REyxfu8sOIPp0m5r6jTvo+wwmZdlmoeXevOjyyUh4UIfIqYvKCr1kpo4l
yEYrbFDMSwBA+8SHxo1i2JKNJL2zBKrdJQIJK3vMhKHn7yBV2GnVjcOxKqIa1q1e
azjPhdGirIpiwQSqRcOlwCrordROrS0IJHwWCq0H8f87RyV6V/IIWjobzcWO5RB8
A0pO7ZaHXJFFnvBkX/MzmAgj6RQ1hdixPdU3SdrPuL4u1jzwbOXMvAdqOHUZKFBK
PkRnz+2RlxRH3gPBHd50aGN4TCLuXqWdqCCQ9rKEYAuiAWed3nZblFGZ5/sKxxKK
1EnTc0kF0agfsdhw861phTA9vyIfbRVc0RCjfs76kNsLBaB4qGOCfoJobs1iNxzj
i/RFv8E5VKvC7s4gPV/0Z1Ctxn3vb8SDuXYHFgPlOnNJJ3lDf2FaE9IiN1B4xNZY
JYepT78+sNgcc6c1LK+7WKeQES+8JN7y+dFqmlMiPTn69NLNLGsZSkoTF/m8Mpth
nUvF06fXPCsrZ0t9UQPY6AYw4mk6SZ74wFfJ1y8Fin3LOGq8N/AcHGUJSBvThRNs
r6RxChrEALJje4LV4jTwwKwPv/13EJO03qjtf3I6gIB/UYJNFhoeX6vOVplidLXu
RSpbewAjbWyV1ELDlA8ER9wfETkNQJQzY486l+xGEA1K39HEExku8zWBkp80F/Ih
8qdBD4iM1hpGblbz3Yi8sXLOX/Hce5Ew32l1E4PF1VBLlugaXm72RNf1rUSmVPhg
BKjzVIdT+6G5qPingGSFLdWyaDsV++lPuE0O2UcKsu9bHbfosSlUdu9vwF46JfgZ
OjbGZ03wgLYuZpMeoBib3z0T0yILNyBWLtPZZPTJZTKfLoxIOUo6enalSCsAY47A
WZQ2oFygzzoHeXCSsvyyrcmi9HU9IbFN6FpuWEnqZJD8QdxpKOBgsy7QrGg+rg2T
EXZ/FXAYZ9r1CvyUj4D2w317ibcXzvEIDooUKII+AC7mI8+Qt6H0jCYoTidkem2x
KZLZMw4HrZ6o8mB25/YFFC2bDKpxyJxNykGbeTt478i6/Tbyz3gwbHcFW7AjVuKA
M9CiY91wXOnfVG8Tq7btD9InP60NEwjp/2KqFvKnxbRTPwlb35DEh2vqbKtbq16f
xbp8RO+HwtcfwBBuFtsOmlLA4C1T+3FZZFlNNHr/BsSe6CpL3hqcXqjCguVfiKNE
TPtHPmJiq17XG+qKZbi+UjBs6ztkgfXxhNcnwUb9gDLBoeW/cvhzeBvNIMR66hkh
sJjrAZRfF+HgBL57deFJQ/i/jAaYnudmkGSgq/g3K8xPH6mRk2rHXXzt/IL9pien
fIyCpoXlPEYrFHuBr7p1CUkVr6yWveWMz/pHgloJRRgMEGf6/PuFzdFUX9TyJ8PJ
sEVzhpUsq0EwK7fL0bNvYtq1SjnkctYmhj5Qm7XzwJspCYGRqGxO1kg1okA1iUvI
4rvTT1hj7Z4ZqAyYd3RsdDZWWAIAwwag3TE/1GanNq9pLMOmiHwtTG1qtyzAMr/4
/wkhu6bn4/or0mIiTCR9uSnmmDHAxc+3gG7YBRZJjKU0tIKgsRjRJXtWmyN55VW5
HwbAXSqDjmcEGf85+F7LUuWJDG1L0H8bfgmBTrgE80COEWwgCiJxWsz7UukGDMIH
Puu4Wz8HgNEt0LIZ9wbLIO1Ij5Rg8e5KmhUX+IGwME1HgufIPXr/C5N0D5aYaWMR
A4cCWpTRTeGKWmIL/1bjk12k6HnXfSPN1LJet6BlofAZycV8TjRlBxrUuyakK6u9
ujgapCrau38gGjcIpryuU+338HuSEW3FRzeJI2taSYguEDw6nJFxYLoyYGsVlW50
FfB3eIQdfCsMdifJWjtRaYjqidgfKIFVZHiLiViIl++GwFqAMyCZK/b46SKZNV39
C6V22icwsZttr6fcqA+MUtgXbOc7LHiS1w3oWdT/7tjNWc4zy/N0QSMxiCOtsUig
xYJwb7QfoDODldRCDZ2W0swfKsHYO4ptpnZ3BMxHx7cjd8zHUe46QBn9AaE1D1oh
Af/njdp36vne3GB99jyUf9Lv6zHeMgGgt6QgN+5eZkTHpbSeb/sGwZPLw/LTnp7B
hLTZOytz2PLRuDtj00h13sNX/S9TPe6qMFhd+ilIit4AMqrXnxKWOjz29pbAtpSx
FH+vnq+9qafL8DBVoI0h+CkhiLTWZiS38ThVgIqgznV3wdEPfoi0438C64Z8ZpU/
ualxORlzwMae6bhjNumrCKyFspaJSCnviUQGNWOxM9qaWcLhdBPILXZyq3/K+j5X
Qq0zN0TFQmz9+KiwjWQxlwkpwc8PFBUiNu3vyZQofpWG/O+GC1oBW8mFyohoMKOC
X4B5oS7GXg17PL1p6gxVmktYFxtnu7SzmifcwSDrub93VAB0mphb5EK1KguVERVO
5AJX/7hOJHKNb4C4jgojOtABckHmVhOdHLq64/TP4TnvU8MepYAUxbvO1PfH44fj
BO9z3X6Aq+VgaWak8fGYcrj8dqLxotlxlFCpIELBSTpfe8nVdTLMOaVq3GWr5B8X
MLGB2v+r9eUksyH4x2r0VfN90SYJznA3LbP5k79U1dm9D4xt3VVzrPfM2lKH2/d0
iwRrSYImC2t7w0gCeVN2UuGpLIQ7muB3Mly7w4bohGcgRePdjsD5AZHSMlVap+va
B+9BnM9FAQSOWB/78QIrdvVKDunT1lUBjaRwasLj/56h75hbPfMkRBy8lbsU4i7y
0UGDfVHK8Q/N8MELAgOo0mWcXUMZY24DmCo8qbeq+7qigLxlIXyaBxg/MN/nUVnb
7jh3ZF08m/xdorU41mIxlPAzzoRTYFqfihtsq3Qy9lyVaTa2dFmRALtFjh+g8uHU
JPmaVcmzfJzokDnRyr3QmCITu3YWkv3wtGen8H3Zp6Wj+s7yktBHMiCbLNS1UNNg
OgekBHFag5ONQUAGxbEk/N3XUwpGoaolupZ4wfc0hMuQrRAMUmYRTQJcZycDNcEA
2f4fuLk1rvQWZoTCqpfVWkoRIeQq7267an4gmB7TxPe7hg9WkMxQvK7LXd/ZQ9mW
sdnq8reKgV+7MsFd4+7isShQ9EshG5FoBpldv0dlAT8NzF+khWtx9wk3MGjH3Omg
QGhLRIh5l1vvT2lUGLXLQC2vvU6e7DsDrhZY0i/caoBfwlJ1njM2/aUnC/nolfJx
Q1AxNDOGLCLyCI7bOybr05XbK5bKRAJO9z0U8OZ8fOraCOMi+T9V01bcjab7iCJC
d6iCfhHrMsBsYe9Ge1cUk0fq/7NldyVL13E2+91qFvRYhLyJZDgFBc1T/Q7QCdsX
RXdFsf5AKUTDPUZccy9EejwB5zwalWqxZjxhMo5ujTDL/LxyznhRODTTbXO0/NoQ
ijTRc+tCAGG3n9dppgUD23E4bhdgq2Cc7FGh1ndm3W4he2hmsCrRc2zBipy3+Q7b
tJusTSYgESXL4GaLrAF09Fc2X/vyiPxfnLdI/DglfF5Ac09hQ3lz6STCXOqqz1du
u1utgbTyoeu2bLN9VNloqGhQg0FSeYpQZfZKvK6ws4G5J2JH9yuDq0x2aoY+UokA
gh9tL+8fPg7Dyju8RfdghHwUb4GqK1O6vM3S3JXa040xq/j9HlrQETli9QGWojNF
SbhOcfTgK0eJjxruAIV3/qVmIkDHCMdD+9sZhQQc4SFxIV2trgvmz+QFlzCW41xW
/5ANRDZWPaOzdAJoyszESbY4ba7MDbxvffGBql75ZGXA6VEWeh3QnYXsUTM6E3hk
XGy4iheec1fFFXaUp+VoA++DPWMp/7IjOn59rtMYiDuLSxZnlGdcl3r6bF/QZZHy
hUumFTlKfXMEX6TUF4eSzFXgFQKJZBYnHAd1Ky8ywLJDhmOOJ/rohD8xhVuu50Wd
Lil+wT2ww3/yhA35E6ZwSLS82T6I07bW/dbpBMg+XcrwHYQR3R/oxEFeIB/0q/W8
0CZMruTIwjqtP1imownCwOpAX0xUX97gYDQIHOy7dwbE0Pltn7a/okg4usPi9uCG
Zfmpm2EYs6xHtwLQ6RczLIK+6wFx6w4m4KqfsIQuA4pMGS89vKHJvmmDvR9wtui3
ZYvONXEUiFNxAFFbtLIgEmKukPs+OEvsKyaJk9s7JxgaVZYTUg1Kj7Jbu52uu6rc
/Tj3NI0yixS8oGXgOTDW1U8jYALHlssiHLAq3J56HQG4orMY7cyrp7cBTtvzyB8H
2JCUA0Gu2/dsOzPdtwVKZAeXX2NhruMsfzIUkehVo2GNcupRUCe1qy5Arp58gy59
OGp2e2EenqBnOuNpjqlrZBF0EMWygleOtRTrm0WDI459EDJPG+yfOK1ipya4BZRv
QNZYO+tB3sXdsOh7PqMEEFvslfTq5KItl5Ip9vcNy3l2TDl8L1vYdXqGltSL+DNA
m8r24KaWuRTvlRAkHRsT2rKhPIKe6X2StXDb2g3C5Qq3ui3T6yTBpgpQi7eyfqLn
LZpQRkwRiUzbff/oFe86A2qMexO4V/0lAEblXR2uUvJvCJxD0Khj90fQHA6pyi9r
hEj8jm7YR5JajAky0RauJ7ULan9sYveJ9Lg4kqtTlTwblhQxtBBV0xZHWSzo1s5F
ZIx2UymJ72T5t6qasXon404tRXOeGviVTyvdg54fp7+OPnBDcrGSCli2KzC3wW0a
ht7IMjBbvxGxG4K3eZXR6woRExTE2jxiWU8F6axHuwXt/bsDx9yu2BqmlyCXjVph
jDiTqT5e2NZR4pLEx2OfTEBCGqFxk+9iG37wnlxmWzyCnucyd6v2a2xOVSQAe9VP
LAcE30wIWrPlJUcQTIiTr3H3yZwSf5QUJwTmsEKSTyEt2mw1JO+6eNf/GpN779sO
/pMyddY50VDQOZM6mP1SEmcp6f/vALRK/4+5mZp4cpdB1588rlFYXH3H+FaGHVEQ
8amwbMFFeuRlmMyuuCiFZsFGeWDy1qd9UvYYvqDDAm1DAvCFR8BN9bDdtljmOIHD
49IBL/GgUbXF41ljjQlPezMtDFQsHsp19NjfxsgpcE+y1sOszMAIrWX+CCOZN368
gtrEDqyKgsxX3nnK4OMX14ymgSU6i/sbHgj12SrEAAnDd06QL6hXoBl8Djo9IMQA
IZxriihbHp1yQgwBh6/BsBqrjeTRmt/aNbO5xO7RyjUfv1y9O9LlgkGuNigNlANk
Z9WhSp345HRPlp9KBk4zHgdJlk49B67axH0nWQyP+Z4jTQpOvnvxtclu/Lilffxx
dObsZKNYU3Le4RgjdYDVMjfVayudI01JU9b30hfxmx6684TR2NcuqV5bwmNjQyJU
adHLtbePP5Jsvq/ddcFIcNpGe9sn3L0fo/k3D82+q9ZFcZvlXw7Fa1vcdNRcEKbq
PAwQIdYcZKHVsEzVcRJuYZct+vsUP2z6rhMHKragHNOZYjwuzPrjb+R3z7Bm989o
CWGdsVyn9hyjWyJmRQDS+12dmeMX1Pp5gage3iZQ7MhKr2RVeHnm9AFmPUwamoXr
LdHkgY/5mmlTzkzqqtKT2VPbV9+ZhjBLoIStPU5vyoCeRUmCIuhGqPeWbRuWXwry
gEtDCiS43GIu/JENcTx8MPeAlj7aZR/a7xyDfhmH+1UJ/wUToantAujRrvwAtNk4
DyAmizPEGMj3TvTZWEdTFx/X2OyiZAnpP98obsCMHaOjoeCm7IGbLgcGr7sAbf+x
1GXkJEBcJ++mh2OFmMfvhjerpqOVxKH+c8HFaHoJHUQc24ONEI34AC4IMPIztLjw
myaaBlvkLMfag6w1aPFyFW88GQewqatBovrXHprdr75btfW2+3gpQOoXVGUEsFSY
3MQWJVFv71XVlUTqZLSXvhN50/uj0trVtNtzZ5uvIt4Rgl4wkBADZwTvgUGawEGu
/eaZCUiSys3a1gLJtN/bylq8HPm4WQSzJLcQf10Eriuhgm1HSyyRWHDFyW0jjCOB
AqUSq7fu6fRnFAslkFhQWMaQxNRwYfyineN+YznROsAaq+dunR/GnJHVVTx+HUzp
5Kup6RyniNUehPV6sfdncjYADUJhj9HF0xtVjuJY8wSOiC7gDp/eMqM1B7cF+LOK
we9px4nzVSlac6MVIGBoB+aUzJ/T8fZiNNQ8csBcp9/y7PRQNQcT7TqWui9wEeD2
oCmsoDFUmYm1gAzLgITC6vgLBdBia0CBxsKCiENDxeIPhWverNPhz1UNf2uRT62x
rfaWr7DqJ5dGKkuqgnfQ+vltzXk3tyFvpBEYK7XdQ81E/f0eBIs5ZYvUiUBrlA8O
ZzCy//xmuJizMZraSBqWZcIpzIMTWaWsz0AiFlE0TkCpX6DAQ5XzvS1lgugGSzhw
roc1mCy+c2H/mj7XyNP9A73YV9eMmKlEmdQJc/N5viMtqoKKQcEW1R+WnsOD3kwU
T1V1h+xlMZSkBpAhjFeKt1oOMtdupBKZ1lNTatHy+lbnvVmbwp9Q8p73dPKVDOyv
sHupYiBMZ+cCmqrS/n6jX6I92ZVOJABVuyh3CAqi2iB4ZzAzN1YA3LmBIduwmBYB
wi3Atp6nNLui0b6tSX1TUE9wNdrx2Lns1DuUEpuYynt5gKbwEMsmjqJHZg7N5c03
XmOu8YtzkMVvDZ5/BplMlVpDRLodHvZ3s/QwU1Hmdxg3W1l7JWCV0SyRYOh+YOi1
3wFYbRoELQ/qctztcWHLzSnS4xUGTL7UuNJSWcVgIjA0qYNCnw5+K7L1KW3WN6tR
Nav6HAZDjGTXjX3REhe1ckCvQvi18Ks1xNMPDFr5uUamNq+Q9p+5zKa8F777dxKm
wtT8i6v5YLaBOQVgaz8qT5cnlhPWl/n14z/+kE05KbzOoOThcZQZeOLXbzuzhwoT
YmL1MJKbRe/CFYIsukhp5HH3bB2o4D+GcCmr6mVUwp0M754xseu2XscsFW/w+rpx
cbJxSwjNAR9nLen1XmbM/IucsFU+NCevoUORv9d3lICHhbA2jmqQEJcjMLmRHdLX
9x01+6z70mU4Y2HLb7AVmZDjPG/8avOhqIC120JCiJ19Q1MWi29KkwVseOFL88Ar
Rwi8alhIYyLIKGiYkKhdB9z+WC+y0aHoV3Yc4iv5sLNdxTM8ZGQfxmyizha9h24v
42BvV/5aO2vRiO/0jK4eduWvNAyaGBlNdvvU1XrEGPpfbiPdrkMAaa2p9t3c5VOp
UtU3Hc7MZO4BPeXsMGnMa6gwVBhN8cfYxrva8s90GWTxWtOVc5m6RWXbHe/Jo/v1
2o86mI5TYbw/3FK5r661t4zphmWxTY9/tAL62Cl6t6Igp+5xe9m4+Z1SUCKEV2kE
TghjKa48oAj3NZI0yFx33kGHJemu4Lka5n3KvffU8r9tmnFD1vjregptT5fwWe9I
GAHCd2yhTuXGJQxjOKVelWeHj5o21Yv/cRw1PVFoNMODvGB2y3Iv1rYfdFU+A2C5
dcDGCvsQ9s82MfBxcvGPdaKeZ0R5MhTt6EpkwGmadB5NhVjBAqtPXZzxg4D17WaM
5oC8iIYYolCw97KzQ16jvZBTiT6sSjpUDLUX5jMXZwQxyT5mjNLAGX0khoPBTOKu
s0BeGZ6u27hWZx68l47jqtzouP5dneWjid2g11MfnbokELbk8TDLhAxROFAOaBtv
0dvZIWRxqiE3GB7fwcz4h5ZZFRTwr9VBLp+Je3X+MonJOWIVRKTh9gRglHYgxta2
BkJNGGkUF8cDs6qkeTxRRjqCJXBIuhtbq/AuxYnROSq5Pf4+87g1K9SLg69mWmJN
PSO0vB1/ryTm4mac7ChD/FydIJCM7ZcwwCQj+Ia3mxyR8mSszztWjY/F6t1CTEhX
9qrBWTHUVf/RhrOfpuK9p51ayab/L8TITlyQloqzdO+BDtawubyOabuxQA3CgSs7
P+UOrkdBPcrPX0q1zFdlaaAP7kWm6vWtUdETVZ/vlagh6tSSQ6hHItulqj7PLgju
KFInYnN4XHsIP49RKy+Nhmg2Klwkad2CLOdOylfAk0xwpy9IKXQtTUJfxf5jZSx9
4eZ5FKxhrJoTDP0GSj4KKX+32mfGSGBx18ADhuPeqqr6E0RgooUFgntw6X6sx9xg
+ikgwgp91o/csDt/LUHoIKRIPz3c48oKo1IpM43gaco/OKOaR1GWvaZjQupS5QPf
186XGpS4nQFC+YBIhmmcdEhhjFLRtTtm/Q+Jv7uk5vXbUpEATJiU8VRdtIBuS3vx
bsXXLcWz4dBQtY/dVhg2xlPc3ICbPVqsWrSG1mPcH1S/W0ZcKjtPrFRhbIyJsK1Z
jAMUmnkRUzJk6SMwQa9FY5cJQxb7fAK79+AZwDUtsUjksufameSraTQhKYaoz1XA
+7wm6G+ORrFcBb1V6uoTEhzfed0bplRQfzI/spLDn1EFf97IRNBJgM9rzMNx/eFg
2mt68YUMFwXnp/k8BBzToJTEizWqTLVVM0DX+9bxtScKpejQG8wjWSRlOVzG4MBi
Ly8V88dArqW9E11dYSTVTMG7qBX0W7fx+WUeQ9yYjPpsWCnBN1Na9XUoAVGFo+qK
RVDUfSP4v/zE2mrYCOFgfZOJoo7QKNgXecG7TFpwQYPNXuEl8mMVRBjrZ21J4W7j
2jwiFfzHT4gvqfaGcEZCM+LzFacsysE3d1MWpe1qHlUHHdfvNvWfUT3uQgeFj4Be
r1gnLuKJLfK08vISoWie45k3Ms0/i7xFwFNCcFok2ol6qC9SGgjgaBbpR2Nwh/dU
MsPw6S6ho2ZvYRnNrwsmfZJ3KJmhLSmfB1jI2BHHx2tq7EmpAFwlhyGTIRJyoO6v
zDKriQV866G2BNJw94za9czxmQK//VTZiHNXwqxXz6mYKg17fqo2qooYUgr3Mtte
JzzjloKfZv1LlOJ8lWXjKCrN7u+V5CayLV2NkV0S3hDkIlJnFmd+lqQgLzpNYRnB
gTlXn+Xn1ygWPlcjTBzw9jVj7yxuD9Ya3hUh8qCLZtM5b/8/nSLX649PGb6ai+ZK
OCUIuBatID4kBlXEs+n77R8RCAFAdKQV71+DbKKjs/bU8xVlr5cdNahhMi0p4Tgs
T7i+CsOlsvqcMj4i61eegYz1w7WZM8vBDZNq7KpfR04A8yQm/MnoNFM+Xe8fbfUD
mQVcFcbuaK0KIhRYKbVSPIUBc3PqUPuJt+oZd6BlnxRUmB+SZduBINQgnebX0trS
FTHsreBaO85TwkgQ1i2foSudtb+gm20IG5tZEi6b4AeYvLmVcJjLhKzt9CZRyXDg
4uTbB6PFUGmzGo3KrMMnOJ4EDvpYAu3e7LUwYucAFLIu6ht4OYaH/cKbhqnVGL5n
FxoL3b5ZJ2KjENZSOUQNDO11H/LZa/XNErrHBuinbBAq58klAnBb0xGStXq48ECH
0/HsaLiVFYNPum/UsxpLtuXuJ9c5sfwoy7o5R/nZku2uvhkbmArZ/BJWfv2WxDHQ
O9/wRdnTCqpdN/CowIdaBH+btoRoJzwX63zGpzcOyBevD/KI0H7CjCxMxiyZ6Hv/
F6He+6F3aT/J7L7XSPO2p8VMLAZEgHr6QI9VMyMB7xpdA1XDVevfeIIblJp6AQnA
/ZLAJRygHey+2420aQcLrLLAaggnv/rmvIEOJpMo3gW45/z3fhQhSluU2ETB6292
Y8RCIPheIoFR3xMR4gxIXZPDwRBbuQVgcaAEYnil2RkYrm1kg5JjQY0Eu1pSg4Dp
z9S1WQUmHINnE6UvNTSX2DQ28f2tcHJtPtRmSFH96EnIUazHpxKaz/V9Senb3X2o
dNCX96+5NcSmKmw+4MvwT4AIN6CwP8Yw9gXprVoRjbpSJqqfHvj1+lBfe/w1Gazs
WKuzxH15spsiXO4mYh2B+yZDOa7EM0lrDvGggkJSyZ+ZzCLjBhXD52mApadl270P
qgB5emSjMfAtSnSeqx4dnJm97dIohMMfK2GoMTCRv4QP6nBFhoVp7aNe+mIUaRwf
vp5Rd/VC1tikx+JamyJC5xH+syubdfu3wy3skY2iBzchNEuXnUhdAO1dVl3kyNFB
oXLxzjwtt2gEb7DcoLELNDnRmRvEiHvyBD9n2dYlxa2WHunY3gCDolTf5ryuZ8cg
CfZDLyHDGELKlkYsgaNEfD86kw2imdmhnfalJyFXwC9Yt2um90DGwr8DMtve5AVN
PEprTsur5MysLa+LYoeRN8QvvJAsOBgs3jiYiqCYV+pArNagSpaCCsd9mIHs33Ea
77UyX3HSlHCnc8/mzLUEMvjBCEghGnBxbPkQLmWbsXblrUXwymUtd2HrPSb2powD
VHMA+9wRcSHo+RYCgiR05cYwRocR/aQ0R5HlL7MALWkIFV5FGlQxuCpXvN/cnl8v
4lrUaNBT7TK23DoefQTQHKX29uEVqQmFGItyauxOZ79hYwgHPQCB8PhQQ0K5Pfoo
Kvm76PV8/XWoqTvMRn9X7OOlGhHB6zpBkFLkStCHy8XXEsmXSLK78tfyY2etdoDk
UPg1JRW8q+JhrdKX+Lz6TvRDeEEezKrbvrs2pVC8IIfUgtLK8P5w69JqRJVN4T/5
9rYmejGEn5nvyOdut+CCxo8BfXFb7BBu3iAFfTcPMMAvK6WJsmyU0LSQA81lYduh
IwdEZZkHiPPQauYkpObA8EVuidC/GcMWgIaVSt+FFqdUOF2x9gV1MP6VEUplUFDY
G2myug/P+8zrwmxtdcE+L9uoaDHxQqNe5yKYjrlSAB0Irc3FzOlDg35NZP5RPkV6
mYheA5nJh0fRY7axhp1LeUE2NjqR4UX/TZV441JZVKij4k2a/zsJ3aAZsYSfnYca
ksNFm3IEImzU5oYT+XQgxffKQQA1kH1CpEQG3nDPFLqPq8f6VilqVSQf9Zb26kip
j6ci/ZNSX6lfDbqZRmBMByCBOOEAyqg88eI+n6Lx5cdvFJHkOL/RUajGWTDAPqhI
VEZux+ve+C+/SLpZfoxqicaIFTxTcCfzFPDZBCsOQNw4+Jiq6kK2npoMPdkoUezY
Wx6l+qGENwoAn/90PKGE7hpwPX4rktq6FnJEf6V7nXzA4W0ol12SPBBuo6vQUBCB
jlM3WcmlwTmaKYr+zq4nWznB0yL9P18+Wqxmt50nXXCMqJBvxMlKlNt5bnCDufBp
FsrhinEvWSoKCxmgSGW67mTL/i52E6vYAMkySrM1dd2pGGa6u3EltLxmlkN1rvrm
W9tLx8msqyOK7TYPW83SFzpmtgybpXlfMFspQ8VQL/VPxBBVERWv76G18B4A7ggR
QVy8tIt11ug2+m3IlNrzpAJ9T1hTKOFoqTKaUFYKEgzOTjxHeBJngRzLzeDjhzWY
n41pd0IcyeSq/QiG84ECOYUyndVGYQrI6YEJNVo9Lps0tp/IkD51pPpI+IQCRPuM
LN4/qoVjm/d/GvaAhhF087A7FqbF3HMdXrklF9ZD5trT1UMfcGhVtRn/EdAGRYPR
CZ5RsZAj9SET9Rfa3Nc3j7tHHmVkF+n2OBYK3KmvpkjzfQcfd/c0iWJmoG9NkJC+
kYUIJESwUogrZSJNT/CqkGRs/Zu2GUt+edp5dRcG5UotjyPFuGecmhfV5ESYfzJi
58ASQScw/yRuspyOKuRwT0r8wMHK/uw0XCqLq9mYQr7GEGL/dEETGn5m0t+Ek2wm
J2UfiIgyelPwjU7oskRpKN/+sPsMPyfd0c87cHhecLCwgMEMDWaDpFQwfSrAyLSD
7iTXHyaYCkmYD4GKcQabm/ABUGqFZpmD2yWJdzUaO+/DLo2qw6/Sw15y8pOQX4CR
4O2zRNonqv6+Ry6t0GN5yKEpvxeHAKUahuGWMYNJe+Kgdio1f1Bg69haD997ZbpQ
hE+Lkio6goHvrs2O0SVlqGu41ivdG3cztqukuJ3erVEgUh7x5Els/Fzx80UFwPVk
bLek2IjfCYR4khOBfOIQY/HK2UeUxpitJltRxt4z1FkA8jowhErRlp9C/mvKwz9S
uneH3850mrfl9qTCrxflUlTqfMZsGHFfa0c5ltyYJgIhrINDDvlvT8ZnboQCiDwV
PO2R1xirT/ap6wWXB7HlFUb/J5Af75VWVTXmI6J9psgfCc7ubNgjjgH9IUvA8Y2X
JyBgXK3eDWVLwzK67X+2EkTT3S2s30+fLXXlx9nSzjY3i4OMkY92O0qDsOlUlXXi
fs08lj+s53VYli3/XQHr0LBHEG/FqYBu9FzJbhui8mJyWhDwNwO3bxzCuqOaEUQY
7dJ7F//bD9gZWzUU2cWk6X0E/HLVgqxWHlsju5wFJvvQyJh5OdOOzsIER5lsUf7h
bZSdTbehPjGWiHqjqzkURdHD326dvoiTal3Wkm1YkY/ndOX44lpS+rwS+8zE2VdS
lwTHVTany/KLZJ8gBq6Xi/pl4ph8izX78im213wXpmChd0q2Nst5lWAMSxillw9S
7hVVnZwBVeD8ovH/yMtUiwuMyFz462o0KfJCZMwa5ObewPsDq4twu8ubOfRntVuK
Z9c2xxqRneac/UQDTqdAIS5R1bA47q6WMWMNKd6gkAfj3XaOiAHP+d+odZET9NWT
4TmxniS0Bz8aIthWkqja+ORiXOmirrJndta1oTp+xLUMcKHSFStbHjoybdwLunIW
5Td4P6iMgIpIR6S4SMgklF8sxku0c5hOIS++A0htrs5OURkAsyawyXcAWt7ZYHrh
8WATxGIG87evK99aG4MkN2zkRdCLaEmo2cZu9lWLJEBndSPSR5/lAr8Dc61FmfG3
pjzs8i2s7v/VCu1K0Y2g8iJSRIftqCvtMuupkzHoM3b+C1JJ6ocy6YNf2topWrsF
ds6r9fczcjafFjSa4Zoa7Xq0Cg8FowelI2jFPFPnaOxK1JRbafn4R2b0zb6Ds7v8
PdLDbllaHdjVn+348LICgPnN7OOFKpEwwKgEom3HpvutQ6Epob/yvckvzSbU+atG
j/JVlY1loxG5XrQarj0TNQT8ByllR4sCdJekQRHoI6OJ9HxI7OEhv3AuSlaYsnMx
wxLrS9HaxSw5Dc4rCOi9rOQrwNMLh75g39HtC6J7Wj3/CgHjOQDfnzhh+FGpG/ji
2fBA8wAbkbVYl6t+L1inWniYM29TI5kBVnLYbsS5VKfVGWYLDMzUBIP+4Sz7QgGC
dkSiQsXhS9yXGFNXIDzlKEr6jmRhBXP8nOmD7sn0Ud6VK9cPHilnXVD4pW9N3xEY
ic3XCwwNRvMo7vqHkfXHtEg74QzgfVwaOW4UF519MUc9IqVkxIrO+TZeVkLWoxCa
KNKePIljvaF5k9uDl4eegtRzhhW6OZgCUGPLGFqYKZGQavEosS6yPKQ2YHQY3PN+
igYDRaMSZEDqFvDwJlUQsg3dPDNRTcJ8CIr27VG5ZVB/0Vf2+IvI3FqS+hInuWzN
L9CU+HOblIkQaXDlbCkzYPcTG6qYAgwbWDVNfG0VhM8TTj03GEB4QdeJ8/IyBjSO
AKvBmtLhaBnUIufpbuOZpJ0vo9O54cCpOYwVy+CVS8jwNlaArURpSzOxgUyk4W20
QaOQedrRrEBBT/+eD7A/+NEVWjWh+HC/bx/elbuBA5tbwZX5QngXLahqCZ0pAx6o
hkbmFt3kK4MNCWk2O/f2V6a+5gcrQgCg+XDxFtehZwXDtrYwd5XsSEzsswj/D/y2
HwiaKaSN/R2sjC8BUS5l6WydD1+OZpOSna1cxnGa4Fs5TuxDgs85jE6soFbNrGYU
IaJ3e30hWPRexBN/Xvt8n13tGyPzcm69dkl0ZtuER6oXW7BYbFUX2pmWvl46IEVD
v7w+P9n6P8B4ssyv557tK9La8Pf+8EbTOo5wjLfUc0pU3ekdqRt1pFifW9JW7XQs
jHoeK/oXnGWmyW/4GL8DWIAu28KDeZCcB5Tb1V3yWSgHK2M79NciuywaEQcntGvK
5P1WSj3Wtsc78v/YKiqLDQc05tsu4eRzkCh7nt5oi9ONZgkWBHMEkPpNpoJeUILz
Xh+88W682gPWucf4ardUEMvZnT5QnyL8ii6+TaWERfUbW0dAwOHPgLzCgGiCxJUF
ZafeevOVhTuWEYkdL6+wfu4qck7Kj6kVxZC8T/AhLc7OLXR8IYVRMnCLSXPoOKuR
JF5WF9c5aSONQIdnaSKjFG48/aQ29bbBUnc2mpi6vhPkT5ngpP+fEB/ZlCfqb/3k
JTYghLV2qMmc2Ra01DMRuq6QJqngN6siHhcQxzeJNeQdZuRMkvYq3KnAekSjPuy1
oHeITsG/tJhBhL3nOC/A83Ll0EdXtswAANFwdTbltuYJsYvInPY+blZkcgCMFSb8
EMRPj+75NZakmjgkEWriExs/8aixJQnRs7HGuffcv9xJ2UdWjOzwBsYBu0DQmTWm
43aaF+xJI9VUUdm8FGH0n8Q+rkxxPQGO2Tsm6vbObkqujfRrk6ZK0a/Adg/h9JSC
xoVWNiLtSmoYj46bTek7wJPYFOZFk9eYvD43WuPu/N14rOC8xCmp1MhROosQT+CO
hBNxYVt75wcnpx92pinX3opLAkl32Ot8cVQQ6kHfiw0a5Q/OSZdxuGAbMRmipVDE
KdcvGrx3Z6L8vlakfPgtI37jXkAhEKCYN7nM4GWKD0+zLF2T7kQiRpeav1BR4Y6O
RbFqGRUy6jJaGTL3IbbkG3dLTsnkLUZgmIOC+5u93yh3kEl4a0RQ0UNfk/qER8+p
9dFIjy6/W1GS4lwmCrNhf23tHYIc2RbeT98Px7XmNLo6ZpeZc4bJzKpNipCFSuD+
bmYhiNSm5cVGgQYinWcDPJCFyd7e1/+V8GB7/numN91LeVIpyBnrqVLVh3C8545/
vjEaklLhDibZSi4PnQGJKSFyqHmfXqjAc8OMj4pyGwRNMD11ALbd553q39Rq0RqV
51/gjcfmBUnVn9JOYOrjKbJjyDkl1qNqY++e91yVSVNb7X5VZPAbZXXkAP/lzqay
TAmnOaCFUSitRAvseGJaxBdjFAjbEeg4yPDoSPnEvvFtEvK1ymsQqMVifPbIp00e
exP+r83x8juMJQtLQDooau0iJmRpdJnF5ZemKNKRMlIfy7rg/+au0JvZtMqeuAHo
htjCvAIIG/eCN7qzAMRD2eo7CXa2yu/O9llcbAsG8XOOycTnV0q0cYgNdrk3MTbX
qCsNHybhDh1l/OFB6yQuxiIFdXr/+GLMEiIu/JsuWjrq93wdc54p349BrJWVZbpz
pvZ1WQovawMOG6Z5o1Z5MiOkoaHrJtNG0oAXPu9PPUE+v2GLKdSmZrt1Jz5iExGU
UfRWTOIQAqvIjxjMDbZjAHVBurMCggEvWFcn0OTlR/bdWe4HXc9rBZeUMu9oeGiX
RGSMeaLiRAXIjMPA4jaNfHQg4YxFpYv+qFKI/IKSWP7esPjkGnKJwVttfb4/p5OB
J5NZI7W21iP4/32GeBPnAGjTY0qatmxiqvhZKN2F3kPypszgOijdt3c6ZIewdhVI
4p/krlIOc44BC4MIlI0JybKmMv6ieTk4AnOR1TZDcDuZzlQGFN8uME9GGBf1CKMJ
JlYoLRcBeoMWSXRBRlF1yu56AYsGMumj/9EuGaFk69cio0jMfVieZdyA0YMo2trr
ifzKyBRnr6htgh2eEkgxIHZkvlHeAo9BAWDmT58kqZLuA5fvXU+52yVdPXegBR+N
EIdlKi4mSAqin2+BjeSMqKNf5Ypne6V+5+iR1KBTRaRcFJxQF8+y+sHJzC0EwdUo
4240Kjs2giFnn4wU6uIQ/aTT6toWsKzhrp0NuBXcPyAp/sG/LD2cVkhY9WP2NATJ
fb2WGHvy1y6N58qexVTgCyMyECz9dat2+VlM3mNKBTHp8gN7kYZXiTxnpA6SxrKj
lQt2ke3J0Db0YOOqGeWQqDa3CTaLQrI2Son4R57uGOgyExJTSinl4/mF9HM3OcrD
S6ktN8hBk/mONO1ZGe4r/ogi3PesThEoRcOnChlEvjNx4KYFDFv1HhaF7uG5PBsm
KWopSV30yZp55JcN9kt9foAIN2MaafvEX48QYHI0hDua5yruWmvxGUK22YcRJAUs
p09YX76lOiMDCdUTSUYwobkckzoLI4n1ieR8qL3m6Rwn3wAFkbbYWcMrIMLQm9go
324L2iyrPe2e386abMxI5mKQTdRF5buuRd/mwtNUwIxH2X3wQrvuahoUsTJZQt2e
jFMsFe7wt1DEB/+qsJBumdeh3wFsLWBmAiUas0lM5CLydZ6I0xu9nd0bQGrXoMrR
1ac+rihJBZPX/okv7IOuCIPdnoLRCpf5Jc3EYWAJ50VckTd2dcvUlQ1qrpGc93M5
lMB4i9Ydq/GdTPyaD9pd68GPPsfqGHU98528vkvXJC50J5QRWieHO5a9k1qjXDaC
YnlUBOE4arbvGAP9UV6OVr+fFjiDRvDjikoqGxa8XUudOQLF4NmC9lSdkKQUiyb3
merWhqCz8omgOl6w4uGVCBWBYJ26H2hIjjQDRa5ot56BUQ9DGuDFW2h+pZq2Nkvo
4X6ntveoeTlbb12Hsz5mpRNSnZzPiuO0QbchNsXnmPuHGxjceMmKu9fILmO2rzq6
o7VCdQRXZvKz4kwjd+gVWZQS5a3vuQsKxl48ovwXmb53hbP7irTfCxd10s5f9xgV
GYpkldzVVQjSxd8244DjTVyCZbJ46iyInK8s8FVEsOFezgqtFDzbxFx1GdD/xKO4
t61vwIYQ9hO6b/Y6+OTNNhFYFlnfPxs83ESulUTgS4cHf45QeBUirsUkEDloy5iB
HzTIAsD1Ji/L5IWyY+tEe3bHqaM2gC54fSqTQdCljq91FYKbEtimJAX7ITRjbq4y
GlOibXUY8itaOay4UwNACkr/1xkZoj6wQVbucW8lyXp3Q7/arZZ5V2sSfHZtaNaN
SVejWcALC4TbW3RHnZxoizdn8pf70cgGRXRm9VCLv8cWMVB9Y+MgT1JD31qZRtCJ
vV7PQFjbhwXykwHkLYWIniSo2GIfVUQN0IxgLFrcyg9MUUGXvAg2BU5/iLoGIVw0
oDaZDEMC/2s74AEuqMZ8N5bn3BuT/ZxFMuEs3VBuU1aQv3k9bFHVus1j2jwVDWyM
xKcbWqc+FiWOzfE17pqjqZHeMmSC9r97Q0BNdLza0K/SX2pjZrWFgPqUeOH/moar
TjF3g7FAdT44nrmLg83N7NscvStWl/XtbE1qnal5SZiLyaQVq2vZtNhx2eNugkZG
r+30TAQB5Xlfg3iG91xEINMG/2BFgsdhkjdWQ/Py1OTd2Hevgrw1fmFPl8gvtSVx
bBty/NUjOLL2H322b63fju69RcXGChWkTA+MHN+39FYs+SDt0NpO4SXWM9sTn4hP
rXYIJPoHBSuohvt8zswVXJHUkeVAVZN5IugXNqVITVu2CZzVAp/+VBFp6hXL/1t7
lx2tH0QsNqL0slN3guQWX2yu3JBhkgoOZX6AxlZNueLQNFCWub5XA4E45uDCmN21
O+HWZQnDyGu6UGpmw0OjLegXICgbjCfr19+bggWJVCsM3paNxXJsJvkH5YySzseR
/cU7rUUrlI9Pnjfoa8LyYdphQKrSXAWiyVYdSd4PwYiFWU2sIT1o5hBZQs6rw9m8
gKgJj51glTMc64ShDAYqUehm2Nk4eP2g6cxAOjT6S2kYWmjuLYJfWuRS1l/GM5sj
uW+JLsHDVSOZhZnvNi+lZOK3sQjQas36zMCXjUL7ztx5c1UBIzpGAE5GJr8QaB8K
gRu6w1ssoboX9a5g8zkwUJqFXed0ny8cEtJuQpCIMd2JGscoWNHZ8bcLgymvWknb
RBfaeRQEWjnyN+Q2nE4pqPGCID1QcF2IhAf/mn9ArUwl+ZnYLOpBRIf0hS+79Mfo
26UaJy7r66mNvXMJUAFbf+bSHi38b1t5LAebMNUndeLaBl3OlmU4JiDd1oItY78q
bH+RDy1zE26ZZLN1rcFUMeySWYTzHmBUUtn6g2s6WPcboJ+pIf9WHWWZLv23afON
RIpFyHgqsYDRFc8RIRmrnXb9EnvEb0LYF3PGuc74aU6VCRA+IkVd57eQxp3KliDi
8TdUlxDT/mBNIyDpcgTAwYpaue1QA9h/OG9ZzVVc6sIXPXwx9ykks4Lw9b8EdBrR
0n3xnNjmu7RqVA55pLSNiyqIuv6ak9UhYVZ6XUfxoZUpsPjYvt3BkxNRQsoThgXS
bYsnfGD19ZhPTCBhn23v5s5nFwIcy8obwo9lN+9g55nWSBCgu6FtfwlpsG/fbejh
YVPkKBkOS66zovce7eTZjNOzVAs2K/TlNygQ/zQEVuGlcOt0ALPiHFNBpBozG/k2
+i3nypdSW4W3sEdOyLhHJ226uzUlNn+Eyny4HgJ0m3UvNStkV/Ep9GblYMQPaV7W
fMrTIbVo3NxyG66N7eg55rxi8Q5NHE+/k6s+vkQFkHjJH7u2OoGkAzCf2W0LM/dA
9lNCZHiG/U52Ll0m3v8B7GgHHBz3j5Z/MolmKk+yjPbbHAqMYVII40u9dE1y94Zf
opQczgT+d1R3Hl2kSPAzXfF2D0enb3EqKw4Vg4KeoqTyG6vuKP8dzgIhVDVtv4od
Lgs7AwSMacegGuY1e0AQkaTmn+mjPfbMG5lGJf4HlGmysTEsnvMA3J3YXCbf1s64
ezDaE/qNj8Fv6vJNPP/Xj/x/jjTS1nwFX29cekXS0w6KBwJSX48dFQC08xJ0HKmO
y/sec70ql5n0hAHXVb2wRTyvABCu6IsCOiiaip6HCu8QCsfBpbXXElfQdwZK4mif
4SPhC8jkHuf3Sww5KXbHF5/aKYgDQBbSDGCLokVStOV2DAvuU2sjUtV1gVDJDp4o
VkrS5QnD9TCASHfu0Kpjb03bBxtY2jyj/d4nmLNCcD3HeaDjjTpUviwe0FcTL3QL
o23tsD7kB2eYFgOrye/3z6kbalPvuQWgUVHbF7dGvyQssnoJ8Tke3jlyKA3VZHLf
JR3lesaERYtzlXBDX2kGqIcmNtOblA+CWD9t77rpTaXiaKi8XzUO5IwOcEeftreL
b8QHPyqtBmdbawkE7U4QcD85JKxldFu33fNuuS+xZQ9TGAIRJ1C3K0SM6EipMU/+
kkTZjc8qRo/G3IcZ05yh68/5uY924puVN9r/qhoBXS2VpaqijRbwhuohnIolImbK
XR0z4ghCPFFRu5a/rjmeVAYMuEw+s+g4H6ivZwxQENLGdgypA7fbcDsqTMb6eDbW
c+eWpCcASn1ImTd4XO65xAF5S7rJIXOkuK0WvAT3r9CJ0vipWkbId4+dd5dQLF/J
a8rFZ5KCLESL4kaaLdBppiTkv0YDtHX0nkXwkUhhlH/+5NC1StVuak5jKM2G4e+Z
dgaIzbPpDV3oR2X53b7zQAQuedTbnQ5cgKFUK2XiIgoi0eArcTdfCuHEz3hLgjWE
K2nCNWbrkQD7kbu6BocRTATOM+HmOxxKoZ4byAvAcL0+QouFvDJrKeZraZbfey6q
7jyfLEwuBZqZ+L8ghIdYWE3rvQqzuxuX9WCjktEuyZfti6iJzhui3nv9wh078P7O
fzUXiRETbLeL7qbYzLGwpsUQUkjW595FTI8rkTduXj2B+QJOKYRFLD2OVXib46jz
L+n8gkMK4vg69KoC6FFYPZvEzDZZzFKnmTVSlqvHiHPVRi/KLnFuPgEqg+0anJRn
OrZdCiXFuV9bFyoQUKx/dVRxxQSddqpzG2MgDHOhNe6d8bve5loyNvh/auPL3bef
JaN0UwHQqrV30+YuCeYDGxOrWetjKsXjGQY1i5TVgrLyzbLfiZXrzvp5nsdF07Xx
gRZIPFkE/XplAajjTclZfEGteOcICUEIpuErKhXiuS96H3MA/70yBC8NuBgOcd+x
ve+9kH27JyCyrP8WCEBEe2FhrSnAslrdTBH+y7TvkJGUplUkzgDlNhp2vivZJZgl
pg7Jg98ALkSFWMpMGjvnmhfON/swKatqLZuggpoIm9yf7TaCy29zWVfM31fI8cCF
Ve5/pXCyy3E5Hf5TqP5Ar5Uz0oJw3csLZGUPh7xIRHwdZPX82JR/5qnTl1Vtf84h
oWnE3TaQOuPlUkV63FfR+hqzdXqtTRmPlqYOCgToYAFNHH+2n4PIor0oVZLIMfEd
m1SXv16KCSJtJWHl+FlsmGR/1JF6Jl47I/2n42/ZnZ+ILzI7VhOfBRn5rdVK2QM2
xqQnC6mkXCzHrRhhkULh9gG1cJLMXYtLgZFUuz9djfmxHUkaCq6ejvsyR5TKGIzc
fiMfoMBtWw8vdzghpsVq1OCFSu50nCzCFZEa9cPoj6l6fJ9zx9QNf7ltna2Kexpg
W2Jmrhp2Md78isnkm0zv0kuvAzYNlx+Mh5N8p9EcbeyEqnP5tJ73ZozyfaaV8Wx9
/05YWQMelm9w0n1rRU78F/5wPprKexXCWGVxbVWlHBPHjbLbhI2mWV+DEtwUMIIJ
KeQrtNvMaVsUabRBRZMbl1J4p4FtyJXa1KCsblmBMtL/Oom+Go+YavN0d4ModDxZ
O8cvgBGl0vWnIetaJW+ROath+GUXYC4+UaZqkq6yL59M+a689PCXZPgsVN+LYhSr
7ubXS6grmA+WhmNzCScxescvMqTWAUgdhE2YS/rPvpRKGWWbOYEt11cbraPvBGCi
DAQt/93CoBPlItLRkoM0fP8w9PtFn7eyNrev+Q4nbNqofkbl39c5P1QYpsMfvJhD
q9KGUK8r+voGjuSXQS75FSN7ffHGddCJwyMaGatJ/WUdWYUFL2LwXAgmApfd8iMh
yCOrrN5DPuWMgg3SJXHoArNj+PcLJ8/FwoS/uaZ55+/lTV52h1JEaSZnIJICinW2
x5yUQDuskqi44f4HIzMxiX2FnxGXDcQUoVdT/17erzD13NMx0B3r1YqmJmQ6OHQW
6auk8kXBaJjPJWzwt5CB4EIWwEN3fjzyyBu7N1PcwIsbPx1hMERqeRFWjvvQodHj
HwWfIzuGDB7944tzDPHcg0VDU+JPp1GtweW2Mho13gTiPF0BjTRj8mcNAeOkm/Bm
T28WE/TEbobMjaqghjOHcZgmzazAMxJpUlgO6GZZUUF0B2aU7N3rNRtLiSVnWK1j
jt6zo12QbYnm4ADAdcrCGvQrjHso1BfoU6brnh8jimQhnTPSy7rSvJJRzJH4Q3Ei
az+Y6RcFDkCV0VZdOTxMqh2nFUlUHTLO4UwgXZFurUp2qzYOjtNABrXVcbN5vmHq
n75mKwMpkUqaU5PHqVxeLrBkkxyzM+tSctqfg9bPzYH3SNXvbgOSFstuxFQ7Jg7Q
76h2MPFpxcPW401qRJnOcvS4g9AG6HFMnVvfj6Wm5NRJftoD0PWkTk4MaLdGeF2S
AW6Mbx/TSnFu79FKTtCmXvC7Cybc+Fjom2d6pwkcvcymVmxyk/FLPh9NmjhNK2Iw
bCtxRQo3XVplCcjmeG5xnPhBvXzsjlfckhOz2ti8eaztOJlRGiZTVoK+pUedHMM0
TtNPYM2JRktq7JDLsoq4aTp2EdSKE6jcQUjgZhy2fO4b/zgp0eJnFWX4NkVpoaJN
wEf+gn+PsyIgFncYfpkefl3N3yNlmG3o8wadGbtAJpxKCwc6RQVjH2/+MTQPgy6R
g8H1ULf6xBAxofCgTGucWnXacYeR0j+Gez9MN9R/BmHd8FETXM5YoNoiNxEoa1e1
UZCCYHSvQcQSjUhfomKCz/I5hOaIy5YLrGRXXECX/YUGEKBvEwytnN6BdmRqNOOG
PLgnXTSrjViAPmGGQMaey/LyGf0yC5/yxqu9D5eRiQ/sHQlD3S19P/0Srani7uzz
FmnqKmyt4tsmpFgrJSihZhwP533PjGsbnvSUszvhrfvCQceOb386JK11AYuQPs6b
pCo6WIAq5RW6WHlAnf6uxtvh4Wd9Ggf1MJbD5i16o8Rw7SSxizB8cfD1VTNLvTEQ
wFQg4NBwBKrJTfkzkiXMozmRL6/2QlfS5GLKs2pASmI79Ocp33j5eF/7JQM0DxZY
KpXxzSduyuKK/q9Kgtwl1ug4Wp8gufGKucNxjHG8I7LZ5cJI2gCEuEeLnHXeNc4h
10gj13PxsQG9yunyApZCS6CDzH53rNK2Caf+pW0Qx9KcfMQ38KRqelLTLML1+RRu
uvOtfjTABGnCUvUD5akDZBfy/FBkY5tgorPo/UlauLXjshdtxONdTXdpMLP71uiS
nhX2G0tuF7Ox3Umsn77nlFr4BOKFnX+6i5HbuYw0R69BUXOCNoawGzxB6DZ3iX3K
DNfp7Kp2Cv1d8wauq5TD5Xwm3c4OM4qjqdUsNMwrnowgvLlcbvh2RgL+8F8S/NRK
zjqwHznpnaVn8QURXj3YsVoDGY/pUHaZN/7/DN20546h1qx0EmMllSe7HQ/cMawx
9KK9urF92PCgy2KE0vBPCCFTzfsCplPiXA8PV58zrtEYZ7arCfblE+pAOUqe/S3w
tdRy5iH58EfFdvODrKM+h2GulhyZCZzR8KvPX+bHopigHYUOHtIVYYRtHJ5r4Qy3
8OXWKzPrDiRGjDTk91wopWgGFeDpzEAAf9EYxLUntd5HX/4OWsBZvk7ZWoGMmx22
54KYCC91cQ5l2U45PCtxSooe314V21sAbeI4HN2CsBU4lt01UjG7JNWTVniOhn0G
c3LQ4FJAu01lHXbOANOI6TAIdLkeN+KKVs01HS3UTfsF3xKxgioWRhp3n9kDPCRd
m10mUXHTv6WqJHHfa46dAv3Ks4JAyU6r0eBW6/N/ieLv+c4/fNzaarCo4g7o9Lt1
WFg5RsVFyYGnT2YAXBGbYESc5OPTRGQyCr34j10ydk2zj9uoAy3KDhaB/GewLB5a
iSAlCgktk0Ci+arYcPGwALGdfHAmNX0bw4oAhLo6pFp4LroMqbL6MVyLH1SPlieB
TtaAEspvF4O0KPolBRGbjhd+Phli3q4TA+gnyFGsb5EaIJ/9UAyH6cVDFhHcKuSO
0gPVBO9srKAChgQ25mrapk2n8EwQwCmvwR+Px+ywdynp1UT31saEEreZsg84VtLf
ZXEk89d2IKw4O12nyTMSu4Qlvy6m5B62zdC9erWCL/Mxt5MQLJUKFpU+0FjhyGNS
txkUt0gVdI2WfZpVqWgnDR2ZL7EJxgZA6GZU6l1KLcvTVXghOXeuONMGuZXguytx
PjPdwhAtrjgIcwxzLpT5zQkDEgV7hv1VQXKVCnuVut3Jz3UsPyVVon6vkVGFcDQa
103sNMUvT6fGzCsl9HLnJb5quUnSW+RsGQUpVaUIWaekh0Z/URprm5jzFzevjvOh
ifebTVldeyIeCVV1fdl8zZoD6BCQB3n9otNJYv54oZSyIlCdBT2u7tznRGF3Rnoj
Lz7HEP5bRqGFhiMlrxSSmSB06RpfWImKLEnCdhdyg2aoo/XNuzE8u/4SIRRVVIq2
B9L+c3+Aa+tvXqND38rWmq/JlPnGzIcpSOCY/qnsq8BJd9oHVMclSYMk2E8Om9hI
1LbW7lLKgQ1YtloY2o+O1BrA7KNS7cjm9kzVEM4oQV2ABkDa1Nf94NlwFmTZXOWk
mSfzmhzJFKvmJBpktsZjllXaWvchMkmYtKdWLth31zE+cy48MMrf6QhJbvRB2TIU
qK4cOBowVwPZyp/Z8A02APDWFKCYip+RHqe53R6ceyd8mvmzcirBHWP5v0NybD75
VLtZEUogp1hCvREvyLSxoRokNsJAOopR0gp2DJNBHuVWAksMmFKUbh3XHtOAa6LU
JF9H89BbL5cfL4yfWerJBdU7azo8O7Yhdf0hc50EKWusRKBWdpATIP1vOJdpCXj7
IDiFJSh3YaaUl06PgKrKx1zbmjEPzC7x5he02T/39wwDeIAqEGJ2TfH0zdJsR8PQ
6zgX8ObC679nPm0URtisqaWTXl9CSpQAFOcY5rMP3JFfNpZ5I93qJpwqFHfr6Oaz
KLEpPIE/8Bzt33IsFsJYYknZWrsNuRoLvjrxdwlZFQX0anVXD2dVe/hXBTqCCHmA
e9XItnI/ctaPKmnPA9uxKzpbdmoW873SAm5Sx9NIT3201+iaY5wcPsr0KKiloJVH
D0EyyRaaKRmyEpu4Guw9KBp46VKQv0u+ensu3EBDCk5oZ/xO2LoU4Ahb3YeIz5OD
wgOYDB5Qd/NvU4mSv+szj9UmEtE8D2GushoFrmNTW+qpS8D1bFMJwvXtZ7Z3daOH
958TnzCYqo52Iod8wafgbTONhdmmpVGvyKKL28Qz4a+IuRyA001K+R5ANLEEMjpP
28F45ejoF7WuPMDf3IR7mCpFhx52A4+LipO/twcXx3vVOaBtTHqKUbnKdiE1qPyG
AjlKjmqywAfCDAL2w/TLTXwcQKcbobApcROK+/CoFROZ+E6aU68L6AxZtFA3zWiT
df9emMLY+tI3F6iwgZgWneGrNDrPsp5pOWxpMZFf8438FDvU3fnz9DbxYv1BurrP
anFGFcQi2pKKvL7u+hAdOktNd9K7vUxFLx7MnDwVnoQabQ9xHuIKoN1pd5lDvg4i
GExd0LbkJOFjO9E8ZoJSk2e4nSsXOLMqp4eISzygKmcjKTC7g7XXodKVGK/FPPN8
fYfgxc/9GNAngDIKg0uF79zKjoVEV4gz8sQlOKxgGB2TRONeHAIhgFITY13uefcD
p1UGnG299jeiqqy30IndNx3B4u00u+FvenXTyVgnhgNRjxawhK0/0VJwtJ1qJ1fu
f53oKWufm2+iN9iGmGrhyAnD2xd0Yx5Ucr+C2m/k2sFe1TWaUAO7EMMneRTB76Qj
w9d5QIVagbSr8Q9M01lmFrR05PMgv6Sa0akn6y+PtG3MKPFhZuJONBM7IcXixsmd
bWc6PcbqLLN0okLKSArFH9v8x41xy+WKDzD+lBmQiYuvmMK1uGvHyPzgTB4xEtw4
xg5pKDyfQABk+NVqhFsn2GeaqDlcsGfFlgpKrGMXNQPgMdNxZBQ2vcy/O5FjWwJG
pBhMheBTUAN7LLv13du337TR43RRsU53kviFpt/b8m9J9BgZ/Uoydp9SXbgTv8rB
6OCz0mKrCopUCw6kSd+01zyXJ6OhYbGACEgqw1GAjg68KnWZorCqm/ar6GDGsarS
vjSFflu/OePu2UKJ1TGQAVXcDsC9h3bco8D0IimB+xrAnXwzIbsGHlmJFVNym4mK
7OFIMW9yGSMBTWi8BRU2PlgN5GqCA2FejijgVg/D2F9a5NoqMdagFSBih1gOndAF
UD3mo77rfuIx+T3ZABCyfKEB2eIe3ldIBQs0zV+5VeYB6+b6Bd0htyOaua09kxmf
OdSgAEti4L6F99wFxIvTzyyoVkEP+m7QD9aPPaHV/Q2yU5et2t86y6Wve60OvsDH
NWZebcfZtDdCkEAVgpvIApb+YSQn+DWiuMzoijyWvPJWgYnpe81kjGKVKvAkhvXA
fkIM8m2XDrUwTreekaJ9HVEzZ25Ck2Jw9CSJyI9GSSCrDqCh2L0q+7H0dAPdP4Dz
Tm6PQf6A7rdwa5+T5M8Q+N+X1DfwFtWXHkuyLO+EMubkVqMLbbaiBvdTgtxODFg6
GQWq5Rz1665gnGO59St/peq9YTBassdNamUhoCuyT63+Xbsuw8lXEAOUcaRxd3A7
K3vm3hu8I7zardMktPh5CCw/s4xmXfpUM4M6xmyflwfr6fR4lxFqEqVfWd70uU+0
GkRaVn5TqWnOIhykjVAb4UcIyBTaHm4GuL09F9avYtGNFg4PkMpkaDg40Sdc3tpP
F3T7DCLpDlc4llvW6tuEJIvTa1asqHeuyYk5C4Iwt1zWUxZuqmzcSkqIQbeluefV
D65ov9IxyFs0yBt4RGtIh45dTxGgFNnuIC/fxyQQNy7Q04zaygKX4/hHcT5aoRtI
iP+5FqOitFeqJIfKJvFbIVAn7aRez/dMzFWLQgqmSeqyvQLX6Gjpb77WSR01Nc3d
EKbhC6U0rkTzG1SLzcVj542PEltXM9xg6o73R40G5FmuxP4gVwZji+4G8iw9l7OB
5c7FJZDj94VS5G13p7rzK+crN08P7uKXi/GyDXZ588C0OLxx13vYhOh7OAbK3/hI
qb/PqnLwttGUOyKB9l1KcKiiIMWvzcGMlvz/lplRZsPEUp59KzuKY/ig2uhFqEPA
x2ndlHL7sVqD3+wAdwHNJObNvM+UymYcR59R7ApE7lB3EgpgxbK1dRZNEdvBQFo6
O8JzkW9+oqBt8WELIt7RcqxAip1iEYJOa4lff2a0TIXLMXPtXt99dKvNXIBnEd6v
KuMgOK30EntAAUC6WGys7hAuFs32nMBMWu9b+tCuwxdDzzWtjKu7lWHJOH1N/Roe
SaroSGInw+xnGIIo/YsB2l72bRk0taAeO8cq8U8+Q8+RkZLPQHKE+rjN7DaQv8Om
CILdNMhqc3KqyTGbC+k10w/2UnzhCM/324JLyMVCsTAyceXI6xzyf+O6fCw+Qk/n
ZaCbEG1FbBvN85j+1k1/pz4MY+gJyCewl9A1s8jrpYTgIAZgEqUHd5qj1DtctR+f
UU9vNnFCI3/1xhRK/sHoVufFZc9zZ20y89cegWlgYqsaK9Dwg5R49I8w22bQKQXK
ds56fZT4w1Xn1iJvpLfBzmLu68mgOv2KNZp9n2gqqkY5f5vS0IlqeUCBuqXlwC3C
DKq49355Zm2BYuydGtUmSS9k5gGqzwoJnhYpuVDakQeJI+YVCN3yyHHO49Z23LIj
AZm1o0dGXpFdbTffFEodgeRbbfIo/ksW1C8bxfLyDN01BvJLuAIsvmlPAzs9aUuS
IjuViLuMxqyt7oxx6WFNSf9Iz45eEPYz8HqDil+ccMbXzgdVfUfeLASxfkl5D5yh
boZrdTp3Le6be3guT7fOzVTQzmwe7B/vz86L798SGb9CXnrENujGYR5OAUJXCL9Z
KmlMv0/bbFNgKgsCzfZtZna684TJd7dLBGiUkGMEDDNOncfvy2ZAVAJsFUTQl7aK
Wn4akpST9S9U2NgbeTPNPGRjxA5pWR1lq3PwzoIKtMVe0ODMf9mFJHDIKaO61fjF
A/5XayZyXlbCjLxuD6+aGP01yOeQ9BpPzUviqsHjyNr1lk2XY19X0Tvq21mEk+Mx
15Oz/vAP8G+N0fARV+PpCqOV48+ar9wklzBFRAaRIlW7P/5Cbz5j4vTKQ1P+utkR
aArF5+w/TXwcU4HTfy3/RX49pn7qi3SWSzzLiT+G1umCM/b5Vom5kTImCKHqRN1A
V2lUoO2a8+L/q75ZyWD1T7gAnxHQ+3+n06/pEeNBtIt0f3BIUSJMbtzmzdrZJEzI
Gg4oiJCFj/lfJ5dMbPJOi3ePIGQuhHFu7AS80DQjbzDDCfumW6dSbcx0UsLdX88q
C5lCnJABZA40duiFCreRQS08CtdG9Ax7FWIy7R4O7nXpUVfGWhK7Bcoab44e7/+/
wLk6ZmrjPA3iTNUnRvINVPapAGRwhyMgjHZ8SuuAb/SISj4psZDvGz7cOSNa9u00
O6b4Kcv8q3fkx64iRPUCdkod/FT/pJhgAFm5xmx/yaeMTI4+19Yq2cwXk4R+QVZE
RePNtyF4AudKJWyXaXFQyUx0XQrpLyD97dLMENJyJ4qstCd8irY5HaG3U1wzMHoA
VsONJ7eV3Nv4y5C7wZ0cJe3WXEDNEj7tNLbEJ0k0AB4gBoq7WB0P+73oi4mSCn9f
aK2Mqm/plHNfFtU+6rQl1Ed1TFYp/Ti7WToqDWtm9YENXu1ZzFHaTAJbxjryiMOd
YZU11A1Mhj3nuAgOKIHmf+TyorYBXX6XMOXwEII7JceFbD8MpuHTluKoXrEw8mY4
/2lyOBA3/U+yU4pK4IhBy5T1FS1k7FcLWsz7ES+BYbFGSyGmSYgwqphud3h21xN1
XOed1Dug4Wdzup7srhjM9tBGTC/1wPsoRebszFEWAWruvh32I37MAMfNEB6dzeM9
ZXZzFnh0pYLA7e6BmejfSnqLCKaoQdqJqJ0cz3/u0NuPe5j/0C1PqW6+KCguMz/H
AdBt55pqLs67Cb9IW6/czdEOf0MtwO3fKb5hljJz/sG4YCkk5yZTlXJvo4YWnBLA
/8wXe9aZSjHXcH/qPdwKnhroS2QBQ+N3lQgtd1fShm78MiQyRgIyZKMDt2WKNfUe
6nV3zX2Gbfz+ydEo0l+qlZ8EE/gMH47o46JWRKF3M4A10Fy/QJhQGL8LpIcdd7i4
U4WnVH9NskFxR2uT6+btJJR46Qb6MKrtF+RWBkFsRXFrZZNlF8GNbcf0Tf3p9OAX
pjJb2Cnspe6CYH7NdrfwN7yo3agcAL4dkkWKSeUA8AjZTkrKVTeUEYk3BYdwZQOO
B4mTguB+wKUBe1hjFEEm4zYeN3WkLZunfkf26t5TMWEvVd4NGitkLHcH6JfEOYXN
GU3YkaHbtukHGYP8Xyg03XTL/mheIEu7CCDcrdD6peBSqUml5nOTYvSksHBbjM8a
1pQR2MW5VRDUETTgglyIvcpJ89Z2f6NQOTXbzU7RMXuXCVHVMh5co/pCVNAATSfk
4GH2a/0Sq8atAcVPtFVrRqVwrh2LXK3tPc6ZtmRs+XyQhd2O4Kw3WHwpM7IJ41Zu
GlebyEA/TdLiw8dOq9rrXKpO34L/6g2QyBzrShw6ECNCB3DfSlT39rEpwcgyPiMS
4H5ezMLqU19AECUrgNHtjvVxzYgvYxuVA2c/ByjcBMcQ1S+K68Ol6q9jqSaeGmxf
qmu6+bdhxnDmACng/Wk1azB5ZzdTitA7TltIsskgmgXBX73nkexc6IYTKDF8mgmq
txzk5eIEo4JT09nkGjW5D8qwetseq37ypiK7Wu4vJnNou6RyUyxl6Y2lDTxV6a0f
GrsJcjETblXMsWvY+U9QXyEQoxYBgNN749BYm8AOpzQQrwSeSM+WjInoMRC14FOB
K7sNhPHzYag1ymn9fUW0tJwXUDrNRhY18EIFUk49Md5e6mC6WQp541LCkxa/tuUI
dhSa56SSMMnEd7LXYaG8wSVxEyJQ4dWBOngQGv+XY/Y6tIP4Tg8OjMqe+GzciCJs
aq0aksM6LsC3a51YTnSloVQ/voRlZB+sVxGvQFVWZeBG29FL1c5mlpIqDWBBhcZl
x3oQeIMB/9Mvppd+jc9/NyPBNCjEc8f4OTAHPkYGV+5AdRUuGiZYlyezS0y36Dv6
sSj1DDmzDaON68G0T7Ye57zpTAUHS8G2QMc5aZlcFr8Yp+LYxiFWuX4tFWRbATpA
Awie5+jsG3q8hQZGqL5VvJTFGDPaQ99m/AVA7ZRBgYoqE5TNictwWyDz895gtNOt
NQa7c36OzdCRviPteXcdP/Tsk+p5uFSsSoaGS+mP6SEtLqb4sTDzwIAGphYEWug+
ZTX+/YWuuHVbf7FBiebDt8P07ag/dxAtA7LgUGJSIj3KLDhHH4W0+N3gi4TyXfCd
RrgwNpipnuSjE7K8oKTmbQ8Ti54OQwHgSBh8qxtwmfo25bHQvhRdqeJpL9HV0wVF
33/gDZXQWwrYxZVcjrAdwYc48popVeQu2sl0aKKG++tRIA8bVlBg1K1hJstA93Yq
8imqDIy1v1zwAzgmHtpJ49gKe95P6kskh3iNyWoRdf1qZeRNmD1dJHRWbpbgSm7t
uW5OdpRSaZUpPAOpDNqdgooa/7kioU4u2LDvait2Z0bIk6xp9G0Dr4PdIUq8Z23S
9Tb3Z5a2zKvQoFPNL5gwPju7vnOtBHu48Q08t08yxp+dHuaOtAQZePJQoOwfho0S
9N2dpWf4gp5uMAL9zyArPo42qzT/JyKpf9qAO90CsI0RtbOsZv0fCaCAtEDm5g4z
dZ6sHlpFEANkze8uhrq07dEIDgbVS0poBP2n+UjBUxt7MbkteX45P7Z++Yb+bXeb
NdJ7Z+4KCkoRO+ZXM+pSKnE93VphzEL7QdawJshkYs+JnH6h2R/T6BrW6s4mIvd1
OYz7t4c56T0aBeADvODxVoFSKvazbkUcrLptxSRK0Qs2eRt1XKIUSJsGNty4/Wgx
cEvQ+DhOWhjbxmTIFWTBrMEhvTnygs6qrjmkbnefKJJNe7yMWvQDFwEedikiziXH
77UkCgnD27FfhNk5rGa4j/scyv9C+rl65odomd1+4/D9oDHXIY9N/8OOseP1nBMO
yI5++gMK+d4hofVAa9VAKwDvm2YUXYsc+IwZOFoe5DE10cuO50GtWb0YTWPfOgOB
9fSwzYvyotIF6F8j0gBfMAt1cr+b7GOcO6SX+uwygP/JE+iiEPJAxUkQuAQZwWVV
QNWjfhMtr/XE3NKpb2lbzUJHQp38L+XEMxHBjXlwbbbHmoR45uZ1UFt8WhMXV4/+
O9c88QSOB6LluYwyzLhQNB/MahVe0KW+TrUXtlQmv68kF3aHdMyZ4Ib6+5EYwMWK
qfv0f4XwitHtDqeRzafBfxZFfuNEMhpvyDfvvKVhUsS4lt3Fr5v8/NVaeeyRZ5Sx
kdIF05mpPGORcTilYF2clBE4/enKDntZ2U67+jEZ9BdyC4Q+1+edO7upaEPmmv2D
YbqLLnJ1bBvYttmaoMsfpHfqBeHOLjSNur5MPLCLhBGlmwAQOgPoLEw0hV1SpUHr
Fh3H4PlZpe7PAAfimToS0XqKARrFrL++YW4IuK1Kvff6ZpL4LyqY09pcpQIpcB3j
G1NJYvFOEBXM1bdcw4stmJCuvP9NxEtAXC+FceN8GcOXmSjYtG6JiKvFkeQSZA2A
Z0b2aPYk/mxbKJcmeDkKJcib9dvx08g3mYIMXnyfVjfQVHp6B3kpMwvheeyCoX4N
uM69tcSNRtdFnBpEYy2VZGmKoyGDBiS1fgrNeYPseees4rKqZ4FKOxzCOQYItd8O
fAVKMlbZAz1r4r4OX2n8aqTpKFrivGnsYCxdCKIdV9Eu+VMFa4vH7SGrxegBtDrz
H85cL92H8ZkT/OH+03IBBVMk9cd+DgnU6G5Y5xh20lA9xkxnET0HvPLRZiGcsCnP
77fBTxflwRRNvycSkNaN9Lu3QD/Mt/dcFe+C6zD5g7TthLFUtZFgYLKm22ojWBhN
g5aVynnmLK35+YE3A1nrSLeN3dOYlFT6ycNhOPc2i5cqEl77im24t+P3rm8JmTkG
gBGGTHdyQFa/LIUJcKod+PIdkJP19BZe9RZ4Qhw6CjVSOvKk3fkVWCGWHHP9p2q6
oKsjxOU6HU+vMji1w5Lcu4g8vy2+h4kzQs3LUhVIIRvZxGAfFTZVr3gEHnfh6kqH
/MQRAa6UnBDPDFrixnQPC0W83BXZCZp3ntjx0Opr6DLwviRWITtBU66TFjfhGUsl
rM6U6FnPAIGIYUEW7uDYvWyMpk7xxmoSqGHJqX0+bodF16se07qZehRzdGY+h0Q3
i17hLBErkyK7XUOfdhz2wdoGRpYiwcjMKxFmEZ/B7bz0+8OizBAIAYYPfZ6+MM1i
sg5Y/pAUlBUUV5MEyn4aq4ImUVmKL2puKVB5BaKnrhYS/yxXpONLuNUg/HEgBDN4
RG7bjGX4cWJ/TOpm/fpu6cq9dzal1j6d2VYxqmWUeXwODvuNxGoFf7bQ4C4Ykslf
LFYiqt2IbxlRpxWIEojZgCqH3rfoFfTZJ/yt2MgPHKZwCjRykes38Nd4zhzWgzTH
VyWU7nFDbA/z69qr+FeOEFsNaFpDFzX5YPaJ9iBiXS/EN2v3sY0uvjej0vI9xef7
qqGCsJV+f01/g4zlCNOf0+5a9KZAtwehC1VN7NQFFiZS4rUmhZJcmPJA4OOha7nw
bksR3qrid85qNTITzfE6YHpNWxQiuPFS4mXS7gxDDmrUiyrY2UoFfnuKAw6qkPvx
fj55ONnyGUl7t6ulw8/ZC6IhlNXGpkcZNHroYwHqXlaoh4nvZKb2HPXhBtTmJMVJ
D9eGLJawTcKK0sfJ6+8uLvjhItu1CzVBRHw8fRrQCz84HApuvGieXMpJ7GXEnhRb
ipO858uA9DF/fycgIAnsWYbYkHpXaiqBTD7t/EbNeC+JbxJBuECEd74oSyH1PqpS
cm/i0YxI58cwqcEAILXJUJIio+fZepzaPQM6ul5pkcLAZcwAnwGjvnROdc0ZMGeW
voHEvOBG0rqwqgAAmUsAsAP6L4/fBePU9BnXd8aBOyH+FGeveTUfmGJkx/8DiLJJ
Pc9DrSw3oY1/9FPGEjawCSF8bjTX4142lslXIs9kWjfiwFkecircdiLsCRouuva2
htk9xHt8B7WfgBGyyMSx3UGhP+oW9ck2k3AbepsOxZGW2A9OHFQB5VGi4uHOL1OH
HGuYCwe64S2Sd1xOlsqZsgIG2qFjg+YnDaIRkTrptGg9vx2LaOrHPWEZ+HM45RpG
NpHsaHAMk8uYSVGxqqAi008NPW36/YDFjQLnP0PaSYewG5rB5ueGL4up2dTZkiJN
m34UzWGQD/DlR7VyEaT4SKXzuhcjvJw3oOjIX6XAQTDlzITmZq2EVUXPT67m/Hex
ioDq10Gru6tGut5X3MnM7EGAitthmly6STUv22T+F/7584xMwfiD4FeRtL56SuqQ
PdQUpRHdNs4ThoM8+Yjm34ZkOW8YJCtN4ymnZtQG/IRwRqi/lHRr+XS0sBYQxuk6
hdI0nUFuQj//AfyncycevdC0OZ+i7iO8MATCAWf2UidsNtlyEEm4d6FKjek7X5bB
DAqSBwpfICj52TTEQiMTuiT08pE3JiBdPWmWWkjnMYMjTjcCzebvJPNoOzcPxb95
TZdeq+amYugYbI2MIueKVWFYWva9fljz3A+tSndBuESs898yjqW8pXftkkSyajyx
HT0qkt0rrJv/dyaJBLNsA6bo4+zVd65y/w9wPlwTWQS+08JLVclTSHUjaUFGnD8l
DIzLmUOzpEtNTICjEUAsDU9f4JJJqc/1qeKo5UZuVJSrYL0j4uIJ34+TrIyfLsBz
JLGnpZ5rzMOOc2tpxNuyxrgbrzbwkp1nY8KMObZw5lW/zlcf0EwGNlZ95wImmT2A
YXSMAnnsRblhWuaK1xldXYjSAIZe7yBl1JAvU19KTEHKsy1l8mDNcKnsBkWy9qRN
3oVQmRfR8fDVaoKPXYV0RB0HR6ow65O04Svw41ur2EBEzHqvQGvEAjoUGdbyck0s
oZ4vSIyWj4Poo25FHCEVMJPWUTmag3FINTesYjJBDyg6BMQncILLbK50RgFsqJUp
Sj71li3bSEJb68nL5LOzjSlkrHatjHunXk4k66U2nEZytF7hR2GOnT+m0MEFYfTH
uKWXSVZk4IzFy9wCrJFNjmmRmPNO9U6Fn8m6OeFQrf4rhY48p711TRrAyF1r2FB2
MYTHXducfBMfGc9DfYGREGXV9HDlF9YRja5b8aCEPQHvwoAIlcZPKtXvMMaKYN9a
n1SkSm8GHbma1j9/SQPw6HOaUbg3pSSyj0nk0+KhOs/VB51IFfqcdWTAZ9f+YeZu
LA8VwsVF4iLnheOwksketdRrJ5FgWt+99vXxJH0X1WO1dm9DkG6hHeYruzQRzdre
u3tDW8XazO7sMYFZZdEsQpPDnAk0qWNExr443U7rwrofqIrrB5v07amqxrI4AeJZ
MLclgl0UUY8SYmGOmP2fxKXnpTknOf0E9PFszIJutFFtm1d0PEYODuKG4gjoVvUe
BD74GK9JNksjGH+zzLaI0UDhlJanwAp70qGbIMBMONoWds7AQqeBsaG2vpSAFi2L
GPRB1X7QGWRE+wJ7PGU1IZL1pc9e/OLuvEQvcaa7JxtuhUT97M2Gz1rxTeyRd4go
LQ9m1sH+PKYEM0KzgJoOWeWYCJaGQq8/PKCJ8AJ3TdNzQ/panlRV1T4bdHWB+ibD
WlqpeR3gx9L1MBK+N69IEtSFdMVJ8IojCBqVBty+Y2Kf+CNQaczPjTlGoSa3aqFX
V+A91IsL3etB4+c/TkoJlZm7sAqJEG645YwayPT249tAKcd7dBI37ySsBW7JQkMz
sxwHR4grjwCdvvwW+eqA1CbpFCMqUVHQAeCIc1zjOI6LGNXJDcPIAH8Hw1CGwxXg
1UaGa/8yOyh8P+wPprmL86gKzleHEH2ZBfxY9AwJpM+2s1vfNTcWu8S4AdYpIRI7
gdc+O0VKxJ8I9OHf9dtUBU+uYfMjnGTSoHM+QYkj532nTP0Y2x5bP8u2RBVM71JK
HkX0wxWV86sfor+OUSm3gyHyo8F+0aH8d1azJcu+6xR2W5ME9gIcF9duaWU49Bzc
SgDWZejXJ3UFWVbYXn5Nsob/AQxidwhQngflGWMZoP4FFzvdMHrl7QjV7gFIrCOj
8DKln64i/FYqKtQS61JM3aa3eIaJ/nO78O/+TlbXfxLJDwfo3bOznj4RJR1l+ITK
7O/sTPW3xzv8MnF37C3nND/6xKRMeQmFKqCN5XMz7WT0V5BuVJS4XGDPGpAYi6LW
BbCbSuJKmD7nH+ZLARLRhHpJFBgf7dK4RLyPY5249VqtfLlQO8O8oS/nnpWKOO3i
qNAjfNFzrgC3Cc1anCJiAnxJj1IN9jHd2hyaStOhd0kUs3PrM+ZMqkLY+od2EWi1
TAcG++rQWJOl9QDde9ssfWuCadNy0v/Dlj8AaaBDJdAzPHSLs9/N4ElRdmwIteiy
JhzwjfpPyIYB4AsxZ4dV++VSqhtUsUnZ+joUto/hVqMVPFdJvsTkFuEGmA+LHkNz
Dc3Gyx9HzZxJtAmZED5jwmJSvPopbCBUkDLMoMVQfMWSXSjguZZe+O+qGGkIGIJJ
9dm7ckAZDTuoN0uoFc9/37tb/bqgSb7GA6b9v/6ixmqmphdtxzqSeEbUAOt1s69v
jaLmt30reMkpSiRuc9SrzEeZBAQYszQRcdvp5mLkZg3tnXxAHI2qZqe3761r6pGh
vgLhk894tGZvm6z1gqf45vDdgbL9vZZMH4Feazty0Y3Zkb9Irk+SAxcWvVzKyoGn
VXNiAXHRvuz7rO8p1o251ymMApGHL2ogtUemhSqpWd0xHrXIKNO2lqA+9PCffZK3
W3/CFkzhK5dmMVhxKwsv+NaHHpCZGH2jNgoRsUW1uL1bDKgw6v7HTYx9DnXu7eHu
+McbasOZJAS79VmJmd4cQJuuSQanppPxzsTc6gOcfPxNrJiKpGBzXigzcJH/S/Jh
v0necQyjgmyFDq+AWVE1Wq8F1AlDRV+4EtTthbpLfEC9z2prNw00EV0Lhz04sMd+
hsWmXx1ANPSvPC04yt20YsygUueepLTq7BEMGCmg5vO+7FOpfvOAACvyt/Flp4zF
rd3FsXLBG7orgsDR9i6nqSs5fDVdlNzXygiA0PJ4l65tS7Zev71TuPp+tyW7KFXH
15+ezQ+NulW5eBE+pOYL0ZHGH+wW8K36sxsqwzR+IK6TMjVuS6gESQBspnlJOyZb
hZtvVBoWlfbd4KA/asefq867rLIotlRAGQQWA56PJE07QuGirlmNZOWJCZSYEF3T
tx2dJiElVLh9I0Q8VEM36eBs95RmgVRMJWUKZ2p5VcNcj3r2WcsyXxATGFqXOKp+
y8dDK86tFpp+pbtuSnqbmt3OCPt6u1aI7Yw4NdudtJdIpurBD6NIZu+rXIT85SAN
zF+B5L9dhOpHL3H0SOifnjrgU6Ek41iK0hj0LIDdWhw2LQKJScKcDallY+QYjwRv
OVS4dKizb+kOG/hyVj7YUJ9wFCWwumeiRu7xvM/PWlFn95onKJ+oGYUWW/h0SWl6
qGKxhXrvDFGiEhVKNcy+UcoQ6/IOsGIsuqlXspWy0hS9CBasG0nLy3R7z3znpOMt
GonH5hyBuCYpFWlLxo4MdHOZHALbmhhVB1pTw+cDV+URKWTUvF3SfHU5vycSjDys
fAFNtIFz+OSbaPUIhmf9fumcUrq3uWQhLRZRhT3zWgV6bVKFFWdb0CAW08octJhA
/L57+aLIzpKyRcj92lY8gf96i39h5wVC4aU1iGFEZW4QFdqW6CJiuJUmZpN704kU
8mcInWt3ynDoaZ6SZHkRym2cISv15fuGai02wQf9BfWxxKwWyXr7C5UlE8Som5XX
dGT6X6NlhKDWNP0EeGF/pUyarFTL2Nn4dPQrM095juGGtApylQlQqXINoZa2vEMI
OO9PoFhh62GcUl1sFE5iGF/7u/qUiXyejq7NPVLQmn+uWl/Ol2SkLJPSerU6WADq
RXlzaqUPOJFwkjydsaS9JnNVM0pBjjfrJalpPKthMzpK41D2hsB9lCf4lCi6BI+X
NtFt0GEiUrvoPaELqN+b+l4CN2kYWYEe6hLmZbjo4w/RrfMYxiLulo/LKyFq1Rtd
FtSxQ3Khn5RAG9eDf8n+5DJ50jZJZFg/SdbqS4uz2RZowsfmElGgUZWr+dt2HuqB
7kZte9PiQ4+IYQMIZOpVBIKnGaZVTYmdeuE87E0Kv6T4IZ9MaOFJZ/px6yA6Ez1S
heOGaP2y+94miv3D/CLlMK+Ch3A1iNhtcgOXDWf1yHl3ToE/4ZFYCFzm15fv05nl
7WtZK86+Gs4UwceaNtT1tAoecTp4hBXGJ03q9u5aE8vsCt7Nqn6koDx/uidD7dXL
VWsEb3JKwtcBMDNGH1B4PPtkCAAuEDe8KRIKRlWvcSIuOWfPkkJ7NhVmvWw/ZzXD
xzCH+lAI3Kbb7JoJLFt0eccxoSZUDefnM6nkeEGoZV0zOq22LiGxwndL7G9amhv/
eoZFbRStaAlRcwwKl0nxLbky+q5129+JCdC9QWAvAv3CqghDICJ26iDXT9YDjgMm
WDPamIMeIfns/Evj70KK4LkOt/hUjxI7Jc2yYRTnBa6qJIdwb2fSNGlSF3EAIyhi
6U+cIMqHc/cQPM8A59GLoWcXNyrWkXJNsJmp0P6bl+dUNJ5agi051th2U2TipJMp
ZImQpZuHAvHbGGTZjdM3wqWoHOa2Kz4v/1110sybH8c9rBtrcagG+VwyacMGa8Ft
6IJbmq/pcr/JCmXrKGsXugXvyqUdC5a604s59qKVbn1aAfW7iGUM89+6Ho2FwMIS
Y3fetndjIGBNmAWPzWyETtffCU6dDpvpHWgJeyVDKGd9TDcu6tCZ1aX4k9aavSqf
2tPmnHKyismSYPr6DDE1hXUi8jyblbglZaCQ/LGXx7lqQF1mHT5uWGRse0v5kxsE
bnn2m7UxlRnhEI2f5T8awzMziJS1iV8beilMOLeZFd8bOz9w3T1FFsUnKXBpdShr
elB5VNkCcXg+zpa0xNoPXnrXoiXOvHhWYhCRCBlrL87bu5mw9EGzMZur34hRRvsB
R1QgleTKJoYbWk0/oAHshLw/GGZFp5pw6EZ42g1Jhy3u/PFqai3WX2zPjZttR0aI
MYqqmrgr0RC0Bp3aoyx13WDzzG1MtbazmiLZ1pfJnJf1jSU2CofmkF8UBoFaVLst
1kFWnXzJeW4Q7d0InEW97nQ/1WN2G+mTvzIWZUuonWOY7cSyL/kPihDYZ5JPiGKy
8umV0kDRHu+DCpRBujmkot4D0s3unJyx/hQTkJ3LqDrThPxtTbRVDTsNC2kj8S73
K6ANpsC+PPD/XXSEMBzXWeg686bvEtoIri2TeJ5A3ZZEWs9fSsJAH/3JtXxyzBAh
6M3DPLp/7o6Cm1jOGsQfIgFrq1E6TOn2c424wqm4A+0bWvDkaFqY+bcLIwFVuE4D
jkKR/SCNlUlo2J7TeXNsMGpTpFbJooErlUEHyRPwKGkko7x8bAmvXYEq3/DRVgV4
iyWty7dUi4X/ykMgflxYndtPlZiD2cDI68YkyU782s2gCyINe8CZKuYxRYVliKhO
8PkQ2mPK5LFYyiQL4aQmGfEO2RXooSP0iVVjilASofjB8wGWlktg2AoFbGBg0qTx
6O3X2Cpfjo0emQt1wix1xA9zcsu/ahVmZH5YJa5W3ZjnY8ukMSwum/cY3AVZhpXE
hpVxzsLc9kXB9SVVWUdZhqtrOsahoDlNfgFpkiTuIRedRtsBLYABvWzJ1B2xbeKi
xg/yjnzP7XxkySDIVlgXMCIk0jKa/SLDVUsXCLYC+HoqvzjD1oaAkUScM8quLwiy
9UyyVmIr8g9FHapgoUD0ftzfzIFgd4zSups1SoNs4ar9jGATXritrdusBoVRVb3E
s9/0yRt5woCRI+1oGEuTWDUnj5PwM6NZkTG76Ju6Lnf/opICG2VDrEciDp5NhO7w
+Ahz9RszY5tci/OfVuREr43UkomJe/C9QUdNGARn37d2r2fIKWIaMzySVeL220rU
QKaWpmK0+Wc6K1wvi2QQHYIpRyu25OV9/K4DcLDaomrq/mWaUPVhp27Xnicqrj/y
nQvP4e//DuzB3p/9Tos1wmGmeVB6nr3DIsWQPlSlrfwMJWeubD/eiW8LxIcnO5N8
M8zVWL2v4Jo61E+fmcZWiLQdPOVnd5MqzxHNIcT09eIwNXh4GA/Oy1gqHQOw6Emc
WSVDmahktAtxbtd0vTiqsNd0pgpY4VV1CbgFUpVssc+woODaQwWg85hpr+rhEk5q
Bj0mFzdjKHjwCmxWtDLBVKuq5mD4KCKZzCZ8Sk89zsylszjph+VJrkStA6o4S0J8
kvlJy8paI1f2iisEeRm7/FP8mV0d9oCp403UN8sBOCyVrNixyH6L7pwulwBjUe+B
MCAueWkMGgwhtqjn9yF2aptrgVMmf8CtuiNRBFdN9Rb9fdvNnfIarqK++0/Xhbxe
bJsZIKz/thfqCe7Vh39ez4JJ5fVNN/zrcachCPoAmwC8ieP2Mrta888fs+tHcUtR
8vTA248uVsMtqGYLvn3OChV1O83pTIXh5PcJdYShgXVnoQ6JcOR7iPBV467keUF+
aS/ssNRogrXVUAsu67RULqO34UFPt8z4WTw+hsetAUCPsSF3UUR8xOlG1imt20xq
UUHTG67fFk3mH/2klPPy9EkPcYn5yxZcViDW1MSFLc6zRysRqA44p7Z7dxCxtrPy
M/L/fK9qwwFFkLT/pny2n/f+jviikmWiHlEuPTfnu3EsrYqqO1rBhnD3lBPIHxib
4nAMgryzkRwe1j7pEedGyo2GxeQS1+N5js6J2BcPfFwmjnqXSPycHMnBQUx+36Hf
pG1tQ9kt3cFOR8SDnwmmDJaLL5z3xZyP1y7YEiZdvgDYy9PFtpshgK0G3QL/0owM
Es3/QTntK62oE3zkb4YUYZmTAVOPwIe1lvIvyJcYMPSU6w320qhOBce+65VSExl7
w5+9uaXEP8naeeSi9XxTyiuJogHS1jm/o1/C7kKgdUK2YFvjx0JRrSiKeTWp1MNS
mftYHMlbBFV6BlYA0ICPtbH+dPh0cvuUNOzEtiFEXhtJdwDryZ9lsMceNDRyXwJW
s/uyJyM7m83bDmSSe5/gVIKJ2i6XN6XTD5flYm9xb79a35efhSTyP6K25oa+XPa2
SxB3TAm28DC5hKLN1q0nOzLAaUoMfV4oA8N7oZRseBgbRRSuZi/vTmmT1TgEVVz6
o470yDGoWG0b2KGzVKRCMtypEnQVU2Afmf2UagB23e1PaqGC3IHuDoJ4bLSbI3lW
ZL3HmQ+tV1tY5+Xm9sBqWz7wXN2z7ej8LH5UiaS256cj+79BzqvAa7cxxe+Ax4ZF
93VriV3mSd507tq1D+M1xJ7cUjGS685D1p701EUjnkKLwlut3ahTa7lqBAcaW1m/
7H16UvqQEsPNXFllulDowGHBPFsDv7QGLEdsDByq5YqhA/SloHzR/FcHdK9er+F/
uAH1QWw0qVpPfsGMQfgnZ86Xy8UuNY5TBBeWVd4e9mHzphNGDVmOmP86/8LmEnCU
mYJxpS3n5UbKxO80f1b1LVnyl+IzgVwb+Y6rT6iwcdnA2dc86WQCAiqrc6uXUx0+
c06S+DTo0CugDhq1YJN7+emC4sTUbqkDpLYMMztUN/oHes8udOxG1m1vsqNLJ4p7
JKCLXn30osnOiotUZvhWcYr01eHKjcicLJ6Dr6O11x+J9CAoBECjT6iggrp1/aeW
MSxGsM9CWKmvNDJ4Iflh2OXBP6FrmaQuBwi0ruzpM4LmYvWphFePYA3bYfNnfBE0
6ueGO+TwbD9alFCVldhgS2byzAo4/lT8kwwLuHEFkqntJhU/swVnwTtHja+CgrVC
Y3klgFBVIzC1lcHmmOPR3iD3N5QgekWGOPxuFFvaz7Xx0PjE4+QrKgVSFjhdm886
iE0k2JYLNFfCCIPeMrJsWAb1tLON3QF+WG4PLEzgTgSq3ZVv+goU0Nhfu9Lxbpxo
yDUfRzQ5w+hnoGtkgQjnE9fDJtWLol2h0NdOMGxs4Gq4l4M80bnRoXcrn0qDewMl
tk+3YAW+7IqEsUlEsuamYcr70Gff1oIyHJi9+UDSHKvvqQ/l8BRXttGVipl2Fqm3
QP2Dmtv9tAvGdeuYORAvGI7G3Lg9xnM4AZN1olv9quobEL8XdPmAFDK3GAGIM0qd
VMk8XOhSsopNPh2+0jzqh3J2V3c9o9/cvtBl7rRBZS8DRICdQ6BUE1XOEbiFPXrf
lLss76eek3ZzE5S1tww4k/i76/Y9pkQHET4cy1VLxIUfxcF6TjUr7CuP+4lyoKoX
I9LVNZ9QHrYOKBhSfxBEhMUNz9hhe3yQ93URrYtg8jHqPaMmxt4QWUxZH9vrobsS
y5+3DCz0UxWwGv0ciCXMypNHcS51j8aNlUEAE80VxI2Ulld5ulkvPL/xnI3FsSat
L1CB/BcUMsn5//RVLyhWR+ecvWzC/lZ606u/JRDRfgOlGmiN2B84VzMwY7X6B386
69YmciZql1bUa/hYQ6CQjCLyMtedirVhTx0eUnlj/TCWUNlFE7qp1HEgGq/vZYpz
53wcZd/cKfWs+2W5nZNcRtJvCyERlv6wy5FC0m2U4z/acS4uy1jxzRp9CxNsBQpV
7DQHDIazGbvlgcxImhKWeRL9+ukLszlSKdM1rHEVVLuEi51t6WvZxXBM2i9sQc8d
TSRj4/GCMPtMMzWRkbkjCRpBnauyCzNKedu8chEeLPbTrs+0+uCLfd9IOTszTTNA
dlH3HS2ws5gQDnwMmmaoC8faxod3m80Y9Z1IJPQPRdrDdSR9GgNX+TuWDHrSsoy+
IUG0uLj4RsGENPV2vX5tUf2adHl5YBpstrdEIQcx4CcLfbqW1DaZ35Sya2m56vtO
GV6i1RMvV+rpjiFVKyLfqpErmxVP1JgnFRz97IM21nT8qgsGrijwj7XrpcPkBjJ4
KFJIZT5VpFCUuvZJLAOsz8a2e3xd3/46CckmPv3dilh/8QMu/QYnd56zuMshlJgO
HYD52sfi4JHwArpJzMNBLKdt+uXXdMnetEjuwBShRwEBSaBquEyUL9DUBgabDkg1
MSiT+7Ch+Vr857W9yTxpbcE6075PD+DyVV1I3ou9AlnfAaXR0HodccJ/Mj2Ao/t9
enwNM8E1IJsEjUh2FZQl3sLm0Av2T7RqmVWHAVdviZUU8BWMGxZnDR1elIt0qFni
rW1kco2t580VLLpcgEQB+0M5/Ard3CL39FOF7Jy8JJy76uWW4mUx4DjtK+Mprn0u
KBpkl8BxJRcQ5PLUoTRgX2C08HoKJ/v8lpMANBTOoO4P4hNF/DTONwpugpE9p+qD
QwEmfX0XH8mFC/POieOPMb9oa4xTKunOqPf9UEmkafoXqkQI1oBjDrEbjBCuSjjz
tJTHqb00NNgbxmYXy431wFuS8uvk02mnxv60RVJd0Ma70v4dGFPKY8ZCCOUB1uJn
ehgAg+XfUptq/025voqMKA0iQUUKOan53avNZ4jEaj80oZVrmNmsFhSMp/pJ3kXt
liyy1nPcZCgIur9qpsggJLLDS8FL8jLch5XAElhxCzu50AjDlt/JSpNThQij8sAL
K6bl2A/wwX+/sFgxZfWBTboZEHeLt+yWkRADXK6SBEK2KA3jpbnXNNgtCItnyFwl
nLGObWRvd4vag+rSj6/nZ4ZpY0Bl/rO58Zv7MFuicGeT3W8Wf/23ryDOCQ0QMfO0
KIlFiw6Z2wTFMgl8m2hLwF47F9IXOQb4blCh8Ld2XgbEqrqMJOsHSqwj06Wa2vSF
chz535L7cqi9lWbOyAVpMtv7a2HWZqIm+D7lpae91wdjK94uTJUpzf13yRJXS9fJ
Ug+eg6sQoh2gcJVSxQWvSypGydTi3DrtHCRPvbjx9eICQ2YEs6ystLe8YxpeDb16
oBuFp0IfJHvWdlT6FqxzY8XhKAPFP4dlSEj2ARoKoGh0C6etNNb91g8VsCHvniWs
nXr8hrufU5Ps30EGbr0aZSd1F/Fx2Lq6sY1XLOYV979bLJ/YpMMcoFaz6TfEJgzR
rN6z6vcgsVPv9xAursI6BgW/6pKC70S7J5xuCpF1SsvfI/0gAxw/eOVbKcYvpxCP
ld2reZ5vunQrY4MTT2LYQxMgi7O9UhgLC5hhH1bY2bRubyhHkMvrrXJ9O0U4jCDV
u7h1a9gEyG5HSDspbGpMK7y501mvf6x3+Z6F9ChAKdB1EaV5/FeFrHqz03rRGOJW
htugD6DgRMSnqHIGf12KUEvM1AGdNkdaJpSaoqJJjigh6mBT6v1Z8EZQS+DkmMBR
Nv2MylZTeVsVOY4dWvPQd95By5cFTjYckv9n7UDBwJ95UZVK7qGz6BXFsyAcamHB
5H2vQ4yt4SrHhuorafgk9f+soDLb3CZiT3miRDHuQczOK9SLyaBWRuM2FnI+og5b
A567/dIS32gUUk7uIGhZ6cpxLk8OVgfdYNpg4UeoA5lTtNypSpaGKytNangeHDyz
ISB7htNNJLYJxLqcoio+AyYkTXfGujF0m/neOeiMFOmyI1eQzD3pOMj93LTzOEiZ
c1dyOUMx0YR+/5VTpKg1kTJUidbVmPY92wNggX3yeQ4yh7mJYOvfQU/GhLN/L2Mr
4o3IKR4QO/njkmzWgAxR+E8RJSs5YM7dG8cc3AChQqUToi5/bnpGzuPgQW3/InQH
qUED7Cc6R45jx7m9K7Xqc3+YljBjVGK39C6cN39NgpTzyMV55/Js1/aYqLgfNZeF
SksCrC+Bt1KIGtqWUxEziD0A8h2FO7JeY7R9Y9gFrBevZiwsmbtmsN9hmHMDx3h1
ddIMxTv1hQOw00g32oV7IJOB2kHSwmzFMOEaXUWqv8ICHe4l+ZHcyjZBRIKDpZ+7
LokrxHfM8OZ6mG2AYA4BCF4q37xuMEbl9hZqzuVIz6ccC3zTcSB6v7Bo0iGWe6fz
WkQ97UIIislFw5W9fssf6PF0C3SQH0/yriYH7UvNC87XK1xH/nwwuqsUHa54pVy+
yZBd9EFmwSub76jF8oOyUQZrkhpgGcm8l1P6cLuZmMjK0D//mjTea6XkWH967QEP
LZ4JF8OrzV1ZZFnXqQOQi7S1w1nH27DF2nbDgyABa/D58SQGXypK5IN1RQ9ApTTX
KJNTn7oPD06TfQry4GaPjjfZ4QjOTF7iGyogl4vG4SaIlXuZnUGb7T3zCdTMqEBz
peQ13CBrCnx2nSK31a/SZuFtspg1CA/rRT/NAcNdrEtPtxIl+Ko4lQ9U+QVk9Y55
4Jg8oyjWiKD0vd5exS+PW4wpnEYfZ+GxJrVf0o1P9TMSO5swRzPxEDdsGBSG9sjr
1TDh9nl96/BmvlrmJXcfOYbgINjo3dhrBqemUvSSRjTC7cAdzdgPlReS9/2hAcrr
Ubbi8uQHicKXpcLPQRTpkgvemqDrifnx64d2xlTwCg8e6I1ay2O4Ci0xfDMt0Sm4
e9pCmqaa44Gnp3PukA+YMXCXiw6eShANU1zXrMk9bqkZ7+afFIuYblm93rreoACE
OL6N9FhryJzWj9REQBI8Qh9Qv1lMIa0eLSTazEIjZhUSJwy1G0w0V7H38AvMrWhS
n+NFOnAm+evl6XFg3SB+jut55HGVR7I5Fd1hq0HsUiy/8y+maDGuVOLoqCqXgZXt
0C92ALRDZsGrylIhOrx6fPyje1OAuYIKpFDjpJYli0844spl1NS0UwddxpqK8YU3
OKCvUpQ7ek0otZ08N/OJlvLRguuUKYZArQZy3lHAmzwHjDA1MyPwkKUw/da2229x
p+TvwLXmnQ13h2bXu7NT1rlfrbiD4Fiv1pdY4H3JZOXD8W7lO+5WpbOQrX5QF8bs
KzbWYI5k+lEUWBHiThagKeRUMPy6/MAol5KgmqSO5NY3ln1oERVT7m//Dt9W2VTo
w4uY6lnQmTjcuogIi+BMIqeBFuzs0OrhihG08wvgNxss8Zbl3nwu+ehdByUecUKu
SWovfwo8D1bc4D6LpnsxCuAJcFeyRWNh6wYVM/p0fWHukfbMnLfvsCNvwimJgs3n
MaAbIbg63NmMHGuUGBi6fOV1QY68m17HO88oby5c0PcObrbUNYCxMYOmxk4GcSTe
Rz8aql2M/QnwAlc6pnEVAFEtwNcMFMvVEle1Z2UZDlvwj6z2kGXfFxEdgvT10Sb6
IIa/q+NPyUeEF4TvXEyEEjw1laavuYSq1SgfGwYFI1wD90Rm66USREpNRtSspBMD
Pjjrg52t7TaUe9dc4wZaxuPD00P6OrXYuNbOzA6r8ezdv2/3VUFXm9Zt6Y0igQ7p
CGEh8w7A7I4e5i/NbDQzjPWe5QgRTVqEqCjUAHxxdaMckriFkiIya3s63IC2jFEZ
50DAeg/S41u00xYg5TBkxx6lRIHKjlk+5MUCxbNpA3HSnlS4hsneOtJvNp9tW+EI
k5PdRbGkcgwi9fUugJwyVoCBs6KGWX7P4zG5Vr+KO94xUsqeT67ZkVrNV76lUo56
BTyS9tEXGp6KJAj2QE/Z1f/Nm4cQW5hhDttEVDAYR1DwX/gIfnYQ+5U4sRWX8oSK
/vPFc5qfsEMshVF2IM2yEIsFMtjSsdvo1ZPiMYyADFVEGaptIxJVQX6FxMKqbb2y
Gwm9Ldcq5+ssUsViBM21AKOjucczOvtZqppq1mUjE5dHovp/WrjjqUnldbHB3ZXu
gzfB857L500CWJPZ+vZpZ5uK2xjLWxxpJ9pwmC0wDD1Cxtgu0XEOlJ0OhPpITWUY
UyUut3xiZbtTbIWvwjw9zWAUfLKyCXMP4nFtZx0cPEcwembs0W+vNCb5IDVzGbSj
R/bDXOghBbWemzwU7TF4CT3uxtwWZwnYTTXNPp3RoAlMInJDyKhRC8je2x5fdhJr
u4zpg5QQlBlfxU+zF7wdy0Lwf6JVQBopavEp7IPPy+5pOhZo+VZHZ75kCO8jkkFL
nARmJgKXOsqQdun14TqYD4E0ckrqXNifVOZCyjct6YoOWQCj9honqErj0n/YA9X8
SHpGWS+jNDs5P2ApMEKgVcAx/9NdvQrH7DEx21AfTpVGk6H5BVS4C6CHJgdnip1f
G1r0AWmNXh9H/+geHW65xMQAjrampp23m0Q3tR0fCAJ6sbCFgz94B/eggSU8YJP7
zw8wpUQEpdwsIKMz2n/Iw1r0BUuFst1hhTSV3Q6AwrFe3Vd0Hfee3C2sdChOtcE3
cFxzBRB59XhVi3naHWKSA/X4RUSq380lvDOfLb5Bc6Bl2aKG+cL7mFMGRx6uvqrM
ekBaDjDUqL5tSoBnReCFF6DDsdmpGLFpbcyB0btrZ//pv1LrorKRWiq1nAExo5he
psPxvGMrH2svn0mm9S7bDSx9T+hXlRy5Ndc3c4RTzXJ1Vfo9JNznz2XbqP5166zD
CMN0BEe2VmHMA43wiy6mm/tEbu7H6ef2KucAP0OzLDJ9BJd2XkdDMzqqf8xfRAOa
P0EawE36hfapxjX8On94Vs1IXagsGYrmS/j2msWhiUe9IwCOIZygOV0Fd1dRx3yo
dXvgGKL4KHvlV45BCsdknoLIsBOYtFJ6eoOMyQodhZIxabS9ERYwvIq+qltC6a6Q
C6wWw9luOoeGVyzi5qtzycsG7mTMru1bv3F0K0GRz735H6WGQVSjUx7b/8hUFuIc
dQwEBCfWN14+ymNNTsYcXiMszYMxSB13demSaBKUXtudqLyukE4A6BcXxEimvQ5M
tgZKcCTCmvVcF+EOi5j/VhKVTumiJVxKpsIJOtTnwV2aU+TguOMyE5WFIfdYZh4D
QasXO4MsEuUc2seSn+UMrLn5aaFBpgzoWhBoHjLOm0zPsSqHIPH5p/biA6/h3lOB
VHUVsg/opkd3MBzalvkKHsu0HGa0lXUHO+DCbObqEck8DEBM6Y6qfkPqKwAzh5zg
suNOqQ2SGlrac9g08y7bRCN4OHj/er117gVXmM66jMtuYBXe0sBA1nd6gkamIb0S
ButBA0m1zYkjfJ1sbkBLWklHQ9AYJIqtHEa+CJ8toGeCixdiwqSpeZxS/0XcCIRO
vjoJocYFx8H3SOHpnxMdNK71HSgTnTH91ttB2B3C5/7pPBJ0v3+Ccc0BJRO3scC2
CG1mkfUBm8G7233G6jDJa3WNdEts5UAhVI0RhyxVfntrAm7b1ycqVK0KSFXbhV4I
tq76Y1IxKbi7/Bt7WipbapqsQwIo+JcAgQ8h/oMOTqrY67+i6HZlaRQJOKVzGt27
nxxe3Tbd7Eqg/nawyB91gUkN7azuPD7jwEaJ/lkSuvGQXR7vtB7CnBRSjf1h8Qmf
ESFoSNrqbeSHf9i6MycIbx59TfHcWXH24eMklHbWTCqtGEF5ZGk0wsJaCcUbwy4/
aP60ixTlvlx/cA45RVkwVtLK8Vi5Ru+HUuxr6QP17AaJ5t8VYs381n5mSKEVhbOs
NEQzuWPGl+56B9ABXwm4+nVf+A4rPXtRZ+6QBk/WiioosFkgZKTF6orimbRsBjk3
XNmxitpPVZ/ECWu+lD6hy+2D/+X+akxBiP0gwPZhJp+iST0ZJFPYqwA17GgGt60D
A5Fg8xOQsax9cIzCLCiMXjgFRfROdUHZxzgPCRldOgCk3J7IqV52H0RLzj+WWQsl
ZCb2R/1dGGxTPiaeo4V+yEICf4tsKy1N7X2bVHldBklQngkh701aR1SxvYtnhc0J
ZVPIKjvuqe85TrQ48c0QLl5z9WSONPyhFD08mMiPQ/O7+1mN6TfMOzCw2kwojjWd
C8R7Qa/epuHe6eFXuWIx3S+5jroAt71RFQpaiuCJRU2MD21PykaHh66kmCeDP7x8
qiZiZF5yg0DeBIlmPpK0Bblof5tCREG6/PF0korahW1iXCUc6iASrdsMEAFK6UE3
rn9fCzlYM5Ubn0+3UFyKPFveAgeY9MEXeZYBVqJEbj7Yk2EDpgS5E5oUi3Hi1w2a
uDhX8bdnNwl//yhnO9Gu1qIcX0k1ptG8ZW4osqZ3NV2K7X+ed/EYt6FeQa2DM3lV
rGotjFyuuJOtIeIwdnSy0pNbX6qnudWwY2g+LwSyhXyXVrErEogLzTCzjykpDLzb
AQMOlPe6ujtwinLVV2vIfmgb6frUJMdjg5+6TFVWs9PBrw7hwDRo2vVH4bJfsOK9
hMaw+FXOjpTdpeP0tPq6Pgxy/h0QgEJkDLakeRSzRtLy2MScBEmpHYinj0WHZCV7
eWsudRW0gTeT1ST5BJknT8pdcIUeeiLly/9a46Gyt1AlnCgkpJIqyC46ew0cV7ly
n0C0DRxV+LJnrYWmWt4rhXy95g9V6I43MptiuWr02171edld7FfSgHrwuwChWTQQ
lNhdN8Agboq7bxtZxbOg4/hSUbA5JgV3+AcJWxBBmVx0hMyQeN+ckkxRgATDwKYk
OS2WxpS2hLlItNJvvKFAI5gm2rk/L4yJ6n3d1uVryFu8ngLdUKkIThQm3pYrDlF8
+d1hmPJoq4GjNfnTEIQPvbcc8EczZS/0hvUy0T8YNu71VkCubU8vHa/9m2NiZw5W
PCEod3uNLAjHtCoSJyHik+5dHqHgCpTT0jolPVawLRYrttrCt9amVliE6BoxpxyD
JDfR7XR7LpS/uAmWfxygyEJhBlncwZrm/YEQTbYSBrlp4mrkdubId4v7QC7/qAHE
OX3GRpVn+liIeZiEf6X8pE5LYacfbuyjPYf3bvgdq+n5XjMU10uQW1fkDb6h550s
06kCIMtxI5muSo9kQA/P2gGNPHauYXmOt3M1rsqcUVbETDSBTU6P185tyEmVRh4I
L9+j8alKhXDaC8VJBHAC5jlSAxnDBDy+rIh64zNlIH5lTXv3ZiyL4mcliZS60QVj
EOVe3opsNgqpYusq1cgGMaVxVimGVqEfPcydD4DFLjBg403JsEcVuQKcl09Kz+cX
elc52ZLvYv+LKZ5X+3yT4I6FA/OA7h8nA63SXbeDYSF+4OJn7ksGBFMoCTAW9ahH
12RZxvVReUfKDQkyLkuoGPnoHGUdbuO4LunEh/MxaqqyGdDwHlW5/UdIYXsFHuha
Pq4Ehu64+6prL43Td/iS9hW0Qz6yCTMSWTgZ29pigCNDyLbeO50O98WV36NyYXPP
A5RK6gcWT0N2QBrCj6K1ACNmIJZUo7hRfyzMQZk5DvFVTuzmNt2KxwIt9J4mZl8G
PBqW2kxuuSJMSJI6t9sclssrSDuG+7k4G/DW+lPzS0aeYvatduVcovYkDau5U4TY
VuBU/ktT5awdeTOVqr/TY6sPiUKICplpnY3wZ35hIFH5Bg0KH6HPqEs6okvPERGx
IK19dRC24jbibrmABpYEpU7ywouiPorcwJBC1wU7IgSMkKI1nrDVlx8uPonI8n2s
EZD6m3nXoDCnxTzI8t7ePzlwbSCVAt8xC6WPXAde0GiUnLhhWzzDgsFk+Qx9ZHie
xDcOpA1r0NAgv4PZHQjYJ/5r6xbSfx8C1PIgzplv4gpJ0TWbmdpdvbNNi7CC4VCS
lFnO7Ne5uersyg1BbH6L4j+e+iAI1xrYOsbsE5eRcuZKeV6b8YTWk6t1wcNwLn0F
X70rTdV5DxYepOwiFPjldqFoIJidUS4YKMhBHDmMqEYi0kDiM8j0N6adUanX2E2i
wvwJWjViHQcumQ2FjmMSY+IvUw1fWeEj0rQhUn5HoYjTwCOaCJnvhLUyCMLJxB1b
55HzpSFMTz9HflC24wtXRiuqoM3YK2I5vZe6u+2kT3bx/3mUAY2YJXe72H1ynvkw
8bfOy1xPlknkzs6CXMXugtbrU6LjgMQlSr4NUk25stt8QBOq8+Me9ZDqbXrVc0GB
u1AnEcJq7vuY+4tafh6STpPXpTf2Kwec59QZc5VX6j3BpQHy7KgDHKBVUpmS/lY7
2OhzguTaUQHSld44SbKsXwM3u5trr/gI0yvG9T0q0bjREvY8+Q1MobvUpMTotjB4
22GmPUZN+AARXUS3dR4kI2BvS5qM/uEXVibZ35t3FFJoUy5gQF0dmKVXjCVLju/2
Do7sw7gkzhaiKcvuqldvE9FhwZ7yXtC3n6f1+dv6Up8P/aJVoDoaYglTKrE4fSKz
P39C6hnYBMvAg6ad7EmzZpFlbNLGeyIA82LDYj/7Xa3iegLqyiqxspcMA/quQqhu
OD1DSVX+PjT1rNk6XoFCU/qHnxlklDpXlfq5BX615jxOg0ploRiTWdG7MTFWi1ZV
cARMRz89gAOC/7A9XCgFsMtjrD+sALzz7g9gjzRsvXOLO2J5ZdqXkGrCbvERSViI
CBpjHI5FDlUN2F6GL9iQs/7h7f362X297FTuFMK65DXXDB12+IzXYkt7Ag8voC/f
VHYLPTIue3oMYF788Wnkq4JIt3A9cc8JQ41+4clWiDf52sohqpiN/JuEUcu5mjHz
yNC33v9Bpu4WjiEGWU6HBBwzEFfsy5Ns+IwFeKpCuBFd9BFJvaMTgv4jx6U1/BcZ
YZq9lm+f/X7qogtqsalwyrxI79i+dC7xJg5cSuV8qlhP3VG8AFk6gxcUsQiecp29
+7poTEqJbxEcr3cj0uJUaUZQcEC5o2Wa+Ti3c2Jo8lavjGfThSiHs+fGYqxfKJnx
8X5E2MIj2SEprErxMmQGQkT3UobW+OaDQ7l+u27jUo0PtPawfPLGjJHsRP9i2kqA
CIny1IBXDohwaqM6yiXieSmcEU8cEGNEI85JW74k4++gAU0sYYDme8BFOMtnUMoK
GWdrXPo6idS4FLeCCNxD2EFgIyTyRyeN3Px0oONkme1nzz9FDWfBm2waRsn7GcBy
02DNHWB6/v73lP2vvKlyHlp0FFdzkog/hy5uRbCLtQf6l4EBi8LWy+vpMs/0Svnb
qSn5l6NUROO0rd/SnXlbaoZtpg3LX/Sa0rCs09o7LrlUBESphku5bDg4yOAXpLKT
p4f7LicETHxKSl4rVgDG6qxyNMdhaTUvRywv231fS6KcZhdu4i+UGTTwhZrush3C
hp0fb7fhSpEGGdlI7w5ZbT2j7koDL9By/1ql8jUY1al7/mPa44vid1T/i3gujugV
tpkjR6QtJspXKAf0m3svu2Vmlr/qP+7SPsDc748c9u5/8T+/CsCPLmkIACxhHMSM
VZGAvCwrjxbX8XiDKtZjNQOHbQsvLIu4RDse6sy7SWu+AIZxL939ybscBOuket8c
44x9k/lEmRRn6k5ziJYBdWLblhCWPcHmBCLisFljJegNFrm9wvF2z57XAFAyPmJI
JGUUhIoVeoFMdqJCk9n+EpZPWjFggCdIVWY2u8TP/lJHGAwESGIenaBJnnza5rOr
BhMCr6ZPM/YkQEr4RBJDn/Jl9q9k3/gAdBfskdfxv5WoQ8+SFTeiTsyupaskxqcE
T4nujtaa4B0DHQ8g8/jSNDYJ6UyizR+Sq4t/ZEJaSGO27dycAAC/EFMa50LwGhA7
QlEcI3o9IybQixCzEWM+no67JfUJAROZqwRRZlrcEDuRYCDLnlw19kAeuiUuYC1c
tpohhQb0cVLTg8sqA4Bvgi5WjE5DPBUA7Y2uIT7BRMfbzHBgXNKf2EcERfQgFfsR
deXw1YrDVvxSapm7QCRwpdicy03dGPacFtA1l9Mp1AXJqcDIgZ1IkeThlhpxgnRL
iwAHovUHAl/RofPjHJS5gStwond+dZNBjtJELlU+KfKFiwQVy04LN+Sikmnv1hof
tmgoCutgWrPpNTvDlP9dyp8YWIHAvr2D1OrCgIl6b2nHElVc39gXNm6aTmFTG4Mj
qTi6im50iX5m5wiqJdFREdvpIpSfKTheAep55HLYq+LT0q3hPftUWAKCfOPpHyQk
VwmvT/+3HXD+uQ9i10ORZL/d0vLH8KxaHTavnN4/VIHGc/ytNehHxZR4oeYEXf38
X8PsCpM3NX48YjXm8cRNO57RFVEpSYmK3Sue+0/54nnyb9VjZM0Or5pEHIYPgo6q
ThnOrgAFJzh1O7cgyD4fM+aBqZeCE1ZJ/MmGYCHEAFNMVArUgIxQAd9lRGgALyug
kxRDAyVfbci8PBAGAklvtHE7wk+WkXSZsO8hVdHngY7h+VKNqeXrF75FOyaQL8u2
8JnMhJRGaEDXWSOm+K16o05wC2W8ZoGMAICSW1l4Ee9A0CQTBg3FbTjQeL+vhzTq
o3rxNmWwvVv/k8sRPRY/HjqYtCpCLmAX63xCR+XS5iffxD1WI0ZAazxRazt20qs+
1HQcHKnbvdufOvmerXdSLSUs6ZJu1JeyurL0a+LL+vzX+K6BGHm/NPtviOh5P4hq
xoL+iI0LiYTrYljb0uY+GmHbqaRZ938LyxJ+dw0ItN+czhSw8vTXO9zFLRdoiftB
qW07JZgIQBfRUsypkXgdbaH0ESJmN8GBtlxEHodjZZJkxY77QdVSQTP1YSt5Cvcx
CD6GaN+4D3Zp/GwHIedrOdSagJ1KOFtBeJlCUE0zb2iuDXDXsdkKQGyJWgiCYzG3
u9McazNzG8EylpIlb58E2DvBGs3/1iSuOIpN/ApS2jBUvflaLKR/+9u1WyzhjRO/
Q485gmtSfMiGig3M4asznoOI1c7S35dKke2w2yld+jNYzkX2CWblZTTOURqpDi6G
KVHM30hys4Ag7fJmIrD2k3xSDwYVkxoGpwrKdJmbuXueV2bvNvC/8FMyQAiL9RZJ
W25x4gmrcOry4rAhg/iq8PEnivpECmGjEbTlUWBn574h/3/lsG2GPaMhkf6EPlV+
v5h3ijQ2x5oH3fGeaFu/8C5sDQO5jvd3mINpYxg+DuVO+ndZ7llsnJ75ArQEKLtm
+xcFyQFcCKcTW67876Jx6bvdqO5Hx/jN2CuHAHlURD8Iwv+071+ytL++OR48wtuJ
wEJD/NG34wMJQtqQP/kzExpPnz7S5MTzKzU3en0WKQNx2EmwMd1nIb6lHPrZXQrq
PQ/NWc/DWHxTe64Ss8ZaH/EiTxz2yJIXfBkA4QtCZz6P+apllCIsvItB86ejZRPg
Nvhqmb/nWXo+2N8790B3UZhp83Vuf5TCSU+HL3cudFROJKL5R8unAPOjVRzQo1ae
BFPyKd3/gNK1Y9Xvx1k3t6yljYqvezgI4z0QuuVgc5J4dGhJGRPLafVEKPCn5Zzv
hNGhBCvSGv8M+qmD9nIJAdugBjUQ3xgoL/8cFaNrzxJ8LdU74cF9Yyn2FlCVYVh/
wPC64TQT5CdAAPhVZ2BcF5NHCkrgDr50gpLgMRd3DwWsXpV5bCH8oRbxFY6YXPT6
s4W4d1+67bBIit7xx9TvED7NWViPb9N3Q2wNGhnJtwSyIlQCDrXpfY2MwVZy6Mo/
m2K2CeDVG7WtfotxID0t+8vaWb+6HJSbyl3EbdFzQqvn7u9EivTxSwrxhMCEIdAU
IqhjCqAR4k2iQGsUDGdjxJ1AsHCTBV1fj+pHC5G6ZFucd0JJ2qoS2RLYP83nja2e
xyu2TJXPztQEkuJglkF2iiy3Vf1OwwIKHtpSDxbwXKFLHp7D82AK1MV8BuREarTm
hALQ6L+CYHT1vBoDIijpyOUsJ4evYSTFygbs0Jedz3FxP09aOFxlA3lvRHN+2u2D
N8DjLK58bnDdby8a/1LqdVCIK7A5wj32lUaQw32dd4ZsWWFar+rXkJBhD/FN55VL
va+FP4Qe+l89epLHBGP2W6pJ3Fkjad/NrmAE3zKrUCHy815a5vk6QRY8dq69ttnc
vSdxipa8wV7LjYlfwmd8L0uPVn/XX9vAkphpbNL17/PTdQyIu2xGxCLasO+IiEbr
opeXzyaqq0uMs7dhc1Re4HipjL+yq1MGy/cUnqFf3zIucDX+MA5TvxQE9Gtk+ogP
SinnD5lsctjjokN/dYAqdhex4lu1g2MVg1q9NGzKxWCxksnFl4lbffoB9jCndhcL
Ewpcugfb8k2QXJeqNzFNftugYjJV7rCdLFTS0z80qVebG3Vz5JP7a/tRze7q9frq
S7KufCJG+2wSgXt717x2yeG3Jg9PvjfwOTNQ4U1oUH38yXt6+g8KtAslZmAcBWqT
BkItweZxGRiIOjWIAwSE4azwddMRFrRdMNJy/rj0vTNkZcTDsRafvRLmGmLRzv4X
kKIyzy55YZDH155xRzr0ZwhRR97w4zU0Y/X4YvDuV9zM1H0y1dIaquTHUdjcxeFO
qxq11CatAra2fdSsNXpytQKPh0w9B3Vt1Y6N/WkAF8rSXCYo8/V0mfux0wGWF7VT
SeK04qKTJNRBZ/bN1J7zGfi8MIGJOiwNHJntxcZPbaayEbzafYYt9PMbVS8b8TKX
TGbGq5PmNTYRyC+rQ2NyX86Pl17c1W3tcsxZyh4Wc3Q/qgxbTeteQnarGpgsR30a
Yq1TUMmMwmzZ4w1RdJffn73rqA0kv5V0FvIin/YAMbRhFSVS84WMU6ClCAwiiAT8
tIMjtm5xV8SLoKebD9OPElE1lpfz9JN0HEtguwDjtAxozVABZpOocdUjtfXXJtTI
Vi60FcQBFyIhMImisjEW9IHshgqVgv9nIMK3LFv90g0hHdJitInu60c5TYbn/xP+
Lpg+GiqvDi7Zd29HBkjKRpKukOHY29m/UQ7McTKjWS9OfylFsJB2Jvu3DIubK0NL
T1y1QC1yw7ZWGTomho0dIhDiVh8SV67OBOfFfcYjN/9hAjnPdeZp4mT08NNbHQMR
nItkmEZnKZad4NHgBocWlufGlhzfPJBHE1PikGTRG+hs2yO/zm1jE3+rx5yhzjn1
30Sop/P0JgG2KfN+3qsq6Kv/sJIbFheXuTcJfX9FfnULtF8/G6ZoKltkHhCK9zLL
a4QdHgBbWVjuKgrXGSLaegeXgbC8W1VbN0wt0QD5Sb+vTXl/g6CmS418JcPIaHgP
6sa0t0ruhOEv5Ex5jZnONVzEoPLgbvGfne8jGQv62U7xDodpPN3XWvXvQhrhX8Bm
VHDlm2apEoHdoYi07U+4kCgDuJP+U1fkr+gjefiZSNNADFsyKWyIs5ycfgxiyPjN
IINuDqtYymuSGeeBa0HdzP/52Y+uD3xErpJiwE0rE5zp561bHr8VT/gywOEUieIb
VkoO5y3ErZrwZeAecGXb9NKCBHxBsGLlra4g7zh8RxnolqRAHIqf9qAYGPEfZD/a
8v0PPO9ftn/DgcAC5Xn/sEx5tqlSKi7X2BHOSFfxpaZPplay58w31TjJmruw6M5O
Q5aoMOh93F4xcz1pH/DokYuWMAm4o2a4145lcPWh5Tu+J3aKVWz90NB2JHENWb8Q
G+bEmNpZBg5WOc41Tm1aeUvc2ZrBCNrttkdQFWnLcvpzklN+i5XYFn/AYg3VU4TH
DRmbXuLnLr1I5WxNkBwSMylrjOoRrok3b0py4g1VZ9JF2GdfIvyUErup/lVsa9eV
pOyKXntNVO5gJC/i3XjpViLjqLNOUTAqOmxEiqwHooWcwwo+5WAkgA9AVvSQm6wm
ssDXmZUOMOP/KVET6ynbY2RAkjG/JDwVBlnj5SrX13FQmjoapMX5YVrPfv0VEphA
/1jRXO0CWq7he8rUNaHBSW9OxBai9LW6T++JMVnFrBYdNBRDuM4jontJWV9xsqll
4wYBlHbMIU7PNJG+eZ6O4BingsHjZI7hvN5CGgLnIaDLBQzwFeusaBl+B4HBoVgC
hrkMRUBKGGoZOaOtW9mo/8Ev+FM3Ip2r4wNBgUW9+4d+uvN3eOAYodqoZF+8bgnk
ZHoMULlFGZGVspqG26+Y//pj9dS1x0hNDz2SsOjhZKVFEzzxFL/VOgOlkliNoQA/
SdGdHdE0I6Udq2vhY7715T0D7EbkfnU/8iibUILGelcJjaU0hlyk/JW4rdPfEgFg
a/4wAb3eYPxjmm9bTGVhraj0icUIpzM1JwGZo++f02Q7ZZ9tQr460EwqtYMhh0oZ
KVmuwE8pLD9B9PWZjv3bV1EQMzj8V6AuEswuAziehKX6q70CO/0S6eNtVIqK4BpE
vT3+5GQSFaA3wsxVvFf028zn9LKf23J7MNWTZyDj+O2YHeYw+rhv0nAzBUMBDIDf
1nO1z6PaP12huZej+bULX8ORF/fM2AXs8m+SNQYw0l2zCYeBU8qK3hIn+91le2s7
4fZWx4OqAseGFB9CNxLM/A5XNv8X4C2tJiBRJLyWAgfucSQ2akMamQMWS2nXgZna
UGSL5ZeiZwEA6Ximi8NIyKetPQwmaMsqjZGvNUuz8lNKTS/Sm56fVQLivxuxpw7G
r3Qi/B81O4u+IF3X/9XKov8nta+kuIHZCq8Mr/HblWRZE0EqPf0gpmXdngKdujSI
YC4FY+8OzhHIh1cg0jErhfXThv3G0LucqPRP2LusqWKLJft0MCImCVGr2JIBMxLU
tili0g3oJlXb6W7iwX/rN/qsAn1BIvy7OQLZBtb4CtmxrHjCzH9N9fENR7UC7v9J
RTOsO9iaGsYG5xm17pzXCEhn2afpdMMIAyz7oSSZ/UxCdQreddojKct+OzM/i/6Q
WE0oJ2kZoH6JJRr95NSNpYSL0eTx+EI+njcDmothsbyrhYCrPWtvrhdoQ9fXdNUT
yWOzu87SYv+HZssI6bQjpkLCZnM60lw3ChS2P4VlBM2LxpM/3MwWqodtGlcBHtQ7
GOdQEaGEWYSv8URe7SMy5BFIRQRUKT2wkleeOXHwDzqJsGQ2L0my+MypVz3zmw5a
Nco9eud4t10yj7srDBSqXrea31cFGM3j8xWNvyTbQHkf+AxSgOl0SKmJCUdeZ0v8
yCjkrlJQfHSF8eAQ0wG6iOt06Yhdj9IJwwemJTLnciU1MQyzZBSWsjTzhzhJ7O9D
I6m9J7fILohlwLB9djvaNQqSG9+GDwZZHyzCV79wp3bsPeuU2kdjQ3Lq6kCG6GTU
V/mnt4/1aLPKxyXke4teKT+BY1EYugGlJu4+6B1DoUrecxBv9WhSz0zqHml8ErFl
a/1759awf6UPyFprK9J2LVmYB4EZ0ir/osrOwVW8bMjWKgzd+dWkO+ty1Z3fhgiO
tPO+/6eq9Rp/CuTCNlLeZ6Fc3dLqQKQ/rLnECis+AZRX2auoWcvOCPFEUgGaTP9M
o83ejwDWrsbQhVMELNLISNHVWLYi96tRgzXvOVai9psdDLsHEAyou65/ez8pxiwU
RtMA1wQO8b80Nib7rKQw1pjNhbitV2L2XC2YV6a5xfjme8YXxUTba3DFZ9aq9Tm5
tQSdZZUMJVE4AUhYc3UqSGmr3G0UXI9MmWTiXpWoLZcy15IC5hMYRaxVfqOytspm
ALW98gy+YmiKtNyKKeMoEPDHBsw9AHtYpQV6rXgtJMxSyUXV5mFOtVI/ctCXEbKZ
FafQFNVK8zwNtuCkIruFdZWO5d3rOGpbPTmznKiloX6dS/Od7qSZTEMFEBhhiFc1
eTNu39y3kOMhH2cRyh0TvfWsp6DXSkjOXdYVgxkw90S/etcSda0uFOXOJpSW7bPW
2Fo+DFIUZ4shnIt7oUQ9CCqAtsBnLsTvlGAHSbu/w2MqfOU/Tpfg1XR6IEJr59zP
259PDQ3zg4K23EVC3IuwjROdFa7anf97iE6XEBbNDoj1kiKxs5YXeGcgJlPJlvZL
h0P6XLcaj3xNeSIvarKhobwy/LA0oX0ypKgnnUvLDW4OQd0fs5OTx0uPK5/IoAiq
qKz5X5c+u19Tdzf3zQMbIT8rZZIyqfvVhEbeuHlYefYpA0/eMrUC4kAPTnhcJav5
FcUpdqB4aAJgGOaAcZFEms85B//+Lao9J7XplfNvfqszkuuWBGcgOzFOvuqNb62R
vCBwjyq1RG5kRCLhQ44e5MIx+DX3xH43Bz2NzH0Kq3ZgGzzLKFgAt9NW/1FRya10
+gOqQCvWbob8ufNF6LMs76vCUQTbwaJCIfN98cvgk+OoiNclr7NfKqOQ/nLZ7G3l
l51M5r9eIxWanF3PXRDoNWjFZ92lA9BTGQ+iPP3EuADHg6dRrUsw8sXJ97yZnt/W
MF1Ki/TNlI1JI+CbsyYiAey9IA0t8kqp2Wm08I4wSkdM/cO3D1kI+vuKa3Vd5a9P
OT2jKA/MN8MbGbIlRfeJgzIqLsrKasaujDGgMdM+rR0YHVZ5Qgk8rVN0Xe3ivc1O
6sofLBLN2DQrIJpomQ2/e7YbAZUKHSB5h+BBZQgR1oBtSaW69/lYQTvM8eaAayBn
dmJ/6fRdSBLHJKm+UbEOOrUDdubLQW9MrAbtE6vWW/MnGLTlCk2RJm+vNh10SLwY
t22XxrvwWwtm5+np50zpyvxR0M0HWt+DpN7+flKFMbXXAYBJe8K7jrVwza6Ii5yJ
lQtav6+IjbHrDM3VeZCimVaTZlfcQTmBvrEskdY1oHrx6bnvbcGh3Py6YyBAMFQY
+AG5POH33tiTdFhP7Tx8Y8GGmG0rGuxmfX37QEY9pNDh0f78S1QzD4uwnS8lAOim
9LoA/WSY61fYG06+4WDFEnFPWvg74oZzQcCBieG3TiOR5Amuyr2JowBMFmyQfK/Q
m2P9wC6IqhDuqsy0vnxzT7o9+5NGBvEL61E/pkjpS2G00JnOZrUz7V/4NYBkPoqY
JJSUugOjtRrkPne71H+o5Gd5RTyWCASVPrI0NTErEKhArsn/PNBEH2vOvHETG6/T
Ff75QBPcI09zetABqm7DUPcR3939wVOi1YRbiTCWlgT38Gavvlm8puZg+rFR8u+2
AzFCGaI3ias/kFcWgobW5/oiOaXYw58AbULqYMbz1CAx9pT+bDx0jxSEURJpgTCZ
i/Z/7NVxrxVjAXz6VErQ8/B5Z7RkqphAQsUhn2pv74aiaD11ctj5tgKvQISK20/0
gxUJeMdv0LVlhmJWw7K1ZtdxOB+A34+Mv9+Cv8Ce/S4L8dNWRstfKv3jSDdqh81H
ekNGvw0m5GDcRVtpw6irZZKeUw/7bsARjjVUr8ggmuWvL5Ej5uS1zV96nN7uWgzw
GouizgQNBF4rV2SogtH1pmhsbpWs2+8APH81aP2d8ZWcnRSChLPAU/uReGN9Ucyq
RNT+GarA4cn297KCumZfAFpKjIsPNxD13UMkYgW3hzpYM/xR33JLzby6hsnLFZHw
F8GyL6bPkr6zr98UHUWYPAz2Nhwky9JTyQjN6sWu9vOZsDgsx4rxNRqymbVBBGlD
04Njm8VW1stL777OXzj9QQpbBUlbhZxBuNPQcQKjkqMGFoRTxrftnAJwtwSR0yr1
/w8LuWZZTgerBi1b2NurdHLK+LeFpZTwe65Fcy7qGdNAPRblztBhkaN1QKpgY2No
rXglKg4kcpXXoXa4IVZZA0Lkm/kQWTXdqt/sLYp5mhN80E6RT03EKHCz5NbPaOBl
w30qo+SMHUEdiQJpJ+T25BTwwVu3uxFW8VxQc157HSAAFjI015JSr6rFvnWyVqQK
CMSdsKXrRh4rtGaH09HY0TYspZooOcTuERSCIos6an+ShJ0t/I9b7waQxR3x7Wni
pVcIsq3fSbjB3vMu0bMAvlIN6bn5xO31BJZnm+OukXovoRpysjQ3+x+oSlVJDU5r
ma8MS5rpSqhQCcYquZokgY8qVs32BwkTtA37t5S5jd/3Y4rtYI7qNyuSxrkjn6xj
IAh93W59W5PgiUz1qTRupuAQxle5LKH7AU5UNhiK7xVV4dBjnvbsmLR+mu+NSd/B
bQX69Njpj9lgZuIGOxGaL8kw1NX/Cn0wHHMFrS08PCc8nh92CTj60CPAlInr8zy6
c9creg5PzliK5w+zyUeXg9lE4Ji0nE899TD/X6bQKOfipFfHiNshSC2igry5160s
A6Bg0HQBfSxmiyhFH2YymQ102fkTrkaa0qV6xKj6KxB9YMmeh9HTlHXzu7Q77+Rl
bcTUP6nxnWa9exB8D1FTUDdI123pA3d1d6Ps35BeqpsjRO9l6rybFhoWHaLLSZ3J
n4UCE9/rgclg0QXp+cOmWhW0qf/XAtxBZnwpKZqwhkCH6pUhIUlt2F1e8TZgeeFD
rAQ0AL9SE5PENupK0yZtZDbTd5tbC8fdGVTrW8LC6ttmaV0+88XUS1+9f/mjp61o
Nhe9evgs3bUZv3wUER91p506LHr/y3mBrm9BCzGThf4a9lWcEdRGmbTkVSxDlkIg
6S61TOY7Hw1qKKqodUGh5mpSaMv8ktjroz1OX+axrb+yQm2opsxY3937gp0HLmLo
aZ8jTpPj+ylAOItFOeyx+NzXVmM4MMMVhkaLZSPn5rz9ZgUiCCPwc1sqTZMzkqcc
C1doEFuRKE5yNgXBM0nAtqoVbkb2v90j9ZL2N9InymZRvUvYtX/qE/dslze2QCWU
1MHdHRc/fMAznV5RdfhehNYs2N42HmWyrV8qgXyTEgm8cDUhOrhlry/QRwSkbUwx
vDTMa/R6tyH6kUyIqRJrowjd4ui8uJl1zkBkqTRrhPZe9JHJC20k2rResjqZbhe+
9bzJH34TgCRjd/VxtwrSlH+HGB1rVrsWgnvKyFfcHGcJFDwFeG38uY87ZDSOtZyI
l97zeiZIkIMj2WzfL1B/F810aSddEXC18HeYS6JZOuf1L1+tjBQal+Oyt0TuL04M
K+dQQst4G/M8sAgJTzlNeXp/8rj1I1gKiDefVyqnJxYAXD4FDFKjg+O1fD42dgRB
OVenan/q3hIC/0WB1L23aG0NkBaDJ4wukfdVnWpAVyjiE77v2aiz33FbEUnjgT1w
4MZp/oKZaLVzui5WXcVI0tocjOZUX99pY02bf6LNbfLRAPnpezIYE0OzKb7xWcPY
Ut3yEo0Ovm8E3QmxqthNEudoX1716hR3dgF+5UKjwMw5GTkXsUJKVsxkWrR82udh
vnO60alpXz6rK6kwoVTD7dz2DmKgannAXbRScmyFNGzKrSNIGpNCGPKNAdxDtFDZ
7cInDQF9F3UJm/oesc+yvhhZjgpngCfNAvOgm2/aIdZ96yLptK7oNbsigYupq4v7
9FyFddW2fErj+9el6+VUv7l9YzG704YRWuxGcx1vQuhkMCxyM+w1vrJJF694NSPV
4TC/IR2pvs5BR/uyUFvVudO0vYYSRP8XTnjGzagEDlDzI3dKfSMHx2OjJSoLtDsQ
loGcm3bO4P4W5hALexc2lWD2kugx3pdiWXrZttV1/Y0gXkkvGEpqazAeXxmvd6FQ
tTAu27SEFQAjjhtgwpvBc5b9jD09yGV/+kxuVo2CL21SwStnvg9DzePrK5EGRKTy
CRrECiYIwBkHwFaqptmI/FFIugw8PEvWJfkvGJqNksbqWedgZRuPABnfePnLQ5Lb
FTFjZZ90ngd20dD2xxB+C59gB/Nprbi+uolBYuR2k8lxPLS0LN3VYDzTWe4gsXU2
gGtn/BgDjz0LFMkSCqh9NCmiy9IEHJjbyFfFoQks+pJoDG4wCeXd1O3CNwOIMDIh
suXE1v6ELSDL5BOFDC9KQNlTUOMLMhzb7BdlWq2grog3XL72JtsuJkmCc2ePk57E
cpibdTDqM1Hz0vseN/3jGv+Kten05N7p4Bg1zd3vxMweIMwhksii1e+IvkPbTDDx
WNrBYrNq9WVKFqEvUNV/Nk9a1bwWvO5/R/DtyfXTGIoeYWZrKbh4GRWkFt5FZLxk
WgAfN1AolDLOpj8er1d8S6wwyLZpj9yB7FNG+XBJ/wjnnovall58kN1kLwuv2z2L
PuY9bLc+O90WYX16F8zqHVDJihI1slAzOjBXUPw/qr8PDIOXQM5FVuOwEQnWCOR9
WcXdxagN+nBJQJQ8wnqeRTBKxA1rIPTqoa+GYjytoha5IFpLd8ax4Bc8OIfhEU3q
9SUF7hvhi7x2KALBf3IHvP1SDaKwB1tTe7Qk5CNQN8atV8wvATno3GWldaFdLcqf
RihYAsRZbajViU+Qu1poQcJuJIeCTVzyYI3ZGv8s849pG9zHmcgUC+/Fci86rNzm
8oa5ozQKmEpJgusZEk3Fi+EN7S8oRN4czygv9405gcsMdpOgkxzmp52VLQ1C2uCn
jAZujCk0AKHsP/ZWtveYTozAeuw7cu13eYW9aNaJSB66hBAgLw7kCMjHcbIF4f9H
I4Rc3QHCQgZMNJAquPvXTzu+NXl60dT3b1KDiOPFge3M60qdGP2ByWvlmsptKa17
wD3WXw4BxKuAzH6xfcqXT5Tx8iF25mHeuuDBJUobLNuZLSfTljRtNrLnsUIF3F6O
AK7SWDh5yJ7G/uovIT/THrpEDr4WnJ4hFlYpFF9+ZW40CYgOG3dm6qHrnCrbTphm
gzA8DAIuuDNXFcQ/IZOE8FgRQuZCqeKKTXsOmV07GS/HLtqQyebiwFY9Zkv6P0Dm
wVq3eAQ4w97LGVa/SSlkmL8igj4Xq9ImvUXlTUpi817v6Ga7I+hCLRGF0h8EUXBe
WWkvjwBuI/XmmYd+ku+PQpnmN1KWgxxJQ43LNmPc/LodOKIEpdFExZ/BApzcJERO
ZQb5M2cDTFKObGAMY9Y4BzGHE7eNEdgyV8gUPuom+1jp85n5/MLKOxM6KgZdZBbz
/stGEu7H9PIRCh+tf5hpMIP4FQ76mwGTDr+3VjI72hP1LIPoPUPS3P7NhL/hc0HT
QpaVL9qqm4MxbSaTAe6N532Q8ebDN3EBr4rfJHIRcAT07mXxObhvtwQ6BfSId0Bd
Uj8ARuPkEIWZzHtez8HLmpN7amUU2u1F8ARjHYnH+/fTpXj8l8oThGaf0gP+X14x
NpUusNwJKvBxdIDSXjINMe623TtU6IL0AH+fjB+rw2gIgZiUZXjWUqsgJYNTc5aL
p6k/zF7ZZrqOSt24lYOVSHl2tryTO3dcufTQn0IfPvDBpM7a4ciOF+gaaeo0AtRZ
ZRukU5KjEI4ukc9q18g/xCm2YxlsPB7OPvim0aXENh3p3fGmciAYg8apJVdoxj28
u13Bau9EcyrE4YcBW5ijRmA9dn2gHl2WEWeh0Ym8NSafrY06o34KMonROxvkz/eb
MxRvf2B9zRjtOsGmdozrxxqrJo5xeOT0KfX2PbjmEWuLg+6UmLOlf1NHVZPDmOni
MuulNZEoqAQsAMZwVfbsRtvq7Avr3FFBGY7ozRvk5Fw0OU1xo7D6QNikISfN1/3P
ht77K56+JmupkirV8UzUv7/4myzsN+Wum5MN7/oF3zp9GU1JWKGjHIIu/Q7IyoUx
hnQMw9jR32cGHNFTXhGxqJTbN+bLz111bMBdmoxDP+btPNx0iA20CFd4zy7DKNtM
LrHDUAsN+Id05mvmkTGJmdXdUlIXuzVxSY58btNmuRXeF1UqwbJ+pG+EcjBhUC+K
doYJ8fdWl70m9Z26IDZ2VY/o1J46GbAuPYYW+IhQULQ1xJ5LkK2qw7VPu9IyhQYM
uGOzMrj3OaxsyUIcYMfiM79QlAEDVsuYW84cVvPh0wg7qDiGueNMpi+P7vaZXB0v
fP2g+JEtJ4GVCUJTxhwoNvY3hc0/kusbmRVEGrSGYE6K5xHqCNu/77kQShpJ7FzK
qfK1KVJt63WICpef8X2iV/xJ0XzQUpzDHSP/MH2TbX189x+pYtO3qOh1uh6M7cxL
3SH/m2sGlE8+s+BcAVoSk7cvsaASYzLR7+2l5C/07vWgtoja+Jd0GydNHxstLgf5
58gQqVS0tHpOQ7ed6ZxxK9DC1rG/XVnJQ0hTv9fX3t+OcV5e0Y78ss+MZSPifvTB
nPAOOm2mWkSaLBWv25MzWBLFxGv8KID3OEAzZF0E/4+qdQ/BCQtZ7jsBD19q/Rmy
63o30mL8+jdJ4xAGoJy+r7Z62hIHvJ0K+vDyGQpwOaAG3YgaEYxlWUHdMAzf8jZB
ZQu+s9GCUmomA7/kFFP4cEcDt4y3EXLk2R6RJR9pjurneb4xQStMr4JvMrY9aTiC
9XtVPLKbVsXFHvF3Vy1V+f15JIdTin51RqHTowXLo6zRlhihb7NxFYPXjvKwcA8c
DNFMK3iSl7vUzdFiQKD0mucBOrejRbBRsMv4hNwzj+rgwnsVuOWW8y3yvlDKwOYT
0Pnl6ZmyWIngVFTcusTd1rr05YKQsPbRR/WIZgRpoVIV8snaLiHAnnpLsvRiHYWq
UEj8DWQhMerT3Ts51vHq7Wdtvyb4L4W9RcnrGnG5l4x3Cz3fXhRMMVwl70RtcMBf
ySS+qaEDEl8ap41/1lX98kSIMHwjen3AOGRKtVGGvRkO6dv/sTAUiHXeGQNZlpXh
XKuH6HsQXknmTCl+ELvzmpcHktlWqS+eSiL9QpY4qJfdkf3PvVZZ8du/Yaugyu+5
/nctVgcJ+OwD5SlEGoHogUmgzs9B7nBIQcE7uxIePo1fxBf+H+VBHa3ndoFr7y9W
F/OXKXtQYCRPw7PamblLrk0fxvRUA8zgYUSzgBUDZazf//HjuZz01OPkb1mBguLt
JcKzyNFHw3bVFAnbqIhIzCZyZ3yVoc3QNg3Q24TSbyUEZDGwPPyCyOfXALd/Oa/F
5KaDQyGZ9Oi9fLZ2nSVI50mTQjT/ppoDt0A+K5tAyE80bm3mGkOqxEF8jTF0JoOd
/k34541PJO2ktFMRGFicw8EjGmFJ47+LZOMmCblr7jcil31J8JeScifVyhOCYFYS
CBuo0yQOfhw/c2j3DdkEXhWbYEwtXBpo677wEsSGTpjO2R4+9KtZcw9sRonBfmKC
MAmLopDuNNfMCh/3zhPPHU68l26RUI7lz12U5DBngUu9W/BknvQ9KFAa7M/xq/lO
G3eWYf4T8f+OdZhU33e2hsdiJsTmsm+I2MCmBOZnMvdRCpx1vNcmqReTHcHxgSTo
zfKbPqkVDPHRr8Gv0LoNJit7IvWzhwGmDweitSb3JFuMMVcv3VvypxRTVPhGAQXR
YO86VunizRztUPgW7vaurq5tITqYqJL3Fj2lTmQx5cZO8EdyLlScWJLWNbC1d1vg
MQFEJcBCwD8b1Nm4qJrU5V7tNWiZgihv4XROpn6yOwxKjNooOn2NjuGMdNgUEHVx
u87llUAKYfx4wWXEETWpxzcTasb7/C6vOBJMS0maG+Yeoj6zTEiWcficN2MOiUO5
pZ2Vwg3S/RH8WniZbYZJMtEeENUf0JLyLS34C7QDxIlaPWdtAi/W5WTzebHAoPy/
0ujZNPs6295hTvmPiI/jEkFs3deq4B7eq0EuzBVj5DNpcqvBElRvHuLmrxkbjw4n
WnfXbdRm2j4RtSYrAqdzPci1cCidn4VnY5sJx+8GsuJp9VmfZ74Sg57O1h57ohmR
Io4zEvksFnrDBd7mgLlDEqdx6bzNIyaYU+EQuAPzsqmbGG2M+pANhJojJpT4qqiq
np5qnUX0XIqA++NQTNu7/QPMmYWrzxLKbn/8NQZTxSFnCyy/UiG4xUHYP+3JBxsD
24bqRw+8eIN8vF8O1780DRVpq2MRrzFFsD+WeqpUyfFFOG4xBVN2P00ubv9i/9t5
EEuTFSLTjqjii723g6ekrA2VEDUPxhMcZ71ujrmQph8jwUTuq0/SRk2x1SgMthei
Xegorj+ybGoJURe6JapZtskzo/T3d6amCriPkm5F/dClrtWSE3RrWt9wXjp/29L+
jXenQn3nLV7eC7gKaHgiVx6xJwx5gC6oTHEPVsIhh6csVBobO2ducP45jV5N1YbG
KFP/HRvv/bh6IxxHRWDXe3TAD69v+arj9MjpIENbaOaN6o6wVzZKIzWfNH+d2oGY
J1Cs/NKK/BiAcnk6kpP+DCOWYCss7k+ZdhuVBf7IUpUH4ywKMFerPPHuOIfDxoEP
grAj5DbH8aF/4bvltMec7iRa0ICfItZJMt7UfshQI45yfsiBEJ/8MuDdsw5R9jvZ
/e00j08dyY5IHfdmsvA86xzi1wfJmnRR+zSQfYEoGQAMmyXExxvXS5G5+xVAtaHA
tTjfpF2JLXY4fSeQfR647PL6k+vku/u+OtKF64RxKpKEHuPTeKxvyv4m8SWvTkRl
qHLBhdGB/F0ZWkuTJiRG9f8DcEJIzhofR37FgKYWJqaoAt2YHG4BNpjQKIv9BVmA
2SZOBI3lSUZRxq+aTiSnJ3m70wQ0NzeExDeH7lD9bzUgQhUiAWcgUEVDg3GngR6Y
pnh72BN3xyab6SP1zfcI9drPknckp2JbVRzo8xerz9RB5WTkNCgxlIOlL1vEqjcC
30SSkJxcpUDBgegsyBdIWqN7HZZO7xQAywcF19QH2yS/8CbZnYUDvkEUy5Fb3CqP
3J78lPMHBi0o8fn5pMIhGx3himzPRM7dD9V0+HDf2ZnqbXGtot9+Ma3CGbuCd9MN
f5LytFIs8n6RWw2zzL5HkZGg284zzO1j/IqrLIYGhMezqxZIYZJXwNCeVoiMePRE
mwfe4CQ87ksDfGNZ/8awdoJ76yet8TmRx/KZBbxDgRBWiztcdUGCmE/tQ68MgVW6
bbtwWDzpZkraYP1EVfzNbfhjZ7nldE1N6ubn6WRO+l9DavrQlmg2Z/u1rjKi7A+G
JHrInwCuMNndufnQcf50L5QoL9OZmzztiK1qJRhWF80AUASL4GDAUaOyJpAwswfv
miAp6nF/IkeVcd7lvcbfGtxXu8o3QOojKSrf9a0+nnNCt9c7eZgMSAdeKFzDk1hM
nefmRXi7P8MkRwzVTw4XXx+PRwMaF5qGljRvRl9fPjlrzZfo5C7i76S9Jn2Qhi8t
DLVh6R39yPPRAffIjRpAnIeASyZIWLNBb1tAqzhQnm8/MSvzIAxnSbOV2Z+HDA4S
oMKbZ/k22bXNslddgxDUr0GlL0qv5ra7k0Yhq5omkYhvyk8YSDHCMCwql/rQX4x8
2CAtpMrMthUSh5xtFshQzmBP4sMEawRvGkStRbLmEPwSxaM+GeU+60m0jhhQMTHV
bZdo7OlbKFzbyQ/aaPOoEn4UsiLaG3VoWgPga4k1jHD0Ta1Am8653L3lc/5NM8BZ
bv3o9vKrN2irZYR2DtWP3UvSc5QH4tkbKp0ryPIw1bO0/RkFvVLYZzEdNKYdXGFP
ovZ7kc2oDRClZrQUGnILrLL1HC9JvQqFsnGK2vcVf59lwGUJWkRjlATv4+lEuRJF
+WgSbxrh5qvU0OjoJEcW1boEK3x1S37hJeaaliYljBOQcmz3yrpiGhdWYl3mSxgY
QgDKSYjKFFHBNmyqNLEGBBqAW/Fgl6VGdU8564R+siGFKJVu4Lodc0xyKTJEdPmm
M0oevJ+9H4aRQcElSITXHUBCEDJdyHH7YW+ctLEnaLTvoBy5FQyx0mK8NJFOvxKf
Z+3DDWjOqfzKVjz46ald8v6fLeCg/357sCt1lxosTsDghZSpNDJw7SL+wgQDaEOA
5UNhfKf44UIojdz/GctlGmMtq5ZaCnzrhqGoYW5lklu1bD8aXduPXC4lDZ1+/Xee
sMnm4svw/l3AFf0nUCUW3epYXLPLkJvVDrcwAVLDjQgoaN26vXNcr0AXq5KZCkKp
pMIKkEROQoieonvjZ7dfh4yeehzJD8kwhZNF6A4B4ZijcIAS2/je0hHLgvsga+SI
xnSTzC0WkXzFvdjEMS/Lwc13krpIfjiMjeH2/fclS+MNHARIEtvEijlzAJzGYhPk
0CiMX4Pax1HlMPELaU7/yXVSxzR3ngzXafBmjjlsKFITkt8ko8BEt/cnNT/5e1px
S7zNEwOCfI3heJhb9Zrdd+P42PEdxKZuqkhW34dwGrVGlX84HRUaN0k4ltLYc9E5
m34Pq85/TvYxHuRECVvlTyOnfXYhfLrZuljwG7tiTGYyJjILaWZPZaU52zxTMLvV
VtrxwJO0BwJpNtaPh/rQCUOMKQr1vDn52W3ZVB9ZJj+dEI22HWyvzo6AtR8Uz4it
SI4PqUaHSrm6Zypsx3/FjuoWlZi6yqfBq2Lj54T0BBEcVC59OwxBIsMceZVCHiMH
ff0ytRm1lMlfla1GnQnqnhWUiDmc0kvoSe1qbyOyqp8YrGHU2I07wPGleMRVhP5j
5Hu1Z0fR0zaQcprxmhyRf/fpduKsCPreqmsd/a5y8vhs6fN4QRIVbF1twSp1U1kz
pHcY6UvfQ/nVbQQoTgHhf84Qu0Hljx+MGyAtUENSWEes4oi57sMP8szO8L5do9iJ
mN5VjtEJuX8DFCJUxbwwE/Rjm0gdyoTSWHzg3e3s6iReKPLM7aq0cM5VKAhiDo2Z
fk/bLdk/GTTBCZqsZYLA6VayfAjsxG4E/AgP1TjVRZNO9Gbc0e0EZnXqfTURxh+2
GslLrs71P8PZuUjszZkDIGXxnYAVc3WWp6unsMgxPp77cNdfmgshjYV4EElUx7vD
Pq7z3byyIuIxEzGuXtdNKRcKQ1wb4Y3jFAOkOjaw13gxuexsejKA/ATB10BmF30v
Y4DT96RhEkldcfi4HsoKXfCGCotoo28ocp6GpKksWv179mByI/n2XMSErcuDAWNx
2qIasHjurFhfgXhzCg8+taefxyBb/q03z1uMj+bNYrzmbxjca1SLEm6S98Z/KNUj
cTrwVb0DmHMdDRKzJJ9xdazhckdHFNlEJ/tlrvi7QO0ooWOpaI8YK6pHCAsl9+Zk
v4fGmGE824wt5PppW7d0UAQ1zD8rTF49/hZXjXoQHrUQXWxS7eRrhzYKiBnmpDZ7
Rk34Qb7kM0UFwfEwpFItH0rsmxPaKePX6uz73Qxb8zioQWi9k3k6f9eYysoEntfu
wcMtPdFNPP5MvCYdoenTzMTLUv11OEzp1R0cJE58l0MR8r3go60Zv9osQul83Hai
WLZDaGgYXxHhiIEokJ1hK1LZ/z0RcnBB2gMzLm9hl/P4Dz22agkDWlVCn5ML9cO7
Cr5bJxXK29DB7LoDqRhyseGJoFM+M3rnyc+kpqy514+Y410cxKeuDj8wn7k9SRai
UPuuEOx/bRRCeuSvoSpqq5pXHOvd7gDBV6VMqxCaljnXxC3AKxGO6t/6Xi96u3+M
KUExDTb1Uj3meYnTvJf2eboDbTO5ToVDdNtT0a6m3BJNacoNPuK4krSybulb1eCF
v2G85a1dhaJkNT4ULLkENkQqhs5jB5T3fR0t2aAMlvAXhA4woPKPBFHmGSry9DuM
qjV9nG0q+XqdXdMQbYWcIp3GJUb6DXOvndtzoXk8RkEmxPNHsE8+AIQA45nABIu0
HtYo2T/UZYunM9qAYp42EM7kYiGD78NXlV6yOQ3kKK09lvYuKKYsh99KKTHTcaGI
3oG0mmR2JGcpN14BbJnRo2m3bGzUIYw8yfUSllJbb/nyfgZrbDnGidZ3VL2INF7A
0Qu5KKaGQt+mYgbX7kLLammsFUbG9BaKhyxoWvDUTUsvreg31CpWRGF+NWF71YK1
YKErCUZn9NEZ1p08+IIaIoCaTDDtdwR7ZMTZ9GFh9HX4A+/81EJoxnS4rvhMVYTT
sm6mCQCYywsYdfJR/sGkhgzGoV7F7TfMnteS6yzviXZSDDPKf1ZMYp7T28e+OgaA
ATV7j6aUOmm9R9B6dUU8byOefdDEDB8014QsMnUGCYqZKeGwoAR5HcX7AqVNQYxI
Y0Ew5gxi48ZTv9CphrgCLoWZXGT5ivXIGXtm5kl/FRXG0BvJV2MXwsURqzBQdbjM
3+LPsfZ6F22JBXlwKpuOlfA5EdTUYptfbrYBwJA9R8sgTywFEl3z1HvrSZIEgBSR
x+Ohndz4DNsqgfigFE5F66zfmTjBZv/vZjRee2cqCuznI0Zr5Jh2pXkGUIV2/fjJ
d9xjbZ13GLWP4wVRC1HYLyRi3QpDmuHlq4Uu8lmrmykBwHoTFq9XxJiDvyE3FZrB
l7gp5DCeobNudt0ZA3i+L9WDsUsR6aEm03MyCyJfr1PZP3F8jCZD3JljPn3gGR7t
t4zTN/cDYkdczGJwHMxliBNrGMmqWK81zKNoQIg52ZarVfNM0SNu0s10rYuhm9+A
o8it+QHe998pohSM+PHSpg748wclSLrzXVhSnifnulC7+Bl896hm4CeExgqo27pJ
r0ELI19rv/Jx9CGsNUl92mH8OkBp8ZMCs2tJcHtVofy3pvYy26ydoN1Fm5Hd9I1R
C2hc6naWjOwILSnAfuUfNctvfzjEBhO+lirLbBEicNwqiWmbUXys+q58euR3FL4P
0vlj9ivSdE9ol0epPNUaC6DlFLXJE36mfZbCIIiJQtLpqX58geJvZwYC7iFnS/vo
hazPxaovkHwoZcq1H2/7Okqc/FrMCL+2Ci2zFpxeLjKQZstmYEo9KtvDwlPkNl2v
CUnY1iUpLcmNIhrhw+qtGOcTYt7NK0gynMmVBpBa8Tgbjqh4z41T5J4tZ0atdZ9a
EwffXpijnAfM0zFgy0Q9ZMVIKjsEvGRDhsoK8biz26bPZzIepnipjKMLr3S2ef1Q
AxOSBFnRZFIEIYSV6R3fy9kCTKFwN40A2jYuhQ/JyiqyWZni0w7G/IN1eTLQilUc
vxAp1K/zwai/zWk5zaL0GGSicNu6+3KCF0MQB8j+NRk7Ba/fV2g8aQj1lBavTWQf
UtO3im/zT2/Dh2f6i+3DcvWxUQGIYrz2dO2EwUpIyQuCm1VaCPAamLSZb2tZbBwy
f1qmR6QJO0GW36TUtaUFUvV9QpLs3DkC3YzoMBb4jCoaQH/qvxNfDi5k6GJ0gOr4
Hq9Ito3enU5TxFdz19dtreCrWV8cPFsLmZLOKB0dEzy4SO+oVCUbSLTkbJxMEkM7
AqVGgEOBF3C/nXdMKlqvqDHkDOdgUw8HFkA+3QoBMx5M2ZwUaLyf+YIq16VatAAZ
49AwpB9tXp2E7wbdh6RZzWPZpI59nbNAA/RhqGg7cmK31oMaogJh4QtHsQ0N5UwO
IP+bWkw7gVmL0+XjNNaBTs61KnAdbnXrLTnjB8q9OgzAnwujGeFAzXLY8125fVVF
MPIblVxxvoCT6RKoVWZdDQABECbVlCTqnTj6P4qkhiu7FXZ5hS+eaoaJrOyyTia8
RwIcZ4xxVRsNold8ZC2jipy8z/ZWfJVXvLw/WRNa7MHP4cth/paSB8h/K45efhJe
vPnQ3dEUE0LI4ZNERU+mA/ioJt55vwEQPpqjiueq93vRz4oOGkI+SRUJHvtpXLMF
FZXsolKFSwO8KRy40BV9yRkFsYVRACAoCqK9lukkrNu/bXF1cK/J74cNRoH3a+8o
L6VbSr5S2Ew9au95SskuRj49elc5W7uesq1xyAQIieg0syALWz/9B/2yQt6b6jAI
s2Nu/QvzoTsrQEpY8Vk/UZt2mk43TWc8W8mqiCHUx0iAxHXoXmiDHH6tMVWo0nA8
2w7DlfuvVUKmePpgmpaWDItMayGq8xgSocUPF8bLBzW0Sm7PBe3s7lPoq8fHYjdz
CFysB1asPxyZDWbGnWMcgozZ5mpO9zUGVCQHOAhxFNIBQZKVl5AEoMij5oF94IbY
MYkxcVyVzqbzLrGX6OGEFDnij/ioTeA0TQE4Hw/mwPw0QHZgIsRJFe31IJ0oMb4S
IQGUbNxkV77qx8z4b/6JLLEiQuCnOEXr5MzvMwdCFq6l2qp9vfTozs8LPR9ft7Lo
3jCP0eQXxz0MbA1VHkfF01YIqQQ3i7mI48kdu1p4ElUnYdMDyONPJpGWvaBLCRTE
IkJDIQOjdYkH8wYjtV5ER1KMWlmFCWB5hLLUc8zxZK4ayGe67n1yfIMss6Ik2fh0
MtyvNKjurO01NTWkCHhfsSkZhatCfnipHmOgAtTgbwg3V9ydXz8OGC0xxKAw6Qrr
5zkrd9B+68rMPB+4sU7o2mDFCcQdqQeE5t4utLYasYfhTzNnEzJ+lB+NVYbAoGXx
i595M0cuTaqm6uDomzMQr3RkLKQGUyFskmbyWZwkKD/WtA5o8abm4cBT16OljCNy
VEN2g45TUZH5aLuZ1s9PJ5MRQ85yO0q4274p+6gsRnpw3ZMqIMCNsPSjmSdNGbP3
QJgf0STm2NkPn+QcRBBA6KLPHHrEkNSicYudSNkMhv5tkrZtZw0JBPw3kN6VKbrp
iCYTLiHzct0cZF083UoTkTVwqsqXQFR9IFD1kTISV/q2+gwW/nAFb8w+i64GRM6I
0zByE++xc64Mjw/sZgSaL2T4debMuXyhxrmre7Ow9zXbsKU9iouaxa04/5HIQUkv
Ep1R7kJe6oirH2Iwt2f+E9hB9ilmh0Oc8YZvcRU65CA4DGO0b2+PwkPTW8Tu1M+3
M/Dz5bKP4cbU2odv1znqRgpEowrwOjIOqCOFvPzir9Fm6FZ3CFeYaN9GeG4INeBP
YDHqXgTz1TdHTd51NfCRC44ap2Zp4PuOoIZtpOqWMPEHbqsE9H/J9U9QZ1R9j0em
Oyuyn3itsAwfhwd6x8hmXvWf9YNPnhEapa3TrL1TK7roZgmi1dZ7n1+beVKs4Q8P
R16WRglsoYGslXTtWkoeH8zcbmCxd2BRKxuHargpfi5e4rOZUWR8++UU2Xq1K2FN
k/poDLMCJ9ZldFBboppE5Z7vpspHpH9cX6MtTmGYn9xdsE3dQtOMjg5KgFtlUS8I
Lu/uZd6MOU2NzLJ1wtN/ClhV63IH89fPtg58aS+s8PQT0Y0ClMugEbx3FJ2UIv57
yi24KGZL+65CvfvyuNSNOBYewTtI00/b92gAzN1axztbgiWLd+/7gU6LhTtlhq8R
7MpvtTwaUFQI59gKFYaOePqLT/i6raRcHhV3hRqmN/hC1Psg00rZeL9l49ggwKpT
Uf1X3BcQDU9VFz5R+iyOyG0iXqdUz+f6B8dm91/cALGWBb1ZEQIkG2sItyIOP28j
EIjlqgf/N2ixEB1RI3r1IN+czR4/AdkNidr0wmTUnsm3opa7bUvUYZXTcPl+ko86
4v+8dPWGIE8Hk9VV3+Aan5y3eYMrQtDL0BiYlh1TjgmjPwCqJu2y/DrZ7S3ci2Ms
K93NWN046sm9rDzNjHaFumit+Qnzfcp8FfGENRKrGLY5gajUhMAaGydT+YM9InIj
yh7YzVAQ49Ry6F2jo5RGz9lJp7Yo/Gpv2bF7upqEBJNqoi9nTemYe64puBU+Sgoz
OGTwRZc2EvwQtDoNP26V1GnBFCfML/W2AIWfglbVJpfVunonOifaSjBcjLkZVRbm
ERAylVxiDRsubBJVPGFCApDgiJ/V4hxOIvS/jShJobKQBmSoHCJTKBYwA11njg4Y
DoAkr3J0MCcRNYds07ubhFhhmHwIxgxrhJqVCmE8Usz9s8+N61qnmEHhmjzyRSaI
RofcCbD0DHfkQ+iDKcPd0F4SsRk3zANDeklyJwtrn3iNRyfScu3/onFH1+4YaiNP
do1h4SAgkdvlHNMeLnH3m3l1hn7YJPNFokPT/6R3yWYL1imir2QM3CQmAIT55D0E
NDIVQdy4NuD4K893eFD+VAntDQ0dBgSoJMHHj0hDzK3nqYfRWfmxjudBrt4BCsy1
TYfu5kSho3y5Tusv8KigqQRphTruLzchyRDf6z0fyludN5GO1zEvA87nHPgZGrNm
3O+UzBsi2ETK8CMXLkInHdl3Bhkk7z+rjj2JAuSyf27G8AhzSBq/RbXYqX55bWzt
Vin9c5Uv+kWz3dRD3on72cm2qzCNHuRWjoyXUmTcmRjbTUSFzGodPEPvmU5E6yDC
WRKDyw0ErISmn/I1JIadflFYoA6pbjIVaK0m/pZlw/gyqCP7IPuYkE11r+Zf/JYA
5C8xjW30RUdh6XXaEDFLnZKekTlxhvRW6UR2AsA/ZoZDPqylR0WuIvrzt82a0eF/
4ukPTUBkWBs6k8hvJ5QMnV4oWV5vDb/ipQW/SyJfvXYK6YDIDL7zkv5JhsQ8anJH
na0093A5ZJ6pa1IyMrKAlvZ27PM8zkjNKLwKsZzQzq04me88ecK5PienOVy1J4ea
ebsX+7Nz3LrEqOd5fNGFRSjRCO9FJK3mW7z/xqfDga2hRz2EsIncZ8UctA/ZTRdk
UsZ1o5AAbUwBdcTfJjtnvRBR6u/0fKrqYmSu+btXO4jzHlsIerz/0M2788jD/N6+
/tSXO6acf1feKuoi9YeNcoYpkt1yzF3qNICBgtORem+Oi34jsHLFw+k5sSHFqBj0
sQPgJntdlmq2i1uUuk+McZS+48xRpa5wgV894HZ/jBxMVIpep3NGsuZSP+fBccl3
+oIGhL5XGvQsAZ4UXKjs/5p9EnTcfJJR6QUaGQB7BzibNob/aEMbD/YLjfky55oK
IHokvfWpll+njYQDmoK87COlO3w/cnlS4pfzUziRqhbVJ/kbXP/liAgxEQs/FFDi
SPXXsaZ67eiLFZKfryWIQCmBUkN7js3yn/BUEMpiUxvVM2YnOr37+9fK8Q6tLzAG
14ERJq0Ycwqe2LZ63PMMRbRvBLEMbDvkrnWnBGyvwVCcdRcjVmDgliWJM3uWTAPf
Ax001NZ3dazJxhWg4Fxwj/cJ3ep8MNLpfXQkRZClinZKBt0pBaoKu7tjBFogAkyh
Gm8+cVVHiTrk0V4Rew4wGZ1QBdsQjBQcya0syfG176xvTpSVWnkjjLk8kI43YJXR
2pv3+1u3Qv0KD7kAE/vfdDYRtg0WFpYXU8hCysNXEdERCVgqHWJyTLgGWLkm31WP
+TJnUidWsxcxLRB022qoDpnta2G3KB30zU79X4MP+azkIOu9DI7rOfgLV+c7D9Df
yX1AqUoSUvn4AOVhfZnS7MLBy89vHjWjK8WYKygbbVepgreDMclKHfG6CD9LI048
h1tK2Nffi1FuFLhufvIOe/Iuek/2r/cD0DIxhyELXySH939a7q4CF4RpLpuhhjTN
gS6xUG/uVkJlfmkwdxekgkQk+GGu6MxHeaigfoGA08zbDsf84CXTu7gPBrTDddUY
+YHHxG+zaDzj+Hh/3fyn/dMz/dARufpvjQ825BKwqt44VlIRkq7wvYPlbiN+Oo48
JkBaA7Jr90jUB79l1ijVCrowXfIYnaa1VUSnhuv3cshaCQZYbt+StgLYJwC16imh
yUjzsF/cZ87gOfVHlInfE8UPKv4MKuDJfKEDBcv0Acba2ZWJRToWUuz8vNbC4mIT
Pm/Qt5MwZsskHyg4vJEsWiWeg8mFd5gSxDFOAv9vN65H/CLcoLGxBPSHAmW9aAM2
OsC/E5mNXHtRA7YnZmhY4lcVhrme2JcPZhVukXsupX7MRHOqjOJsa66RhzycSoJM
6IJuuQcN3X3mx9sidxh3Zr3K62uJfnFr1oz+zhq485Tj+bD0TODnfElyNhZ+MmCq
PU1KHkXpvGZlTcTigfvIzbsCUXV7IzKaIljwwi0r+0V/GOdpngbdAHQydW+i6Thy
HxeoTzf32swmuZ7MXEQw6A9mgfWWiWfY1QXp8jHMi8L0PT08N5E/DJ/XVFInzHC+
SEU/m+8sMvFgtpJcb3g7+JMfJNieza2MXhIcDRsBiVZ7TBR7pfx5Ju523of9amPP
8vhPtGGZAEQRr5F7kpE2994/MER8UWmZxMiaKpzmDYuUIWJKyUF3/D+AJ9JcWtn8
FIve0QvDzkRsTO+gThzLu2dBjWxOWp6Gzb5XcW8QJz0C3sWwPUgiQSK81bpD6XR6
UVA9cphSSUL26/EhCd8qLEJHppo11/C4B8cFCoTPOjnQUXnWMBwWGoI1NROTcbgQ
y4fLgjG3gSoSMb0RnmvA9QYy+RXOhZPl18gk17JQk10tC6a6oUsWlwdFRbbgi8r5
bpH6zikUMZYrez0WZih5ANz8hDdUUVQwAmLGf0+AfIwSQjFTtrrsnjeVQOsh+Izd
hJi58AAHiKpjPYsa/WuCsIMS1pPKVfDygzxPiyNlUZlmTltYD+4fqIG9sQ5rF56Z
fX143d6BtjwqbuqPWACLH4ONMNnKwMwj1HkJcZ0EN9bT8ivIlY5NXNIG0UNcNDvF
2s7APNYUtwS4FP7l+kYUqMHENyu90ZDEx1H8DVcn9TSfeaI/Yy8oilZgj19CK9gB
MvPw94yzXZ86Twz60zzHEOQLfslScrdFBYIOQ7Mluxb1BdMR+PpwnjgNBr6abx87
yge0P8ZSTKit9yo+nNkfxUbGY9hVioNT5IohHIaw6XFIMCARCF8mD0lAoD2zdi7c
i3viItHBjdi7JY68+mRsI0e9em+lQ2s0RlCxffnQzYHm50J2s2Mx9mHYucIM9pdd
ZQN9VDwDDPk5WvhZPVMsBH8L7Xt/v5yFV1j3Id2CBh10E3xXuVrRXIYXdtJHQdRD
/gWwMQdh9jtK0eg7QhvHuMaAEOdMNmu8nSH/izuIy3uK2+E8RxSqiRhoPRf5MV6G
ENPJfTUHK2uZFpDIEzVLa3VxC4NVhlIjGqDqjsnSm1uU0niO7vWVdQDQsIgnkXJK
WlS4z7onF/aKkQ8E+CGhTvzJuCasPHiKaBuadM2EGhZ7pR39WgJMWVftfwoPuSPY
EKD6Y/4eY/zmcraQHuPvkQsk+2i3AyVbJ4vhrzqCW/KTvt392ybpFS8A5KK100+9
6aOeRu1u61otOngb5XHfLmIK2mfti/wuDtf0ttG8CgCa7IgMh+XiupZ/iheHjiN3
ffDxQPRcccKGAj5h/cAtirn+9aG2EHgvwUrQ1Pc7kMUIc9uTZqGdOvv5AUiA+Hwb
M3fNbSMmJwKCa84V24NNxXAWvs2JGm28Se5oUDaF2Ox7eQPjBYVXS75GTikdFdnN
lor84v4PzjNGM+Oc3hHKvIoWnUA0zJENRU58rg6LFYpFzsZ9mVHVUmG/j7AyTbCz
BuRNpzpXQUicUTG+4j5XTYOd4LA9a689oP/9DsHdC9nUQyds8gNHXYmCzlpZIbra
h94BDJG0txg6d1bklPR9AkLCXiUcuWgngXDGrPwY4Kp63aZ7RgdoC7hfFJlnDTqq
7mnJO8jSnGxtcDctkWX+Zci5iU8TpB3Ec3elIfXgqL5QLo+6DiGAUTcaICkw2p8I
NWsR69PI9sSDV525EfuAk7WzatnLVM0bstCoD1EHM4OTMcHBFB5miPVIFEJWtMwE
7xQTHXB1IxyyJdo+SaApJouhS55WDCpmL7uIB7+948stCTrxPFMxmcDWTJ9w7pyL
FQdODcgaXGhnN/6xfWsda/zeHWaWtIkfgAMyRZkkDrF3YJvlcNzs+snSFKf1wPQV
G73XN7tbNTSKTV9nGWBjoW+zfEj+VepC9V+WISCXF8KzzxfS3Gd5nCfEs8hsrm/r
x0GGOQGZ53Vqn89QyvoxkneA9BjARxD4xQS9dEUdVZvu16RfHHrovZgA7hke7WIo
o1bD7hTQ4j3pRZQaNcfokLbkWxPtRiZqvqqVoPTmJY6f0x+ekNp+zFJqqmmDzHkv
YS4HAhLHKIlvnYxnkKCygt1EBVx1k0nksG9upgBIynDjV0BIv6PEvQhZcrxTz49e
xTmhKzB3J3P+WqMDJN2XyRok23FpHkVMYxNAuAxfVC9zzHWjFCCawURNTwYxKAyE
b/2mX/QP5+ED5kA005eV97z6PNjuXjn7/tv4NSPexgL4z4TVXA7yi5lIOQry1mIN
vruuCLTU3KCOQqlWFUjXrsIEhM9A/wJYWJgLriQaQAnQCd4QM7CEecnkzIHuDe5/
KlP/4kAXTz/17lSjYqiYWZb/nRF6LxK1QsQv1ABfe38Ap2z4SxL1tGiQvhI67it8
QJDbmSPmU9pnkYoP+jaisV3tmsh3Lp9AoqAyfzphUl3EshimVSxVQ0PU6cbTrtAk
dFuHh1lYLU0TUj5czy90B8qhnJOFCCvV7INcqEG5ai19sz8MQip09wKBPBEyMttT
otWkXGnOXCoWSyq1FvjM1KyP/F5Bs7tJgeU6ycddZdn2UmsVf9evM8GmJ5RCgQg5
bAzh1TcJH94ZgA/C592cUzmWcguc1ke3ZTB+TVfSPfy5hpefEoO8k2cL4yDLRajQ
2W9efCqLSGA3oVtGby8haNan0SaYdaaL3Lhd8l+6pHyr0SCemQ5gbTJDAYVZ4O2y
iUi/URh0icO0WATqiswlbZoOy//lt1dFt7vEy2wbSajaMjCzwhpW7kbfpQ86o52J
9MBZHsPggHm26NiO3tassJwp5EaSr6BCb7t0N9KW18aXFXMyNHHKJPQkM95hrTyB
1daowHMpnVkotwN3uIi88yzOBkUz0pdeX4otaaRr3AIV0m43ivAjTMbISLlq8dkr
2p1p924P8PvXjPfAQayoYBG8igsLiqSvLgevD2fLJa+GrVKmZKiNT4uqQ/61BjwQ
dVHN0EXS7bpeXmvCwUy0vzGxr9s1u4QvwJHYiw+Kw/A3sJE2nDE4MqvaoCME5yEv
EN0umH3Rmv3YjYI6v7hfLy40tHkUHaMqaJmGkdPzi+3pFvrT33S7cZTbRrQCZ9R2
wBlkQf5ZJsxFSOgCk5LLWlzc4rdmLROTwqNR+eSPxdJYkMz6We2MwX27YqH5kSTR
AoqN1dCTY6z0++mzfAU2ZvAg9aSLHNxJKZbRkZ2H1W8FI9Foe8clp2Stwbje+6pk
c6JDlvO9eb3FWmYC/c8ZsAJN4aeYhzeTcUWJrUqED2RqPbsFZCKqBwpZ7Cx2UY8h
9jYTpgVlhAH4LBO8MQw5xKVCGmJth5cD4c4oWl3jpcrgQ/KWBQnLTia8bZYdVfu5
CdY6EAKxY4+KD9piChDJaU4GJBwlilxbZ4sz83+yB9felfG/qyu0uakXSaC07hV8
svVSJghoEehvdchu8tkZDyga1tVDqu/gn4lVYWtwhyCxya8EtPAFnkrbztKEfiUv
yOF6Y6X0NBLhq/4x+vzCPBlAHWw6xHpEEY2l7NTkj34D/Ps7ixCB2YSMRgNdwZa3
k3PM5Ihc8UZ/eNCTHfZ7OkEXwG6zPySMy+o3t5J8XNCC0sN9lxaZSfAC06irTstN
KCpQVoMlhBjlzcmuqOHANqEe2oq7u5M5BXMf0/rZdRXtw05xPNZPpwFWaB+ukNBN
WjOJ+mimIG956H1Wne/vxVG9Pw3FhMXfoiXXBt2CH9PbOFH3RWdMCD/VxC8bbudb
cN1EdReGofnlJle/4ZnoDg9vAnK+sNc48PnKIdsMR0Rm4nefjMobHPzl4S/NqLJC
lcaIpxIr4weUyYB0F6sf+cVMtIV4fUzyqhfFQQrsIHuIYvkRWVlIcA96q1d6ceEm
FSoU5fJu+aLkxf6uAopBg9na+Pb6qL8mlT1aUQXxjejcTYpf2xopgGBS2cUUHpp5
UEB+5LsbiseLpMwNJLj5KvkR+eSsNGAVyRCHNeGcOnIQqYEO5ggW+ek6ixnEfcm9
NnLLrW5DSJ0l/lTuhqmvrDbtblNvCCK/PMXqgsagWK4nuA+BJXY38xFwznFROP14
D6CwY3DcuyDtQ1JAQoaYApbC18A7BBWxJtGib9kS2yU7UUFutyhEJp1SU3V6wOpq
3OdHntqt3r2tTkls+itZp04Yq+bqJC9/eAuGZIK4Ty5aHxG5bJdJz23PyeTQcua4
J/8zp4UjVVgdeO6xphvpfBHYKedcnvBNdSkmYyDGD+2bbqcyggwXpe7oYA2t5J3i
bwkUkEFgv5+I7i/RTyyrB81aP+wuIFeeXVDwBBomshSBotzxJZjyGvA8zNsMIpAS
MzlLvv6uVsSGzpIP4zcZ1ZiH5xJdOhzKHWHoniFcauPogvo6BByeIjaHRlr303er
8lFLmtywVQ6a5Cn2/Ue3vf/xEFwVFn9JPRFE1J4JJIuShS+r3vhZylst69hSHQxS
ujCSlMLw+G6eYBKiFjj68b1d/YDQaexPVnR73sr9Ty4Cl+o0QxbAwfWd9Yyeeti8
xSTGO3yNadDR0lt5W4U1elL3D7uFaPmL0qAgDCsC2j/ug31OxIsV6/V3ZWKkTOBR
DylOYeXrtElrxF+DTWoITIAFcO3ziwm4Ds/bTnmka72uxZ129BrULBsStaojZDNZ
JvNL8NTB8Oek+8zpQSzaT7FNch2Gc5iHezkCdxbp4M8QxwKncCa9XfJxxHxdLB+9
ocu4L4xMupR5BsHBuCBXkaFBbqvBVeSu+wf5UujDlbb4+FKqqIlyyeJh/um8Q7Af
X4htu2TMPLoko2BoKOlnXaC3gFo7nmkDm3wx0cb80KkPPLWsW2NtaFa/YAFcIocg
XxfhOkLAgf5f9Msfyn3nuC20LsnnwNCYG+0a4reLU3sL00FzuByfdYuE3EB5otJq
iAzzqwB6UEjQ4l1OrJTk2h2hR9m4mdy2PQkKtrlmWg46+VO3ln0P7hWq/I0aqM7r
gCsduK3/wt5k6Om+7ZNxNftiTOnBpIACdb/QwW5Caoy6f0ocTbJ4m4IuVOVd6wG6
geRa1JZld7uH+1nlSyMv6Fr8x65ADUd6Z7CTkB2bJUbsG+vnzyvUI4/T2gtphh5T
0Rf7vHUfWZCCfG0yUIo+aF/j7ZC6HtSuoWMKiCYiNHVVcxPJRimrvYpcU/KIw9oZ
rFBDyUFOV6VPv686Wd7xoKmkAt/yoOe4RJ/TLhIUdYWiaY9EciU3VbLtHS/D6FP7
e6KVXl0+iWWhEx5n48JU0yyYNMaDED4RC0KR43+Mxhxd533KC2/5SGot1cFSQS3t
rztUhCqMpTcvroRKnyYvOVteSn4+cu8I69swtanc4C82RJucEZOjftZSgHB4ZH3c
380TYwgZEyYHJLzCyMDpy18HUDxxfS+shKWhuZCYywLywcvjUhCTR6boVf2BwVxv
MaLpsWpBcl+FN8dU0XYfp119WdZIcTEhM6xPgJLrxcyh9u6FVt2IhaEVHenSxsof
v3FJbaNoKcNKr/VESDka+pVFPj0a3qBOmjcMfjjKauaJkJuosUqF0DxYR0QKAQj/
4Nn3rrLSVDigyFoRoUDBYN5RfFYCcNpYu2iA4MEOKgmfm2GzQY2h2+qYcPF3YUib
Joq1sacKhlm8gswxJ4/JisyOX5oN3xfW/2GCkI239hXb/auGHB43wLrNa8sFXBqi
DtDyw3EvGlzsMNGHrYMlCs4lLPtdC0qIpzzA4LfTytTWfnTv0FHgqPpAxG2McR5k
x4U7dJb9i4bhrKvX/IqQhFk7BkmgmGDysnbcrIzIE5oL5+0xtWl5UTptJD/xdGuy
p5iDuM9Ztkdvi12Mxvk/p4Dcr/qlGBBbHwZo+6K3u33E84pdJ/GiUblVdNOWEx7p
Z4PwSzN4BoJ2bNjWOXODe6ouBnq+3wnqjmJBWonlMhBiysLzZcHwQxbvTiakmRWE
vlSgX5tT56ChNTwc6cbQ3JIvhCt3vjqLtXpU92tdBeYWl1zEKlhNe8tEaeH6xiWF
LjW2wYvHeiQ5F82GViWWTaPWHrIX1i8QWCKvmhgvpiXctMkG1gF77nYJWuTwAaPl
Oyaoc4OjQUYVa12gF6SAJYnNnPsZ+JjcaJ0G3/LUH+X9XbbpNUYCQDPJ+A5vCAYq
TYBCntmUwZFyeFH9BXljyck3/m9UTRlJ7Vd54SKGhU5SKnWN7zTT+QJ/tzbDyH+g
oPfCDO/HBA6TsdtQp5R/DEo06Y6TmEyFeHyEvw/mxIPAt600Bmi3qDmFt2mgVCKL
mmZegxN5FOxzaFdasdY09U6s+iQqyJHijhzAycslkJjRkZCqjk74X53yGRxnHcws
UVuapSgIU212d0BB2xOOT0ngETN3Nj08q3plKYWFjaqfhKucrK6QchdLkuEuZ7HB
WAufOmLklXx0pSWwL9HZSgMIyw/yEwh9/Wt3G7MEmUYh8gpPImYcon5v7qZ0wcXY
NWlFr+ypOVcIPV7n8jQ7C9WTbF/Qpm/Ny9Ee2ZCPmePnkTyWwBYwNohju9VVakK7
/PnMsJerZ7d1rcI4ih03/JSb3XV54Li1WHfGnmxY4hJKwOlfCzmGjhP7JWyz8+mj
C+8t9Nc3Px5COrFTpE5af/5qdES3PC1v0MgiY0PH36SKtw9pS6++3eLrR8z+Me8l
onn7z6KI0uD8egNcpONxWO2CfsAxFloKHTIATApL6zzhY/Dw/EZDAXks/PckxgvW
raTZ2LKYK0Eit1fhN/ZmZBvlqO1GrZ10vsq2c1LPYx08D9WQ0yFi/HOgv/PfPvOC
H5yNLPfAM0jneS9dDet8vA7AgJ1RR9N66Y+b6+dBENVTPb5Z6WTuEYx+c1RZghfi
AbouEqX/bNvJefFs+vqsD/hlz2+f0jJsD0KPC/VxbeTSaWedXR3H0NLZFlWisDZq
5mJhMVKRDsYONMdRXYt/U6BA7KnJKHtj/oMjZtSCGushXWhlaK6pYaaQTESxV+gA
lPjSzxCO2gixtBwHSM2bLpvJC8jDjbK8D68O9cTRL5FWmE6zznKmHENDo0njcw/5
z1Z96vbc6EVSNbqU0IkdXraj2AI/7bF599YOs2Gz+8/CpUgBJAHn8nwPpFzcF23W
2eLyg43+5Z3Sy+SsTHtiL4Ifhp7SQL1weLZmg+u8J0um0pZvyZCiOX0vPI3131v2
PDudG6QfmA5wpR5NCFMvAUMfLxwdypYSKVkXZYdgZBNgNrdRROefiJb32afZE/IO
a94VfqpZ6j8EL/BOZwJLphwovXpWdhReMmhQYs8gnS6RhpdhhSfj5g2rpUpxBvIS
qgkcxYgMHk4UZlxaM5tosEPy2S7AhvJvzak2dq0FlS6T5w3QxOQ8bKQlh9KP3ibX
WrBNG2DbAkF6CBl6XqOr0CBpWibbPs0FFmTR9skJ16CALCeEeYEH+2YKTXR1F6/J
ewKGt3EmW/dC6ORXyX8SMMXNofh2uz2Q2PiN65cdi4LFPydHRhdXGlri6TzkUvgE
r7fiCVS9WhQAJkEZSrMREhRhuvh7T8Md5DM1EnZXmeM+V8EovxA9kspYRga0LnFm
Zkg5k4LTTPCLW7SEX+DU6IkqlhVfnn4EKMHCNcRQkEqcc75LLhSG60sD5c4INEqJ
mIFA5nXD+FRhQ6eRcJwMbzi2fYWm9WEJhUSzzK99GRIWkyivlxoOI0+Nbcnb0IsF
cljTO71kZaqXKXtCTJf0mXtLA0A2YH4IiGDQO8n2v1DYedRM8hLQneNjI2JjVEZj
82JSTmVIED9W1++HH3gXKnnve7yEGPjxIeSmktDmPZkR7Ijo1h0KifkwM5GDpt0v
ZSwk7evWfmR9tCRvKGuxzxS07q3Wz/cuJ9Kvv/u78x6fur2S540+1e+GTcRN6H53
7ss3ByLQKrNrkQ6rXpZmfW96gh4lmkgoS/gZr2ZRUxzRT6Hp3VtwPLTP2I1hgdfF
A/u7ZDxvcD8m9O2ZzTRstHC4q2JzRcVJsjZr/H+rYvAKJpNugjbGYBmInIrJz4xY
rOsLF4nibM7jLcxWPmYXcBb39Pv00ALuAwZmKbC4ywjcwUb+Nr58ZfAiDIt2qI7u
re23jQneb45HKluABORImDhQfvQVmUcKP1OTe+gXohlhmvKzz4wUmwhq0FPA2Ul9
o9sDIjNpAI6+/WprtO/M18g6hwnD2hPOJL+Gga2MgQ+TiFwAjD2YSSwKD4B6c3+u
lNEs9zQqEXxabFR0ps/1JWguUoGJ84ySc01MbHK2jCUhESri5veAD+lpfG1U6tpZ
EIyOp1zQ4Y0HjzNhbvRXBZdDlV3LfLRbI6WrVkVufXzBRqs16GbjhBw8M4GQ8pVd
7AFj8gSLu6at/EVkDNPgCfsm74rou5YC8CbugMwgi54g/Lgxwlw5GvxddUTScaRN
nDWnxSTwTJZZNXoKyRPAJwruOlnY2qPGvo3z6DTCVV8gWlch3YCJAQNuchC7icMP
EeuUbQ4p0qkPtCPn7bFZjLA+dGM+KWJdzejj/Cl6smEhSOIbeV2KhLVCxvDjp+7q
yJkoMuOVEHJ9776NwWsdsdaniI0VdKajr+RpFOpDhLrMaeUEB5Vt5vSnEiM3EmyA
Q36WmZIV8438pnucFufydurupRphkNVPOQdgvYa3mjrKHMcJgEFbRhtbXR84tFpq
Y6mpVxQkRQXiqN4sa7alL7VjwdLoKqbSbkrFuXz2j3f01LhoZDx6HRD39gkFZEbn
Iz1xnj7hcKAuxVmfmiuD+ed0l4eUz9E7exMLSEzAGA+DPZToRAhOZ0h/0SL6aQvE
5wUSf1U67DGPnVoG7/u+eYlF2RErTwhpqLpA5mnxDUTMh5EyRjSaVfc8XnnIViOk
HiaYgzNZoZrJXrr6bDK4NJkQh/FFK3PxE1gmJDfd9Eb0FqpSgEbhaSHjcdS8qtYm
WZqKTmWhOPN+yWNRUweE4L54znZP+N/ffwfOmVabWjtLiVmpOPCpvP2oApSRwNUY
cgjEBfnI/Wsl/GjT+A333y/ILXc7OE0clo6M1E5ZjcCEMcoOXNBFHPixgnzFM3og
zoV89WvFyiNAK9I23ROGfyYE4uz91jhz3pFRGBKQTOey4fXeLgEwiy8wjpg72FVj
6PdEv2KnCMucQb3iX/X6+oiEV9xzi2vhfomVVynaUyUkxFpGFZwBRoc0f8omkkt6
7hpS4qaOPru9JHCAkWi/bMtrswBOnISBJLImRQERxJ4Sk+rRXi5AapXZYuCNPM4Q
5SJZXOx+AdBUjnWCnCVdfSwQUEQ8e2HLS2TnXl/iaHe41BeDgDMuycNAsAdWe9K6
G2l0M5052FWfHmmfKrN9nr/nsf67Yz5ULvCk3zcFNf1PvbK8tngOKf3y+p22Jw4q
4fp2JffBQMAPz8TI0pxzIMeti3xf/09jWb8Xw++x/3LgNbmPBKDe48wShSZnTdgY
9dIzyrOkKOB/sUaup3LF5f4HjdaG+7ulbSnuYSXkoqSbRI+hqnxErqIrW5ZUsLH3
z+uNUdYgMHPg09in/TAKM51rVvAI8keTCw1TExhDowd65ciniC5TFEmD2VrykeXQ
rMHOr6rJhSuqjYhRClLEfa8xfPZjKVM4KE9rSDkG2koRsyQQtmWZ3K93XDeLzfzT
Pbv0QZtxWgSHVSwJDifwtyqw58IiYmPodpr0h7pNKj2692xyVhLHg4cIZmyHfa+0
2+PY0tA0aeEIzchKo+Edb6KAXe1MTo0AUjOKEm5UuGSKmbN+p4liavOEedUEfHTA
OvaLaROZ75N0DYJEZxAX2pVx/Jazly5Pu1nQ34RyQZze75UJy81A0VcAu7r/94EQ
9gQ8a/cFDWPXPPOXNH06BNNz0hi38IvBBSZM8uoXxOh3FcRBvgv9vZ9/QEE3+ize
5PfyCIZIwtR/g6Z8+Bhh1b1G7+L0HXiz5THBx8VNi5OtVoI1fwaRRNKnfpfepbDo
PQ6LAF/XBGJCPrNMRePOH4WRxul2CjqpLjDIQ+xTF4/FfQcYZCsBKdExfZyLIN0r
kmK45m4/K9Eg/BiHLPcKUsuuB18Qhb0VH6IgJPOE+aLYSDbcwPvYTSjaMCh6OGqb
o3YrWs48Pas8haKZ6dSOwTop7qWvZCLALjhfDHYQ0nJF6vLToQZI/Ws0l4fX1wE1
rNdtrIHqGfC4c1hVkYFEfej7Iatsf3okDguAzVO7P6H3TrBh0cuEGr5qXAYlGL/x
lnCzAdcLGCHBfC9YcjvSvL5n+OMxpzv+3LiPUsFVkh2aTnBo1YOr89L0Z87Zirk/
u7W4PHDIxnhJqaKORyM9kH6jx9YOI/Ma5Wdd5Hqh//6HLJSuh++6P1TYZtUzRNbU
5umM2MKiWTaZgd7Kdh3eTZDXT3decWBusVTCBu/w215AybYLQvDsFPaxetlaGfR8
2+qlXEQZk2HybBOAbw+q3Uu/Ir6lNmCEM58Sisv4aW7kMCRxcmmNtSCnlj2xtDJ3
FC71XzJz58cOTjjldkWHQ1avQ/qVQnqP5VK1P7D1kYIO26nPqTH1fvtC4LjY0FXM
nLVsN/vYu6vmlqDra04O6DI0XIJQRO/G+oFKMApdAYdhb73s4sQe6Lbd1joZOQah
6Ft+DA/OkAi5/kJ5JFcOvMZ8JT+9qXInAECrFlxQuJyUFJap1jjacKtqqcGzxTng
UoaBV4X2HXD7BTbdbhX1a5qsBRwKTdB1Knzp6P54Ub61NKZJf8aK3pSj31nauo48
kMRiYDBWGYMT/e+2w/DRY86mGlwqVMZKI2bSlwZvSTkF7ymtY1f898q2GoMfjxDb
eV/U3pkW1wZb/WbOhPxC4G6TgehALHxM0w7QXrp3dFR45x7ugYV4Fh5EhcXg86gK
ljAaQLzcB64AzCILdDEU9YJaRJNcyG2bS1/UkxQXZSSFSIC48HN2CGPUmoJQ6/nU
gpAx7LjRLA6XLE16F48pSuYHgh1ooj/v9zqUgyI6lQVCOlBvHmGfd+XCftpAx5+K
7UP/Z8qmbRyjmDCq8J5p35p0iNyR0FSN6bKF66pPmdTLDa9wZ2wgWkkhbBzfQOKq
DXZT2xOHUtGBWT5w+k8nb1srTY/PB7MnyIX3o98EYIcfaYxm0jrc+iwCzEXxNnh7
zhBopaqHjLU1M4MtD7ceM70VoOyhZR5HGTHeitegMhQjnrXH8A8FeNGH/oWgEXQO
U/XnGSkbL/19NrUt1XqKObQS1O0BHgoe73d/vh18G9/nDD2/cpDsmWHLkkLcVoy6
gJLQuO3wYInxTPeAkPyLAHHIW7CnCdrVHZq20LG73SNt8FavDVoFhiki6jyBzU1l
0qz4DL4eMx8klytFQgD4lZ5uFtmeP2dyzR4Yfqsgq7tf1lpkEG4fSgQec3Wb0eFz
urLLcIwnm6teM1rdlQ3UpIIZGguypBmDJa89JDw/OjB49HMdNK6B7MQa1xpm6CL4
DwLlv6cxPVYWhUShZwgybQMp/a5UcAIKxwJlE7PBm1hHDIV+MYjGTObMJhSYTrUK
PStU3+wlMWoIQjwwxjkBeyxkEc21S8jlX8q+u8q2yeSpOu/PtMiC23fGzUoskNTj
UhCOPhwz9fo0bKBG3pPElHz+qBAxj0plzla02Mx+kV9pmlj/hDm/aS0jHVJHezjl
x+4OSlynVqzziNxa88Q8cmZK5VBPCNSC8+4hYqkHy/AtKi3Ak7eHGTITCnsOfgyv
yLM42J/TlQoqGLTK3/X8g7sMP5VVJzbAcjMsssI8cjNUJnwrvJqOgE4qloZfvSTt
XepwQDNrnCHfOsTRJoxwyVC9p/QOWv47OjSI+emx2aFwxdZO/2JW/ruumNb6sfJq
/xhwHhRUWJmtxETl7noeIq2uCYMx35cTGOmmfvacEWZ+qCMRf1jRzU6fSKmnMfUQ
+DU4k8I6O490885BvE1Tf+b9/yL4uvk2LEio7VMZpP1y1CaQR33L9CMnlgR6hu+u
qswzrIPcUHAX0XZh4DqEPvnSnLeLJY/7N/g/osudVCi05mo/ITYMW1ysagj09WbD
0np/x3vR/ahPIUyj3HiJK6rTTXKEEYqhCP8pClpEl0mofFRESA8r0MyagfQ3/Ps9
O8h9aTUq8QSP4hFbNMb/nfW/pejAUQHQmWsrBvWE7OGlp56+1fTwGFqomGHGU+uD
ASC/Kmkud3bkYYhHrfyD00XNuJCs3UAgOS70t7eY5dlqyjhlLRc/fI0F9jT3tapw
U346Mdh3LzPnO5F4t3WUaGysmK11CcaVcxdo3Hevhe3addMTTC22m+P/KbQDiNTz
Owwnh3TSYsaRPe9CRa2z0XZFKU9IVN3IU+rWGfYaYGfvP6nALrNYrCplQhtW4NOV
OVV/EjlIb8WT9wMAtggz12HGRquQtCYKj2PK3WhrC/HqcN5+F7R3wfHM3JPMQwgn
uum2I8IbbjcaPrz0vcFQGy5k+L57bby/Jqt1fLg2yiMrGgO58bTJmhqHTneZ2BsR
qXF/C9jmChGSsQN0U2JDyhTLrk1AhVP5coNA6EoPNaR0jc5KIXI0ghcJ6/P8xGS4
Fhd6kJ5UwUzV3148apyLVK1KvN0/gmzHV4klPGI/wtN949wMCEtqdlsBFtfImD05
El4vI/2tPMg+eAeZ4m0NkeN5wZkqA6eBalOBcqbq9qihE/ZtK7QQ5aLGZRL0R303
gT7yYOOjYDrM2oGUFw8vVq39IHss8tdm2x2DoahHlYSmReb0MIQK8pTuRchNajLG
WWuEF7g9608vtvWGhNAGf4uMPdw/giP6rej0GyNL5LT5/UbTh2sILpEpen2cgfHw
UeHIAJ6MnuhnPvjq+og3cnn6zqh1oXGs1v7UPZyEQKrebBA5VrNORsNv1TJ2F7c1
Ci+YYMF/207iVoO/oF3MTStQXR52H+PvhWhaYXGTQVUOFc6lbIPWTuM7cNpnEnVp
VrIfB6U/xfDWc+8ZSj7z2JqUGRy1rVhMFN2OzOt/Mo/QYm4exmpVAYUqUUMwPqQQ
myPkKEE8MhnEiw5CVMiI/ozEdKG7ccMkKUz1T5iqY+CQhCeso3vxKvbRuLOamfkV
stZ1VdbG9eys2pdz8RhpYatnQfEUMtHW7XMB4QZg+pcXKEsx1+/T3AHL7Bw9zl30
or5vcMSspOoKwWnCGC2MmS+SP//5cpb4kkNextbi8HbOewnz4XvCnSznsdV+SlV4
Qz7F4g+dx74gf4hcaHDdycVgzbwiq2mkmGckYUIHP+rcMzGvAxiC3VXOUbSwz4sc
gPPM9nverrqgn3LmUZswYMPqcYm1NPnCalL3YKza2Ip6fD7NaLTyjsfFwZzwlx72
hh30ubU/C8UwrlZzotZ8p/ZVhXlyNVwcLGGIBPVVSs4mN85xQ3i1xJMoasha/sU9
liIUCaS4US5DiQQQOZEHczOXjrBHkxZGMvE+q9Gr2l7Igel00atUWhe3+IGBdb8X
MovVjnAzjEz/+LkyxxNLfwxM1ROLiECws0Uk9r+EscA1ybrQRRzsH4RshX1C0bc+
fH8rMfLcneAdJ2vwytHpe54FebJVVbWT+EZTIHNUAUlC+nYSZxI5PBcPmQbMhqe6
hcPYyVYwif1gzroN/VNR5YD3PsFQ9BAKlE4+VzTagz/nSugnR9bPm10ATBgiiWQc
uZa171Zt+YcVdtWrMPyOBNcA0DdSq7TxtZbuCJ/K6xSebEyZlNByUoFDMZg1i/e7
tn3GeyROylG/JP0BHAmB7CBjkqivTT++NH1wdnBtyz1OT5UaJitCvos4Kd3PJ9IW
7rAxgEwFBE/r5BDgRHgLCREKMyrQytJxeV5Ict0U6FQIOZuBQuoC4SKYUiNkZiuQ
knvgFAy/hB/FfL0vqfANxIj+ReSXzd6/gqjwv9etgLnFWBzFWLskvY0+bLFt6nT6
A8ii6FCkBJOXysJofXijSqjE/QYtBtivMlGwXgVmHDCnaCdMPLsCgfykSItO/zgO
YWUwbexNXxkZYtPSpicE5EnIB/sKmU7iTiFTPLvw8EgSLjihz+odzbVjQ5BFeT4f
pVIrxyXT8he0vzuEmCUsqH0h/NKDkKWuULlSzOkeYddYjyV7AqV83x+vhft3/59P
oZlypy2hVlxUf1bI9LBrFeUmkIVsP4QWiV4YysQUNGZfYiy8wqe8zyHFCQd7enc6
2V2t+bu1ACD/0oKmPEbWTWBkvAMcVT8fvOkDlv1ojwLtGHxz1rdHMX+W9AYqUiwi
ZoT6OslIlVDL+A9ACG8JraEIH31hIkRJYAJVuM23mHq+W7Nqqxw4gfXn7sk34rQT
evyV0ptN1Bbp/ckpSNFwN6bN8xvjg3FfPkkVCsSY5eUAS2HjnuZsG4vLJ6F1pi20
c9j+pFMiY0IUikKzlPhAOE4B4RrRFXC0nA8ulVKCxFkF7wLMTsc0CxgDR+FTzEkx
k35L93z02eEggZHGTAsa342L9Fp0p1MZrWPqiDZTC0lfNcLSJMHOCnZcP1sUkvZ8
Kvayz1S/5L/4fBo1XXB7ZGM7KKfRfpmfRXWMN3azyV14dHsyhShXx3ILYO+SSoTs
PRarpddr8VDgMS/Suk7vwV5YTqCLWKi3x0MmqTJyr5yy5GZ5B3+cXy5YkX8J4VAE
o39nvCPtsMjGLn/XJ0xi7lCLDxyYnm1fKkNQcQ2Z02VKmljc2AFc1li7bolzm5yC
ZSOQX7u5DVA4F720CqiXmHt7GZgt1GanUgaS5V/46FLJcroEBvIqiNOaEDmtys8v
2qrXVPZkN1HkByzpqqWTuRmGkzcCFSCDIHOx/nK6BiRpR78mvd4I32fKoNO/7G8M
Ls8pgygWr5NDZLNS7hXvXL4AsSozCsU6fNCuySbOspfxm2LKQBRVNk3wD5xZX0px
zrcsQSCiTzFh+x0A/gonMdqSUVZFcm4Ki0bRagVBCk8QVSQExpUJNJQzfYblWLKx
CVH+F0dyJJ+2sRzYOSEvKxW2pGMLtgGKiCLBbiUnxSX+NeVC5dW3Itx4Sco2a4bT
vnIvkARRZftKBWYoPr0+2OS56fBeKJOBDOYvbn4j4WlJ/45CnJZnjIpgG+9YS3Mu
iBhmJ2blHNhgHJIa4AvVSzmFuFFWXyhs0rD5JouuUDYUNASehja8rgWLmJUhnWZO
uwXTlOhI0RtF2wt51/WtUzsILfE5124J2MAIQ8PL/la+t1YYc3TjNW1vuV7vksr1
coDBi50ni1utwWBJ4DEC88obqFYPmwpvCp5n7ak3W66U8n3ovv4gN5jU5bfrEkT0
TeApYlfnIBsue/8aFkpX1JbeXF90ktLMQ/emK49oGaOUaptVDP0w2riyBC0/F8vt
rjslf8gmLAHMmJZY+iOzxZsXsygQWinKGJQSokngGiK48r2I+Bct+4nRfvh4dCzq
BcrTBgWwT+q6J4wAsnWF2KsdZyo8o22j6lf00egABw/yMmrS/LWRxmm9bb/QNxnW
O9m9Br1l5c5iBy4UvqTGZkdREfbo+sEFgyeGJKi6bj5f1C8FQv5W5+81jJ6Tx5Gf
mPbxka3lGBFdZ0Qqv7sa7tCLGQLCtDjhXJrhUdS8r213I6R3tVNWnkXFQOSqWUL5
0Fiys6YaAwKajODwdfodGBVnxQPBZGD13r86I4dexhAlHErJPxQ1ToCaDPrvFb0P
LfY3Lu+X3uIgIuke+lJLrk289xVU7NO5Pbyzm64ch4bRJj/d/AK1ZrT2EK2DOuKT
BPeBknlLGC1CRBAAAMEaOKIWtMdrp0UzkpERAPfTFjrXsirKzywoEsHhfnLKoOVu
yzSS8A8kY8rDXVUGwOrrI2zaemgCCnHB4cTtJ9e44Rg7Gq20VR0cw5WNargEsZnM
e0LmVEetNFuPd4BKwW8yjjdqQoEEueAYss7UlgrKn6hWXrru8Y3+elXqaVL3EstG
JSzCkhY23nJMj/IuUw8w0stsPMts5eXNVqY+jbWDeHuDt/37wjrLbfd3B17Lbn/r
MRiWyEvvIvVJacVGP+A8AFdgTpKKZaXW9p5RNRCBm59Dk7hZdPeDx0jCS94+e1Y1
7ArzebgUQ4nthLaNQeNFQzJTSbaaOoVr1qgiC1w5y3X/+GAgUrTI8B4n81kYKq58
xMXSuGEBsjbWE5sxgc5jGTa5PWKKRxz8juN9vsFVUkBIbBdcrsx6uM7JILZTTsF6
tfW8KK310k6IgKmO6i/FJRgTe/xtUmXAEFhunNqaiMtKEt5eck6sJrriejm4cjTG
LiY3fAhkHsjB3x/jMqZGJO4VCystc1ubjQBP50dGW2Uvl+vZnYULkk/qwMu/dI9l
uPoId2B/gZ1XY8HAyGnM5uM0XagdFm+aVH7jSJbIpZJy8Bba1cCZHLdc9j5HjzCO
gaRcZmOkRku6i2XrkJckG5oR5oX0YBjUdH8EWS39iokhedQdg3qFmgkclaEHGBPF
QbbAZsExsV7Yp+k9onTQTuenC+ahPOxkNNoXldjqC50GsyXlqYHrkdd7KVtru/JS
66ARUxm2R6Bjhc18RN450XxMo+4qu58iP1SnvTjndB5C7bbKPcF/F0DpmD/NajmC
El5hc9zSsX2UzePkv4qJ0LWqfPT0uECFc2wgYaoKPMcNgEMQu+DldaAfItCrkoIp
+5RO2c9SbnQFiyHp0zxqPy/YMRuBGvJ2cqUoHMMQDZBHx+lpC9sysBdWw25UOKur
oh2KbRakofZq+4XnZgy4Cqd5H5k6jY11/3L6girSDzt/Y4UPCdx+J1RkgG4Y2Xyd
pPz1v7Q0PGAbu+t5x1k7zZnI/oUGs2TIvuNVF8tuwFZOJLp/N5xzzOdlFMsxbInl
uZAGcIas2UJYzTQ/bjnkfrhXoaXBoeZRZ7b52r+szPN3hI/TJUeGTY1RulvivV1p
AQzrtbmwSRnSNCJ0JYzk1pdXrDOJ/qCUqU+mJOBkDJ2T+dh8bDm8lDnTUBdlnVkI
kvU6h34bBtDA68ACO2hCwn8O6X3RgRiajQkd0pA4SPyehyeG9phakhuJCRIViBUA
7nZVkYaywWlvIPJkcZdf49MOwnKHcmLvpaMxMv4CvZ5YopBaPbFQIm6grIxJMSeA
pYUDXrciSFgGlV02xTRGiNrTzMEKSJSC/BDGpPIGJE8Z8BS3zLGdopGRb7LRxv5y
/CzzB9xxb3Q87sD239UZJrDC2uLMun+FIBGIw7xPs5Qv28AsC47FE4u28T3VkRel
c4cYmBvcrI4x+ozlcg3MHIpcdkKYYzKvPnMomiN9FzG2lv95PXIJC8kYnkGrZnU8
nxsVSHUbFalHIRd4AAp3Q2gDQeRefnDnxdAhOiwYkX2bXcxeGHBzEC+hzG7aP/6K
h1gLQNNs0bCQGXgO/PgkGvWe687RtQGff6Stsm3UzAzEj4eOm6uvhrtiJzAzfM5a
CJ4vsiFqNB1OE7sQxkIB6rzSpXGIYkk7UBMAdokncHXWaRy2FYSkgwjxOWNp08K7
2Is1Yn7k5IN34qf+rWUf2Xb5NlWxzK2fD4AqZ1LDn2TNgJ96qj6Dl2OGs5XwHFij
vS+I6bYUikmSWTDqUeDy2u/wiWyaGrdyU7QIxA5pcqNf1wiYbgqLNeCdQ/w94xAH
RdfSBlPEQquss2gPfcQ+5YCqbcoejkh9agXTF64JZapMti/rME/zAWiJAIxi0nQx
l9SHSwobSen9Gg+dLP0VC6AtZRzqpNaQ7OaXPcIOuqEE9c6xGxsSpTLL2nE07mEG
Kl4KIjqEThx/FjyMbLDsGAp7e++hrE2vS5joz3R4axOTrrBvYh876SPBL0atgPYQ
PsKFH5mgcgF+byLjNFyygHPQd3LGPO59TLjs2kUPJcTjSDQpt8BrzdoKiejNTJ3d
uXQ3C3whs+TCRIIyb+vcF4QF4b+pntLjoFBlwOfHb2IeLSPJLDTyedxFP/XFIDvU
i0EeFNFVZM/KmBqj66+BnxDDMkuu2vcV4MR3sFLbfhLCPw/PwFWvlm6UZ2bfAggC
plsuzgKFdwGxRYnJRh7G57gqvcyizHfuKd6QwRd5coECp8cGdP/Qh8IApZ9XJUln
4NYJg/adMy9bkiSFAoJ8yJIuV2MR7wPQURkP23cDW9qMvODuX4gnuUf2nyA4l0GE
GraraMZgU85tYTicwoSVsT/9kUMzrlkWBgR7BrUIXsmj6qUj3bQGBMW1Cuj5NX7t
7BsNKvzz1xxQR9sAr82yHkeio+M1+Uw4KCnAvKEX7l9tzRse2N2MTFgJ3wftA+8G
6iOMzheOkXIeS+2Mtm0R0SQzKD0m5lfZT2ZU9cfuj0rYWSXSCzpFsA8+kq/+NE5Y
Lm6PuXAhodaqmeW64kP8fn7eT3xe/am9oMSTmlssBd32Pz4JcxA4zyOFDThEmz69
GUr90A6hHl57j0TmJhN1E+anl2z5JnQ6x26EUtVc5ejbZH+oTiSa1oUdpd8yK2X5
gVLmWlcclmKCK6pa/dojjiUttTOV5z6K9OzvdiNolsPyWqc0rVnJogZfVOrZiZ+9
c8hob57oCR/4lP/79Ha27bhiSIuIj38IIpPXZCVOSuAhQcCoauRabRsByEsvHawZ
N1GH4AEvEjfBImc6KkNSLJyb+hE9hJEe3ShO+/ljSyUNWCrnfZtCHSqXa2XRheYl
UxpxvAq1+Cng650HsChlLNs3gEQMVN1MzudxevEuLNYiY8j9AMDaPykpHhcYpDW9
NjKJY9Y74h7eGQxT4gi+LjDp3jXgzv/oVCgO0+JRKHhdXO1gH2SfwO5SWlZsw7DI
D1BW7Z2MtfHhhfHdtxeZb7n7Mb/GMFV6ey0OU5qHHE4a+nzK5JUPOaqcjCEbdZBm
WNIDgGezb3VK0JJkkkSMFZbfk1hZMurxRnDEjIP02g27NGK2QiGNx48atQeZnahd
2Y08+99LtoXsHYK/cXQ0UFqnIyUpXHRhTNBgINdKHzMK8Ve/iR6BRBvsVLdqQjOL
niStNGcH9uOJuRMIVSLN74eGF7rzCGSSl8cBgOkcpLhRF1NnsP5H7ajfaEEkPgSh
iReHUbd2wlcbiRWmdOdpSNBvWuKYC7M94NX382YMD/HKE8lD1Hxy0pccj77JRIhv
kocxUMI/Fj3IJ0QfultxiYMvAk5oFwpnYkC0W8ws7wrnxh+k9oc+vknrSm5wLHQn
8fZobrFstSlaIV6/Q2cdSh0fD9RLzpSON86uMzPklnOXp6gS0HwkRkcA9VSWkG2c
Vj+I54nPdbP8WFrAsaoTy2G6TH4FJJ6jNcORJ8TEVudCY/8l75uy5yfbZhXCpzAf
XXbjNeHK1w44Jeb2L68EjyfEkbZPD7qHElDfUdIQ8l6/Yd+h9F81A+pAZh4N17a1
R/Sah9LhhIE9zmHznWibOK6cgIWuP8t8jtA50AEeEawtdrOw6rAy55DRYbRAzitN
UCJTaVPExzkjyIzdTnDyHOOhDhdMmV3avn0qTnkZhZSNagup7roNI4oMukT+SFU8
1A9ClM24DwbaX5i2YvT5YEaXGl620K6rmi1MfgvNBWxo3lM/IvE92UCdos4VvLdf
FYVgwbvtavWpjmDFIdmJOaRC1pkZvYWKgiEmnCFGjp1Kh4Gqc9doLl+K0zlQhtFV
N18G3LzWUB5DA9RFXvgK/Ibm16oFu1x0adI9y0CBIDISr3z04JTAa4vp3Q+rksX1
nYsFHIBIuUvEuQU9bMT1mu1B+j5VLAm0XJgCZ3esh5jj7ZQczehofLAjM9WohGNW
c0tSukMPVvnb1FIpw+Sn+CFdc0m5TbOM0Hrtg5jRyxL9fGRUJey9GMBlJWOuQwWq
pebr6Ywd+M74GWFWKwQvMTyzarD9xVGPtOZaIh4HoeAyNbXeuLdOvvLYluL4jVqg
wMhj1BINx55tR2kDRdzQFAzA59UWIZSlYsdOrKN3GCU1JcTQlNYkEOpeo8ZI1B9f
8iAgi6oJUgvaUeq0x0h4EIpH+rFUc916k5UUIGCBq+nar776OxHYKtyk0d5OM2o7
bhbNQMc4tr1WdAs8HLgV8CC5tN5JrsfXHi6nAo5XiWpYylOY6dfgIYbrp5V7c85E
Gkx6NU0CWjdAPjdDQ8zLkEmqznkc8i/lT/FdGyTrEHJ3xXYwaqWKBpGeyBXi1cSw
5qF2256pKRgMdpQecqH1lrasY5Whu+s5cOzW+JJI7BdUlzUsQ8JDGeZWraw8/Y1+
W+oOUqbyofzlAnNz1IuUdc2Jap40fkdnVbAOgvCmHQdFAO4KoXlEroJSERLh7PFp
5zawnT4sJtXkwdQ8cHE3iEWz9vHrdCTuUSgoG19hoB3VGrNYbu0yl0xx6R2rtL7A
VTay5bV40nHw5HwWGX2wbQyeAxR3U5szv8bmKcAB539Ha1r3XQhOoIutFG3Fzt3z
5ff/t1NIjeKmLKxTTofty7qsXkUnL9GH23FEnZBuXQf4DRTkayRF6msLXiTSUDCa
Viq+z1x4CgPknahWYKyrBd53ABuBhE+rUF1LoIGNVkul5ZX4cr1Mc1AFXN16ObeF
leAdU6fW+tN0lWtR9ri4lJ5fn3aKzrMMs56JKbsALUYuYMWY4MDG0l9hbIxvQ9BW
HBIuT8BjVgMCjCOjzGoDu0ZYIwhvk9CzuOpgekpO22CiVIjSwdnQPoeBVOM0ZALq
teYuqQ3+3E58UJYTPZ7GZvuPcyXTBaHuULneoM2Mdr9ikrHZdyqU2OxOSIiJS5tJ
55VmNB/Ry9LuIkgqAQkDI/Vu7KZ7etGNddMuIvT65G5D3hZp+aknozjlBF7J7QvX
uLumipo5b7PKcJ6kpNR3SAAC8lWQkrag9qFagqHTa1vzh0BP3+1BIzmWhJQkNRqq
41Y0lE/lec0+0WgIPUhTfi2cP3RUhhV+whdFwmkaVKGqBEFBBRoamqM8IT4EoSKf
Vcvdf7ft5KQMPKFgGnXoMcrky4jrDIquZjWylsaMylnzjTaSA6vo+EWguKWGTUgi
P4h44wRw/stTiY1dvVKKUvHIcI1Zyw9U6eImjOFZBEMk/VTpAXwuQF3gBtBbSRge
06zW84pyVS0SkUPeUOCfAdnEehNDQJbj016BckT45sNYA+5KBf9rh5ZxxdwCEYAM
aslQ//OS5v4DRhTjKKHgLaJ7gcZsEXncVvyholPmNGzCBMKGbORQ0dHt71zAVzCx
7P5GSocYWhhnPywZh1Tnc6jlGYQHTO84b2kGAzxAE2daUBV3NsKWsun+Y47i5fK7
Xu/9JyJxBDeu/o0do3KtznEvBXd+80xYTIgqUlT7SKuJ0HA+cMotxb+gpPG3LTj6
9WfDAiVGfuDS/NhN2oIlYiFztkQueMnT21NWohGB1GTdvpC2zVhUK5oUK6oi9Qzm
WYx3/iZ9liibNdYKrpKq04oUmOKZP1cEA4iXBMdlKY+VTXgw5vijcCozngWOPBCV
UF9G8XMGBhThVjt0bVWd6bxEjJo4D1RGVf8nfc4kxy0S4Va+Mp/7pNpln0yaj8L2
n3C9k8gAYYD2EI5By4VSQGL9uqEhqA6jQrS0s0hBl7c+mVaveSMUy9OeOshFzw3s
H/kC4waumnlQgqdjxgNVDs/qhq0ki6s4Rcpo1cHlPdxmtwP7dOIuJyIF4hbEPMGq
VXRW7Zdrtuj+2xWrjUvXONWIq/+gLZnBz1YABo307anDXrAJ0pMtA/LVcpX95V3+
AvN2Md1LraebVVwLVxjBp5pgheV0U2R3chz8qGoZPSkP2VjEW+j5UYonRjYcfI/Z
1hfy+fOqzA3Se/OiEAFLJA3G96O/Lt6B/7uVju3E+lI2sMEX6CuqvFHEhYgnR84g
LsYV0YUaieD1J2KMe68LPER+EgPKcJK4bR2KMwzvkBuBzWEXlaFc21PRBa/Y7Hpw
q4Nn0Ffx5ON7RwNUr8M5Tt4bgnI89LpDwdTfrSKNqyCVgnaI5gP4/0ZIL5hVls7H
cKoH3d78EkiUezbD8eYAzT0Oddf6b4Bz+BrBaQ5RHi5uqTWiPsQLRaG5ShN7jUdK
TM+TdrRBepTanXspju8vDHP+M0nNLOaobJe2DJj5/1fdhClHm2En3dTM00XPDGC4
fxRUH1aVlHLa4FGcu/ZnvYDWLC7dJA7Tc2HlvwN89NSk4vJuT7Mv7k9Rv/bNCDBm
ty67U90guTaFiJ+1IaPTr0T5IVC8HEFPS87qrgH+VeY9LvTane6w/CwWE4XXzTR6
YDzGBn8KvJIcu3MGdJfcoZfXUr2qP2Dt0m7wT/YtzgoM2v0BLLzJdwid+8ehv95z
2UJoBCrVIL5xO8/St010I3LB48CJqHX6t99hsm6mMrTW140ZCD+tqQf+pQAL8kI7
4jkoVNW2QfYsoJl8ye7AWcit8CEXKrFDrgAtD4fxa9Lm9/vUhqOzyx078W3RHFun
Ezx+lvasVsIUYZAmQfPzAHzqHr89lxVn9otv/DPKsto77eEbQ2MXHxFcsIomQbEb
PnxFM+9Qlffp+PPfm0cZ+9OV18dasizuts25LQ75dG8t0IHbNkJY2YlXsLr6zoVe
WVE5CM4cyI2MKavp98MOf14frdF+ViMHNA1T2Ei70pML57kT4bHmT99JAe0lT3GH
zEUSl4FcUa+sd9Dz9rpZriBUU5yA4pCyz3czF83rEKftSgQurJS2E828xhoeDoJ0
LAaRn7Fz9eUCFnAdaBxFzbUpX1IMg4sOLIQnC219h7iEpCVz3rWqBmiQoCsMY8Ww
nfY6Imo3GSJ3uujIKZn8EkCQLSHwDTNKJy9W29Ov5TZE5UQMUHJxFL2jgTADuC0L
6dcjj1nHKdG1Z9f8n7OGqS8mGYvmvLHIlOc8OF3N4F0JAUCMUKh53SU3y/LcDDxy
EY/ZxVo3RA+beKjbXyhfLHKdLGGqxnQNxaUGpahqaQ5fDMEcx7HJOJSKvakcEaM0
hEDoEGJC5C2kYromUb+YLAzm+a2ksPAc0hANnI8ruYOm2b38kuNUrbZTxjRPTW3N
6eu+iO3bHg/yOOHLPX0xNKUCqRr0qeyPITyC5sIu4raQzmzPuMXH6UOTT2UZ4VfO
/HDtOFwL9gJZnbXo+3469Q+8gR4H1wnjvAj6yTrw+gyjAE3V7WOqe6NEUOqusLpm
+t1NU5RSxuelui1t3y3adWVvwB+axqthj8eXxft7adXZTIeUyrGodG2cGT89VABm
UULSY5fBsxZnLiRh+fRh6J+BCJNm5XtAFmoPZSP7qx82xlCAqBpQpkAl6z7Th31p
EddHlU1rc20vJ/syTutdZ5nQ0EpblT6BZcHHSqfFjKR21OT+2770Sv/E1H+xNmfv
yopeh4gy/qpH6DQht9JqwvxdQObX3tb/bNZLJLJbsAho7YW8zWSZCc7XND62i/fY
/Jd0Mhp9LtCL6ADmRcw9kjC78mBRBRuSzcSn6uKGCR4vod0fkdCxD/tIEtbywKzL
Dp2cBPgz6RFD5TjMAqeK3y39rdhXmSQMmR7WTOoydvGGlIy0fiWOlegOkjaXro+k
XxBLxq6H7GiguxQcfPZERcq7mycDz9XMXSnc9MO468PSx8kR6FBFyQoiLKAmoHuL
vFgX6bq8gwLqz6xFctoQ7H+xuqE6PdSffIhqZ4vFpUPsfJchid6Lb9wSt1W5RBlD
akQKamubIS+g6hxHJBbwYDH18j0c4R8aAvJEbVAUvAyqyTzVJoETpjQsOlQw9T8u
DnagThnp7tsQcW615VYfz6PEzteyKGjSVPL2FXgBBYv83ztXIKjbxCYO9OyGzl8B
ilBU7pt28q7FZmxslzGgTpRmCVTy30+p5q3fAt4r5aPfPLHZtSXDaokXrhDFjGEw
u5hyn66tNgQJ0kcnO9hcICDNBmP2NViNlqGMkszy0Ib1RPh6LnNYU3N/NZxgWI6W
/4tM3c5mlnzhMUOUvrcj30mrodBi23VY+0hYYQerdux9gWYsn6Tx1+7mUacYVhEZ
yI+bOXkmf5I28dUqNH0s15eUHhnkXRzpADyKSlPXGR6oIL42c79s1ne3VlMFqq9S
SYzH8j4BQv2mPhgFCnSjF+BDXAMxVzA6+xvhEtfi5r41V+q7wWBCIc+swJlLax35
klplzaubQnDEBm8ndN7ko+KNsJnYjQx8nr7NSz+dg9Ldp4rMtTuZgW1XG29wLnOS
MXHFnr0NU/OAFmtCpKoMjH8wzYjX552ywntV1wI5IM9Z9RGR115OntEQhhA07MqS
o+db0d+eGVEOjAy66AD8J7cI0fi9nbo1MC82Msk+oxtUmSu4C93zKiB4uxvLVh7T
Y5a+WqaoaUrRkRYSK8dL1Yb9rdq0BuxgZHQeexX7lwddnjoEAV5+YxPT4UPUt+zq
Iu4VuGRXAitWawiYs9UQGLzBQOOgRDW1CG5JN3XKHaum6Ng1dLrH7lifeJeZeP4E
x6HoUMC+9AHZLQQsqaPWW/fiXaeIQY72ghR5aU1LUvcXW1opU6NXRNu9LFiLU6IY
6dueHbSxLVOvj4HClSsiv8VkBAJXykS9FbfJbhofSpynCOBMxKbkdgWByBB8wM6c
lBUM+oYAivqSi54KAwQfVIwml2IsxKaTYt5GuTJNDidjvsRibMdB2Hd+IEOf9/wd
ufeG9G/96Ou8Nuclfr7D+Yj6acIROZSIzDe/vALy0Uc1TQ37P0WGGlih+cBltMqz
6KXyU1zgOEIBoMu94DL/TF3J9AU7s76NO+/mKj+8weh5mqI3J6wdNCxT0UoTtovp
WiNQ8tHq6adCjJDT7VWQeLqDiUlHMFcvCgcEPtvJv6A7+Us36wcWUWCPCae1CVNk
qzSKHgsZyzD5q8pX3WqjI7HZEAzF1BHv4mJMDDfslSWwAAIu/lgH3HDsNnwHN5xo
WSRHXh7abwqSqxKRedv7iJ8SRxx/7IW91pQr5nufdDueU75akR6vCym6vmtDBSr9
N99OTJEpJYdecTJvIN4UGTgPLfSq9chL/JMguYYq41utdhz3xi25gQ96LWadIN/2
DsH3pOtiPROzwkSVdH6aJ/B0Ot2lXjBH+8QoqmfvfwZL/YGwtMP5c+GDlT5b4X0V
/aYWSNZDcd0EwF6cBbGYE7uS1Tp2o0Akz8kO1l+o0urHDIfNfHTQfo6U0iyijLwO
5AYF94YsaoFL7dABUOVgIeXR+UFEJnTxUEcV+lg+1GjGxYkMMnJLlOleFxcUBCJs
fdqVijR8q69PtviyKICLZZcJZ2SmWXf6rZI6VR625STCgDaJRncCLpaNOsRxo8Rz
xej0tecilUxzDyk6ReP74YVrYDJiSudBD8BPKAakBqngIDCReG0kaBeR+X2zH1tY
9BCeJYXCmZsWLqyWPnttR8zuozkpmpQeCZ03UpTCaPHfwrV9cIXPmttO9N3+Mb4j
vbSitbzgBRiWjfwX76J14bVG2Phb/GZ0KgBgZaecv0FBidtCJi74EcJCe9j2b8hX
VXSb5ZQOnijvUDdTalJj4D4IRHdXKidMcYF1WyiJ700Pg6X9/cCb8RBK8AaWv/JW
ktJJT4kWx3SKc/OWBoAjj6JD1WOj/EdAgZlUG33j7Us6Z5KNu+rjjDjZmckOjCua
Dxgx0RkSCUDYkwiGG7lGO5/PzRjE94qW9xK+iN8dp6Otszq2wrIHgMMRvcLKazLk
AONhP8ZicDQn8eiYg+U8TVDyHO9GHA6W01rcjNc3CwhyJGfc2UtJ9vzH80POwWSm
lQuoQdFEybTmGaUe4j2wiaMvqc+HQJ+Joba1alVsEjuHGDPWIuYjbMUUT5+xVRvU
JyfiPP/hJuq/ptpguzPMfh2U7fm25JqP0Ho2xVJzwW8goamWLkDhZdDHUptZsjvZ
CQdIzwp2IFhBmjLtP3Dky4ptPncHzffIeK+nQsNQVEjKBdXFHJRgbCzjO/4zErMV
of3TsA9aVBIAdZfNlB9ZRetm97L4w+ip/gUxbQl3NAYs6O4xbnbb5RAo0vON+aKM
2iEpO/5N3MqjbidvZizNghY/BBs/lCuMSmxNbf7D+Gug+j+NhcIJ3gtC+fL09u6N
ucdcvJCD1vEWuiCqdQFCZ9rhEHNiTNQNVRS7F2dg1VGkzUgrvFdxygwVs2Z1A90f
X9DS7fpTbxQudnAudQAfDjlhHrHkaEsbWJyx/1OVfd2xp3hW8CNMd0IAdnphqDBc
WejtGms3HXzBlohIlUFhxhK0A8+ImxKdJ0VuhiYWyQdVP+JfNFGtbVmrvLYdhOWk
ttESjvCI7QNee3gUW0s5WkqC2OWNEc7+QHqoRX/XKcmDaZE7k6zq7eSWLiQPGiSH
VC5WqxcbHxeJGJ2QddDK03bdWNEgrAL8r+w6vZY0B0qo+iJsvyARf10IjqbARmI2
xzromYjjs/mA4CEokDdswc7eL8p/aTHq//p3WiNXSx3mL6ChZbYU/RVXvACdyaFw
2swpxzSYcmELBNYdBasfGMsYv+Ekaap1Buw3qipXisZhxcVfua04c0HidIkXNYqh
4SC4rFH87R+g4ktF93h9Ikxx5Op3zgbQT57dZdeSxZ3Qf4COncP7yGJuUq0joSRz
sZfhmLbjmp0lEw4vPr0txQJXvkyVLx6avnqqD3ut27/mk+iGTgL32xLxpYMjj0zX
aXYH2UdSKcXMq+TsUGdp4G3HCfaTN8xi/SR0GX5ozKsqRFpnleXOQR5wJiiaazDi
GCxlp1nJR5RTdTD6HrbIitnY1Il9w5W/GWvHMRML28vQTSJgfZcyTdCy9EBJsr+Q
mfZNe/PluoTQtEdlSm+8RoEbzstoG3Qi09mOxMo97WFoF9f+OvC+a8yxA9RK9Ool
AdW0xha3trxHG4OUWjgxl96+Ea0vh85h2Q+1oX+CL7nFtYCtB0XNeN2qYwv3iJxW
kBMk0DW1c5GgEIylA8ulZjbKckKvelijqHy6mOUAo3Xakps6iMpvw84HT3en+Zc1
QpQCxcHVTWksc/iB7cSwmqt1/GXw3Bui9mENO6SRh/n6I5ILOC7uOtea4MDfxuf8
4ffSYyt2laU/zoNOIm3B5lbNH5bgXcMxaq1Vg2qqIJ7Uxfxukps1ZdlCHoISdDMV
hPT4OYST39T32RwtLm9SD/iRV05zbZwKemNGHnUaKCU9dEH2OCGZpB07WrdcYGef
6JpSNO6etSf6UIn7UssROLFkw1n6nf9LtBmww0ka8HHszdSM9wjC8KAF7tZHFN6T
hJdo6DT/XnFKqOracyzpmpEtWIgFHLqYmkV/kE5mXOEmW2LvjtAR4TOpiERPfJhl
P2JVj4ZfPdDoOnm1wJ8Br9HOrsc7EfFIw9SAMaviYCJnpZ5YdceLUy8UJHK9rVqN
qgJ97duj0P4IY+cC7dfRqvUujHF8jU0hEZhSB86MRViPZ7lSJR5GwpWzWVW1EYak
3qd0zM+kCeqy38SGGwb8peuzevXPB1TKwvded7DUx4XXl2XzMpo1GXuBOTL0kDAC
/7WYLk5HOSHDsRiteLJM94453htFO2mSZCqBm1d+1A/OLh5xlh7w3COvHb/TXUAG
up44Nd6Gl9/kEa5BwCSJNYDPXhL7hFzEyOGZJCLjkYiszeVrlmhfdAWpeOtbVTCt
bI2KlOctuODJTKfhIqFDw+qXcQ86T5wxJhvQqLCbggUUvckwO2w4UMbdiNSTzPfa
3Rj+NV5jQxVtO49Id2bck/sV46BYNffmPtc88+kGRpqqC6R9vSpDbjmMihLBpsM+
lZKA8sGjJW9f1ILYuyzN75bSLZP+c9MMFyN/HpsocKXDzols53yWfpifzCR7Z7tO
o2QiPHh3WgAwR29nWoV9qw==
`pragma protect end_protected
