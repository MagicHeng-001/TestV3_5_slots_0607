module altera_ldpc_wimedia_enc_ROMs(
    clk, 
    rst, 
    in_addr, 
    out_data_ROM 
);

parameter   NB_ADDR        = 3;

localparam  Z              = 30;
localparam  ADDR_WIDTH     =  5;
localparam  OUTDATA_WIDTH  = 8;

input                                      clk;
input                                      rst;
input   [NB_ADDR-1:0][ADDR_WIDTH-1:0]  in_addr;
output  [OUTDATA_WIDTH-1:0][Z-1:0]     out_data_ROM;

        altsyncram #(.operation_mode("ROM"), 
            .numwords_a(32),
            .width_a(Z),
            .widthad_a(5),
            .outdata_reg_a("CLOCK0"),
            .outdata_aclr_a("CLEAR0"),   
            .clock_enable_input_a("NORMAL"),  
            .power_up_uninitialized ("FALSE"), 
            .ram_block_type("M20K"),
            .init_file("altera_ldpc_wimedia_enc_rom_0_data.hex"),
            .init_file_layout("PORT_A")
            ) ROM_PARITY_0( 
            .clock0(clk),
            .aclr0(),
            .address_a(in_addr[(0)%NB_ADDR][5-1:0]),
            .q_a(out_data_ROM[0]),
            .address_b(),
            .clock1(),
            .clocken1(),
            .data_a(),
            .q_b(), 
            .wren_a(),
            .eccstatus(),
            .aclr1(),
            .addressstall_a(),
            .addressstall_b(),
            .byteena_a(),
            .byteena_b(),
            .clocken0(),
            .clocken2(),
            .clocken3(),
            .data_b(),
            .rden_a(),
            .rden_b(),
            .wren_b()
        );
        altsyncram #(.operation_mode("ROM"), 
            .numwords_a(32),
            .width_a(Z),
            .widthad_a(5),
            .outdata_reg_a("CLOCK0"),
            .outdata_aclr_a("CLEAR0"),   
            .clock_enable_input_a("NORMAL"),  
            .power_up_uninitialized ("FALSE"), 
            .ram_block_type("M20K"),
            .init_file("altera_ldpc_wimedia_enc_rom_1_data.hex"),
            .init_file_layout("PORT_A")
            ) ROM_PARITY_1( 
            .clock0(clk),
            .aclr0(),
            .address_a(in_addr[(1)%NB_ADDR][5-1:0]),
            .q_a(out_data_ROM[1]),
            .address_b(),
            .clock1(),
            .clocken1(),
            .data_a(),
            .q_b(), 
            .wren_a(),
            .eccstatus(),
            .aclr1(),
            .addressstall_a(),
            .addressstall_b(),
            .byteena_a(),
            .byteena_b(),
            .clocken0(),
            .clocken2(),
            .clocken3(),
            .data_b(),
            .rden_a(),
            .rden_b(),
            .wren_b()
        );
        altsyncram #(.operation_mode("ROM"), 
            .numwords_a(32),
            .width_a(Z),
            .widthad_a(5),
            .outdata_reg_a("CLOCK0"),
            .outdata_aclr_a("CLEAR0"),   
            .clock_enable_input_a("NORMAL"),  
            .power_up_uninitialized ("FALSE"), 
            .ram_block_type("M20K"),
            .init_file("altera_ldpc_wimedia_enc_rom_2_data.hex"),
            .init_file_layout("PORT_A")
            ) ROM_PARITY_2( 
            .clock0(clk),
            .aclr0(),
            .address_a(in_addr[(2)%NB_ADDR][5-1:0]),
            .q_a(out_data_ROM[2]),
            .address_b(),
            .clock1(),
            .clocken1(),
            .data_a(),
            .q_b(), 
            .wren_a(),
            .eccstatus(),
            .aclr1(),
            .addressstall_a(),
            .addressstall_b(),
            .byteena_a(),
            .byteena_b(),
            .clocken0(),
            .clocken2(),
            .clocken3(),
            .data_b(),
            .rden_a(),
            .rden_b(),
            .wren_b()
        );
        altsyncram #(.operation_mode("ROM"), 
            .numwords_a(32),
            .width_a(Z),
            .widthad_a(5),
            .outdata_reg_a("CLOCK0"),
            .outdata_aclr_a("CLEAR0"),   
            .clock_enable_input_a("NORMAL"),  
            .power_up_uninitialized ("FALSE"), 
            .ram_block_type("M20K"),
            .init_file("altera_ldpc_wimedia_enc_rom_3_data.hex"),
            .init_file_layout("PORT_A")
            ) ROM_PARITY_3( 
            .clock0(clk),
            .aclr0(),
            .address_a(in_addr[(3)%NB_ADDR][5-1:0]),
            .q_a(out_data_ROM[3]),
            .address_b(),
            .clock1(),
            .clocken1(),
            .data_a(),
            .q_b(), 
            .wren_a(),
            .eccstatus(),
            .aclr1(),
            .addressstall_a(),
            .addressstall_b(),
            .byteena_a(),
            .byteena_b(),
            .clocken0(),
            .clocken2(),
            .clocken3(),
            .data_b(),
            .rden_a(),
            .rden_b(),
            .wren_b()
        );
        altsyncram #(.operation_mode("ROM"), 
            .numwords_a(32),
            .width_a(Z),
            .widthad_a(5),
            .outdata_reg_a("CLOCK0"),
            .outdata_aclr_a("CLEAR0"),   
            .clock_enable_input_a("NORMAL"),  
            .power_up_uninitialized ("FALSE"), 
            .ram_block_type("M20K"),
            .init_file("altera_ldpc_wimedia_enc_rom_4_data.hex"),
            .init_file_layout("PORT_A")
            ) ROM_PARITY_4( 
            .clock0(clk),
            .aclr0(),
            .address_a(in_addr[(4)%NB_ADDR][5-1:0]),
            .q_a(out_data_ROM[4]),
            .address_b(),
            .clock1(),
            .clocken1(),
            .data_a(),
            .q_b(), 
            .wren_a(),
            .eccstatus(),
            .aclr1(),
            .addressstall_a(),
            .addressstall_b(),
            .byteena_a(),
            .byteena_b(),
            .clocken0(),
            .clocken2(),
            .clocken3(),
            .data_b(),
            .rden_a(),
            .rden_b(),
            .wren_b()
        );
        altsyncram #(.operation_mode("ROM"), 
            .numwords_a(32),
            .width_a(Z),
            .widthad_a(5),
            .outdata_reg_a("CLOCK0"),
            .outdata_aclr_a("CLEAR0"),   
            .clock_enable_input_a("NORMAL"),  
            .power_up_uninitialized ("FALSE"), 
            .ram_block_type("M20K"),
            .init_file("altera_ldpc_wimedia_enc_rom_5_data.hex"),
            .init_file_layout("PORT_A")
            ) ROM_PARITY_5( 
            .clock0(clk),
            .aclr0(),
            .address_a(in_addr[(5)%NB_ADDR][5-1:0]),
            .q_a(out_data_ROM[5]),
            .address_b(),
            .clock1(),
            .clocken1(),
            .data_a(),
            .q_b(), 
            .wren_a(),
            .eccstatus(),
            .aclr1(),
            .addressstall_a(),
            .addressstall_b(),
            .byteena_a(),
            .byteena_b(),
            .clocken0(),
            .clocken2(),
            .clocken3(),
            .data_b(),
            .rden_a(),
            .rden_b(),
            .wren_b()
        );
        altsyncram #(.operation_mode("ROM"), 
            .numwords_a(32),
            .width_a(Z),
            .widthad_a(5),
            .outdata_reg_a("CLOCK0"),
            .outdata_aclr_a("CLEAR0"),   
            .clock_enable_input_a("NORMAL"),  
            .power_up_uninitialized ("FALSE"), 
            .ram_block_type("M20K"),
            .init_file("altera_ldpc_wimedia_enc_rom_6_data.hex"),
            .init_file_layout("PORT_A")
            ) ROM_PARITY_6( 
            .clock0(clk),
            .aclr0(),
            .address_a(in_addr[(6)%NB_ADDR][5-1:0]),
            .q_a(out_data_ROM[6]),
            .address_b(),
            .clock1(),
            .clocken1(),
            .data_a(),
            .q_b(), 
            .wren_a(),
            .eccstatus(),
            .aclr1(),
            .addressstall_a(),
            .addressstall_b(),
            .byteena_a(),
            .byteena_b(),
            .clocken0(),
            .clocken2(),
            .clocken3(),
            .data_b(),
            .rden_a(),
            .rden_b(),
            .wren_b()
        );
        altsyncram #(.operation_mode("ROM"), 
            .numwords_a(32),
            .width_a(Z),
            .widthad_a(5),
            .outdata_reg_a("CLOCK0"),
            .outdata_aclr_a("CLEAR0"),   
            .clock_enable_input_a("NORMAL"),  
            .power_up_uninitialized ("FALSE"), 
            .ram_block_type("M20K"),
            .init_file("altera_ldpc_wimedia_enc_rom_7_data.hex"),
            .init_file_layout("PORT_A")
            ) ROM_PARITY_7( 
            .clock0(clk),
            .aclr0(),
            .address_a(in_addr[(7)%NB_ADDR][5-1:0]),
            .q_a(out_data_ROM[7]),
            .address_b(),
            .clock1(),
            .clocken1(),
            .data_a(),
            .q_b(), 
            .wren_a(),
            .eccstatus(),
            .aclr1(),
            .addressstall_a(),
            .addressstall_b(),
            .byteena_a(),
            .byteena_b(),
            .clocken0(),
            .clocken2(),
            .clocken3(),
            .data_b(),
            .rden_a(),
            .rden_b(),
            .wren_b()
        );
endmodule
