��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��CN�M��rY���k�d��%�����]1�d	a?���u�P�e�q{�;&nĲR�OL�D��M��:O!����߸���:�6���R���{=I�9`�DW��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�I��U��RT�k�ҡ�ˊ�\ׇ]`��:�VF�'ު�ƿ�-���%&`�����5)Q�q��:��Jd�mv���0&Vѝ�ķ���lGӖa���ynw�4��7OEQ�%�������5)�K��������k�U,c;S���ic<�U�a���Y��I�;��mM����hXhx��#��Z[��0�4ù0���h70��@�܈,Б�+���>c_����~��L*|(5e"$yRuD3o������y�k��q �)���˺&]��#�nsW�bU¹��?�r7;f��j!zh1�,�\���'�U�5�M��X���#he�����3p���vX�YH����������ô?��J�:+��-��j�c��^��v�T*��u�x�:�H�&/ہ#�>-+�0������ub�u��U9�'jf3GNH�2%c54_5�LC��L\�ӵ�ܬ�U�۷�JX�|�f�����5e���z���W)oj�j��'���z�q�7R;)5���=q5�(��1�E�T��J��z�|�C�h�w�$���TD#"�.���� C/�b��_��V�Rq��n$	��O�
!�Q<�ј�pVm1�Q�beq��YBs�:��;��X�+��W^��J�o���v�!E����
�� �_�y(rLL�}�B�󣓫$�F��PE�2 ֛�$s��~η��[�c�]"��e�md ����T����>�q����-�*1]]u�B|N��ګ���愋|�⒗ŝJ�́���Q����������$��Yķ���BR�� d���������B�W+�U��0k����m/ȍͬᎰ�^���&4��1L����>�ȎȺD�Ե�ڗ�1lG(SF'���b�c�Od:;��܈⯨�K����h����¾�$��76���怡: ��@���-C�s��ǥV���*��N�+�[�F՛��u$/��-�X	؇鹓�S���u�r�����Q���� �9c� x�E�BN���l���A-��M�.��n�����C/��A]Ɍ�ѣ�Y�JL�GÁ���I�
!o�e�� \#}��%rů���]D5��zk�����vt�s�@��,�n0\M
k��k�o�m��7�d& "�I#����r8�&I�$v%���y=R���2�.@���Y:L�n��8�3l�0W$��`�S��J�@�i��c}��,׉��e\sy�_h��3u|�Q�Ľ^���k����A�s����8�d�*��||��d"��[ev@��Z� ES�Lgצ��Ĺq�3�4�U�MB�T���Cu�T���?�e15{%D:D%�}+�3�!��.|a]����̘�N�ݰ�!c�����.(/'
���K��:�=���g8�zF0���x)@v�J�}��WV����;�$F��o؁g��4�%�܊�eu!?��`!ˢ-s��Nxn�5-ȧ��O����2j.p�L��UV��:�,�����?�(ކ�T͍�al@�R�~�*SE��B�Fκ`���w ����p�A;��	)��J_-�")�lQ��q��SI2'^�H�����,��J���O�~>/�,�\�
�y���
F��"��/g�Ti)��t-["Z��+[Ӿ��ڒ�|�	�^+1��ݚ���!��O}-�_��jS�BMt
������g&��|lsA��h>��J&y�x;������+�k���͋���e�j�o����&��;�W�-Ƣ��иXԞ�P�@x� �eջ�7���.���b�\�����,&$��T(>b�wXϣ���X�عb�����KX�O`�PFu�*���h5U��$�_3�$�M����������j��5�t1�$��ٟl��}���X�סIH�������3�G��̈́Hi��آ~_kK�$\������lCC#)�~{ׁ,��Q e�<�iq�VZ>\�h��G/J���a��S���'7����g�=�&�P<5OLaW��x���χ�`�mWȩ{��pts�{]jg؄�
�������{�	�Iu���#��_d�L�d�R.Wh]N�ո( ��K�e����X/�3xOxu��=~җ���?�q�P�I���@]��lL=-�f�D�[� �z��̀TR$��c`�c��)���'q��$��d��B�7e���P	�͡PD;�>�� bRX���T���:��=Ƅ���M`N�gX�&�����^uKδ�(��@��@�v5[3Gz�W���-s��}�J)���Ɉ���nn��5>��k��rN��m��+2^OÊF�LP�����E�Z7j�cn�\��'�6�x��;6鮍�)���ù݇#	�JXڠ�Ӟ5a��?*$<�jU5�!��{ �JDa^�K.��E�"AT6A�p"Wk��W����/��0o����3ܰ�C��\z�����NKY)5�k�G�Xn��,�h��4i
Ot�oP�xѴrMk�R9��YX�3Q�Î��3|: ���m���#�����x�����:����Y�g���	<����'r�ъ�����B��\K,����,m�w���>v�����T�J�Uj%؋�%kjH�~.��!J���R4"t�r���nH����ҥ[��ݼ��HB���&����x�f����x^4E��TA�7#��a�0&�y�4:I9i�W�>�w˪&�J']�'��B,�"�]̙K3�&R$�<؏v��5u�Ә��~$
~H��FK���!����`6����C�M�b��(w�^=�Җ�)���O���ZR�P4!��>3�����{	�Ps�(�E���h����w|�gSj�r>=l�\�ݯ,�h'��^JԹ�}�;������x�����5x�V誸��"g����E��N�{��asBVzjXc6��$�\�5���2��B�� �g�U���h篈~]@B[ ����Ux
*��^��>F�N��Ktr,����Di���۵d&W�-��k�l��UW�@Ge�`�k���ֺC<dv���R��I`1��Ϭi��ҵb���o���z�Ÿ^�aU��8N^�I'��Y�P�+�@�/2!���e�߯���	�B�����u�4��]������ރ����𴀛Ji���\F�-��͠�T.�w�	L��$$�/��4g���Ά������We7�3���VWH�Q@M/X���M��fr6>�u腐xT�EC\��Op��4�kh���n/(��������P	��E���H\`�S\�]�t<��cpw����mѱ2~$C�"��A��Ⱦg��^Ǖ�y�,�:�>)2��o���nK���U��t���+]TrY7��:_����:z�pk6��n�r��j�6���V��SX�Q	dB�N���z^@�--TY�j?%"\��+v2�Z��&%W?З%��t�.�!6�l�+�zr�]0�ݕ'��\�͓6��Cҹ�t�&�`�C��?�bT=��?���9ν����3��f��?����4;+5M�߮q��j,�j��U���3;�,��G����D.vC�%>i}{������#�K��\=	����.{�|u���&�B�	'w�f%�%OF{�i����ƥ`��z�b�W�K8N�=U��4�����G���^�Y �p�$�W��A��#D8n� ?����\�Ί�1��ó��Z���7� j��d���w����nx� {��۰dMf�[:j�ޝN΋���/tʏA��F�;	]X�&a@0&2)+�:49B	邕��f��~"��
<���|Y�+��f �`�%a��
�g���攻��(�I��n��FV�T�N��fLl���0q�.�|��r{����ʒ�,2vC�T�Y�Cߘ;P�/�Y� �n0�;}y�[+#�}:��5[ ��n�p~���V�HK�������A%� s�T��k$N�Z��x�-/��^m�t��|H� ���T�|UbB�\��R�}�hdn��/��l�u���%e��~�	��qřI�����'xH	��A�<��cR�Q8�y��`�(o�aF,�h?�)�̑�Ǘʆ�%��5X��̂�L��ZnQ�1��0t7�9e�.ͬ�$֫@�ߛF����1+�zb��Ґ���f�L�EdޏyU�E�4�x�����U����
��=)����u�E�2N�Y�~�xo��K�_x� ���8(,1s�<J��{b����~��z'�0���<mC�#�?��}#So �ʺ�"t� ���`N�� �0 ɵ�����x�\��9FJ?n��5]~�@���`�d����$9�������NL���f*]q��~� ������|*�kTI��!���F$z���h��j3s��#�Y7�M�;�σ �*����^���b����ڞl���O�Q����A��r���z'�$����Y-��!D���>�˅� �?@��V�oꔃ�	���b
�+��Θ��H���.����:غ1��F�,��)�m�����}u[?�X^���	]^yE��m[<�~t<��W�N]]#�n�����كA�~!�Rq�t�=�"��A~��67���U��Řf��N$���T���_g׀C��X��~�p�=p�b������f�k�2�8!T��̗Wi�.i}��ᖸt�c�xb��<yy#C�<�'@��9��8��0�Nr�E�1AS!2T��0������8/���!�)�<Y"�.Ù�W���s�L�ڨ�+}7��Q3�0����� �A�$-���׋��:�������&��pW��2��$p���Q�>uŹ�I\��^�y3Is����{	6���<��9�0�K���Qw2���$�D�1 R��u���ma���el=W��؏�
�R!3�wƳP�ޠ��}�K��m�&q�_�*���A�f����EFTX�Ug��mV��)Β��� ��5��?��K�ϲo=��<K��+��#��:�}��x�|I4a�uѪ=���d���6�<�K���Zj`���
�!�#�C#�A?�<A���A��ϯ��L�E�C�!e�n8)5���93]Z�aB�̖�I$4���$�<��$U�S|Ԏ��A�u83��[��0�7u��$����Y̅|V
9�)�D�~�Y��J�'�Ve����]�U��~����7�(�G۩)A�$+��2��Q����%�ڝg�$��VG�������t���C[�(@a� 7B�8g��0�����+���b�x+ĘRt��B}����v�t�0�J�O$�)��^d�� U�݊z����|��n��&������Ț\N��Hi}�Nj>"�?�z�b%�W�R�ҲF_��0Z�E�%�Q�|h�BG6����d�߃j�sP.�<�԰4���X�Y|�-���CP�����lY�&����*�[_���/t?�2��؄�vԻ�r���NUX�!�n��/��X�5`mn~��8#��j��%p*eZ��vx��2r�$]S4�h�)>��\'Ta�C问dYL!R�Gƒ�pF���+�5�U҇zF�iG)���>_'8G��fmw�$lw8��ݝF&�B��=����9[���ŹO��ځ�^;L`"���qw^��Ah�{��^���`�1�+�1#/f����/@O��=o�\*K���2�[���-��u�{f��.�W�G�x�uo��/z^_�rX��⑊q� 2�,۶d�lӧ�x�j3��E�����R�ӧ�t��b먅�j�z�x]�� B'W�:I/��U��Y���#z%=U�PR�.����T���xY��{�N������+�i"	0�%��*K�u�e��	�h j}���y7�a`1��1w9큿�<�X?�=��v���*�������:�^���$I�\e�'�d��p�u�m�7�g����k�;@�Ʊ,^-!/��J.ʐ�ؒ�u��E�3���hx 
��Y����$S��+~ ��X;���
ߥ��͋�Ly%������m�O�3nKy@t�\l]���u�t�:�����:��h�~�@zȜW������	we���kY�3'Ǌ����+G�)P)1���94$���gS��%RH�7m���*���|fTGFG/�����>�D�X*$��b.�{���x8�ZT�"/��C%���V��ҎH�砋�rFVg
K�jQ�&>Q
 �8�����Ռ�̭�H���F��PQP�U��k��S�I�N<�U�`����c��/���w[��E���ݲ�g�jmG�B	�:�;�SH?�ް�>b���r9��+���<J�4$1ȏ�	֥��Dr�U�ρ"V�_�pهӒ�L�	m�g\��D
Y_�c��v��E�JN�k[ [ �f���ӆ��: ��I�\�!6TA����?W;.�����P�)!Z�P:י���<�_�$�I���,��"Q�d�b�Z�1[�P�\$�O�x�M�ϾV�K��T;������+K�2<xˎ�W��P��%�����v�sŪ v�x��@n&�Bn�xm9캺Q���z�)=���ӌE��{��5�O������?�&���֩>�&��}�C��5��Z� #�l��U���������c�"(��pZ�p�R���B���f�_g
�6�B�GJB�=�*G萃=J۷��Ef�������xzW3&ЍlE�o��
��;��� �ū)��pL��S��>�^�i[���3�#,���w38{V+R���	��y�=-`Cѝ6Ѻ׆kP�l';�:]
{J���2�O�zI�"�O����Go0��7�tX���Y9��~@� �b�����Xlg/h�:��	2B�ғGv2�P�H����!J[��v�@�h5���4C�)'ya��=c�cYA�,L������83�VvϧOЛطˮ�[��{{P��p(Ғk��N����w2h�_!U��ı����+[�����Wj��f�6���.Y������� WnE�g%x�93d��}uڞ��������?P�e��>Y !w��J��&����_{���!h�Ũ��������Zm"�7o���ܟ� C��;����1A�r��IEm��0d��%ވ�x���}ۨ#��ݚ�IC��&��eY:|rTv�=�X�|���jE��<X����?נ��6S���s�g� ��ӱ%"7�@�g�O��wV���y����
����L�ų8�A�[���<S@�}�S��0�3�t�D���~��wE������1_� /�����iS�`A� �.-�W'�O�O�=(���@�G�H�����`�}>��^���U�n+B�+׸ś�R�Z��Ծ:E���\Tv��Z��H�VWhT�0CǕ((v/O�I D�ڻ\G�#(��N�) 1`u��"�_ڈB�2�jlۧ9�����@I	{�Nc�$Y.2���Vw��h�+8�������ã�e�/���hү�v�޴����nn�����BY)�M�Fk��[��c����������O��V����T�[;��y�2�Q(;��b����=�k���z�c�^ ƣ���Q(Ԭ�lي��?��.=F΀U!i�Ut<���H��T�b'�Il�{Ҝ��D�W�(Z�$��m�B�ߐq��>+�VR�5�g ������2N�t����<�֖�0�0�׭?����FDZ]�7�.x�l�����M��-_nC�����!0�Y���LBX�:�X���3�T|F�*i0K�����$7�dl�"��Ѽ.v 6�Xe����H�V|��z�� _��I��h�/�����O�!��s��}�*��6}���]�"�[���Pr�]�.��������o�
<������!tx�U�%�r�T
��e���A�힁FQA�u����o���2
rDj�
�o2���]�l�r`GӔ�"q�U}X9��Y�*4����xw�^�&m�� ����eb�Y�AP)����j�(Ћ�q�RJC8`���/q��%�z*`\#����WD���2�W���
�\5��Y��Ny�RQi?�^8И�V��ۥ\=�@�g�S�O{�����&p����Cy��T�ߵ b���	�E�E�d�ҩ��N`s[��JO>}��ei[Q�`)��x"m���By �&�:'8�[4��UUkL0�a��5��&H�C�ǁRH�a,�m�nJ�Ӈq�I3{��]"�a��t��a�p��������8�� �d��F�n�ֆm���L����\�VR��C�c,x�"�xyl��L��/R<���6l܃C��FJ<:KvV��8�.$`m��/��|y���8��Gskq�o�1�V'���T�Y<���~7�0��v�2ʅ~�p���A���9	�;&�"�MMލ�|_!9j���n��nJ��+�=Kk�A���C�v�=��>�*�\�F��x�G����h� �g@Y��\�><O�Sަ�N�Hq�(I\r'�%� �Nm���-�ȱeÌS=��[��aVPxȸ����b ����� :�U)ï�]�.?�~kf�Y��n��1#��0r,5@)\á���F�tIW>���w���&�-�x	����e/~�� �p�9w�`����BU�{CV3"ƕ��P�a��{�;�H]ڕ�F>�/$�8#fw1w)�{�v��ݮ~����>���א��/X�U�� ��CO��JC--�HU�_�\��;�p7�Q�6U��%G;]~YM����9�U�#��b�ި�Hw�[b�d��� �)&�Խ8�U�����+A�Ա7e��
�:_�����q�[�#�Y��f�5���9��L�����]��jN	Gu[�xom�	�����hm��c�[��M������_��|��M�D�Ӆ����e$ M�
ז#���T�F�،P�<�,��(�}(�?֐�[~E! Z�o��l;{�[-�(�l�\Y�빭rrs%�{%+�^!��q=y�c���o�gs1���B.zX7�
�����֓��aЁpp�\����(���WzE���L����<_�)	�P�c�Tk,3i&' z��1)�~���2��%-ϙ]G]�u�C��ˤ�¸sb@L�k��F���= ��bT��ǈ{���(�s#'�(vӶ#��8�Q1j]��q��jؿ��`Y�u��]�gѹ�;CGtuj���B�j�,��;?�V?=.l �`&uӫ�̠Y5��q�{b���O���.���[�|�fP�4.O*Ĩt��+\X���.Y��
"8���cy�Q�Z-�#��0���&8]"칈�Ƈ�SH�)���6����_�;�@\��������� u�-�B�ԃ,��.��kY�����'x,Ȑ�"�^�m8N���?�]��'o&Z����D�Du]L5�?�w��fh��uQ�F�W��-;V᥿��ץ�0�s!�m��d_�����*m���I�0��-y�|����$[#�D[�cE92_�� '4�S��N�=����W�@V�����d����ȭ�n�b��f�$��/��I������|"�JP��,�Es>�D�٥#���:}�F8�Ņ������w��Y,W�ƚ`��#).Fp�.����V��:	��5c	yt���{��WGi"�%51=:x�^5�8��1����h��ֳ����S&�%���`�d���<@�:����\���:�@t�8m~H��[ǳ�a�pj��q������D� ua���T@���F�����t�Ϙ+!^n��������N�۱��S�I+Y��.ֺ:�)�_Z������8tm�YY��
 ��.�g2 W�ZR��r����K觫T�䮛��u(e���i�<]ġ�̤tI�g+I>f݃N��6����'��3�__���I���u~��zH�I8Q[#,)0�W*�!^�.=�L��8m7ZZ���O���D@� ! W|�̨Ù}@Q�h�f1,�2^h�AҠc�&�2�d��n��'6ւ�(y{�0�5:�/���Ë<5z5b�����a�!�f�z� e|VK�g���W
R��P#�o:�A(B'H��,���6��Z����Wͱi�Ε�@�b��-��Uxn�vOS?jr6w�Yr%��xz���),��y˩|�H0�)v̳T��*%�C���"<��4���W�釢�X�����8�9}���˾kx6�`�lԓ�&`��@䖨����n&	Y;l����׌ߜ����JbȎ��(63Gי�T7�ã��`Ln�
����
�$2-�:�(��P4�!��!���R�%������m��-��9���x�WW�����)�7u�У[���=Df$Ӹ��&�L?��n�pGH~��u��� Q>�D�X�V~l��
��;G�§hǓ-y�l�����%^ �bѨ���>��Yl�ru�M��:�:g�W��8-/�P_(�8���fFp����6r�
�L�Z%�9�l��z�c H؉rm�2T�˶(غΝ*���7�6'
��:�bI��C��y�Z�"Y�h�չS�:�[K�/32�b���I�ə_I����]Q������
��[����F�!Ǝ5��40�+��Q�ӯv��C-o�!�(�M$����a�uka��6�����Y�����2'�A�1L�=�n�!���=��Z�F����*��V.���}o��RdQ��N^�P������_;6�r���2)��W��_� K�4��޿ٙ��3_D���D*
�y����G��o  �Q���;,ẍ̨��� f�Y �U|h�Ql�N��΀��j\p�(���h]�j��bN)0�d��)mH�|�ZaUW��OȜ ^���B8�r=#c���3:23(�����!i���H�y}�mi�Dձ��b���	�;���!�92�|���N<�~����G�f���#��~�O�3o��2��0t�J���=�`	/�рj:��V���o���N���r���c�?S�@F�_C�v~����=����k!)I���� �e�p�Q.�,0���Qb�S�3\z43io�D��;wЩ1#F�ҥ[�+ʢ=��M�;*R/ b4{	��	�$	�B��.��{����`�;r�RMfh��^t��qL�X�����F]�W��l�%m��ؙqL�F=�)Q��k^���Cs�fw�5@"��{}��߼����W�yRQ�.�!��$��U[���9�H�
�}��d��GDT�L�;:O�99�]�&����p$(p�;v�w˿";�Æ����Qk84z3Ȭ ������U"����O(n��}EӅz`�F�b����j��I�t��A�
�p�o6ϊ��_�׌&���i����<���.�{u$&���KGy���ۮ�n�ۨO�ʖ���o4���*��Ϣ�ިs�X���������)	����T@��HG���*��u��#{�h�N�S�A�0�N���Z�B�A��c����q�������SR����'��ɐ�����!2_�@9��j$�Ӣ�d!u��5���$N�h�q�{�_��d>< �T���n���K���4��wxm)��	�`=)�e�\z*�{C�d|H�'t.i �?E�M�u��k���V*�^�uA�]#��v���0�ƥ
!��̀l{Ρ�k��~iO�<
b�"�q0��>����-X��B����V(�ow�s��E���^ �JSw`��@(�h'̑l|F�G�|�7����P�MƔ�P.������ꃿ�/�T��y:�ie�e�?���z��� �7U��^y'�X$�=� L{s��>�<�����h�꒭s�a�X��F��3��aE�ϳM}����5BM7zx]N�7;�Z�WsR�6�ﴢ�ZT���\�SE����� �Ad��ku� �@1K��M��^`�;} �+W�ƾ���0�#�l��De����w},Nv���$�����C��T^�4���pa�jBB�N��7�*gQm�D�n�q�}r~�#+`�a��#!]bX�����IS����n2k�����kJ�ϕ��
�V������e��d��+P"U]��t�8���%g�so"f�:�6��� �����2N���v}5�JY�qj?�1YuZ��Jf�D����yrcIWJ�A\��sܮ��.��)�E޲e�X`��"��� ��4e�an=}����C1�̯)�����gr�R�wuMOS��
�)�ԣ�u#2�B���_�}´�(Ș%��I/��)��]`;�e`���m�<@��d��8Nꘀ�;��KR�z,��Cn��tM���K߶a���Lr�CdX�&&$������7�����<C����[JR�'�}{x��x^j���	����S�#$d4�U<(��$��߱���D_���>�t����)�M��\�����~�P�?�R�a�,�����s@�.i��̲Y ���c��~��D����:h"���u����ſ�bN�>2���w�n[���U�C�[!^P������ 4a[�=�͘�2���oVٳ�V|��	 I?,f�_:�6D�-f��D,�:KjD�e��:���*]LU+wh�Ћ����`�mNT�!�SZ*\7��H�ԛ�y��zat��!�,O�G���UB��F�C�5*�mI�<|��(S<���Aҷ�g�`#��ʲ>�vQ�gclc�٠~Y���96��n�f�������c�=�߿7�BқL�����\�lE�6۱���J�v��!xs��1FnW)�����/�H<8Q^yЊ�q-m&�b/��4)���NTX.��dֻ|T��pe��v���l)'WvQ���m�AsA�w>�� �$��t\�Mۺp_t�h`���ٖ$:��R�/u�����W�F~!�P�Q���,��e<h�6�9�ѡ.��J�Y������O�nڑ��u�T�u&lHk�2j�DF�3{Hl!�1w#�)��]��I`�M)� w�Ê�d�	8�2�T�p#���DU�;H�#�*�z#8i�: 
�{�x��<�T�ޟ��b��[��W5��u&N�>���ƒo��l���a�'�/�Vo/ҏ�(H�[0�
��(���-E&ڇ�ݠm�	M��A�(C�k�JcƠ>��m�2���I�aߤ6|+�Mư���*�3׌Q&?��}����d9>��J��xC�\�<D��ئ�b�xX� ��gB�NP���'�C]�آΧ�Tz��`�e�i<�"GDXtgY�~Է���S��sE��>Z���d\Lh�(��ϑm��gVN�t��+>o�Ԑ�<�ۖ�h0���c���R���M��/��:]���P�˓>��`aQ�#�j�M���g�0�Y�x3��w;qI�ș��d��Q�iT�6�,�1r���;K�(���Ą>�~�[t�Ͱ�@���ⷶm�@A�)�e K��%�QW	+�K��ӵ+"�tNp��!x�A��`�+A�!�s|M�}w�6�ah�Ԗ�q+�-�?�fnr���w����0̒���D1K�iy��e�]� _@ *N����6�5G$��}�M��P/�	���o[W¶(Sz�r�b��ҢN�h�mH����X���s���W���v�ͥ��~k_��S����E.x$�Όj$��Ǿ�<U8·lH��9�J�ca�;1�րy���nţ\WN�U��^��0��1>��p�������vN���PZ]�H�������#�-��fb���+K�oI���1e�̋ǘ�%�i�5��)n�O���Ka"V���n�����5c��*OV���= �<LLŞ�On�r���F�M��#�K&9�A����c'�³oOb�V��rH2��\��h�g�mm��S���$覭x�y�e��V
��H]"*u_��:�\?u�У"w�R9S��!f�Z�nF�*p
�����j��1�J4V�
{�9;.6ҼO��WU{ҭ����w<<-6��ԃݢ��$hF�y �Vy%�7M�羥�4�1���%�U$K���J�,�x��(���v�������� ��ص+��N�EGAw��Z�n�6`A+&֋G��#�~{ǘ�̸��w���t���:�",�<Hs��_�H���d���k��_^LC��Lsr�YKC�hM$R��ik!e��zLvg��a�Hχ�A@	�9:A2��O>|T�Դ�t�6�����Q,K7��L�7�h��� p��t�Y��ώ��nw\�v�^� Y�N!9q���1��_5a'�Mk&��6�(1+�����V�{Q��ca�j��6�r�T!R�q��UHy�9���P8��ƛQ�[��',�L9��)0=j#�'>���>����\+*Q��ʖ�rR��W��+Mx����dN��aM9=�����q�w^�v�A���Zs�`�ݒooW�#ќ]q����N�3��+���"��,�@���¡�1��!�צ�B�eȀ�~J�I�*��?����(�/i�C8�x�yn�Z�.������5|�8�a��g>  @��]%����W��J�w �sd���@�HS��بvp���f�Ir�}h�y=���]��dV�-�=�; ���gBqκ�gn>O������4Cr�p
��&"�e2[`]`�M	|v-��ɫ�p�gf�+n ��D����15������B����x5,������ZηH��Po��|�!���$z�j_��mc
�.Y!	���U�D��J�U�ڞ��d)w6	^��0�bQ��j)FD�������M[G���%���g�;���S'&���5J�|��,O�O~�X���Mˑ��{QQy�բR:ddw��n�n�R'�tP�j¥����=e��컕�הӲ�8�D��}�\�L���+�V%�Si�rU^�1�_�t���-��C�樓���gG�Wp|��7 �5������n���w{�R+��w�h�aVs�6Ua�AC�{x�;�X!���S:�5����"L�ށ>�M���c����������F%s���h]M��>���Ƕ��U���&x\7utą��f.8��nW�k��=��= 45��/�W�JSa�y9������	*b���G�`�s
8<��kߙЪP��b �]���p�urZ�7n#c�ޮ�OLa���x�6m�&o�*�a�u��G)*�jF\r�+CTB	��=�n�M�6���M���~�ib�x�R����:\�A(ct��H�������@�rɢC��,�PW�����t�x|
���+|���Op5vkY�I�jX�*��W�/>�Ζ��yD9��>N
A���]6LZpA���R�Չ����	x�Q��'0d]w���H�N���W� �*���25�i�zj��%eK4�@v�k��>D
+J����T��K� ����??���l�A��o�ȆjlA�$��aWeM7�c���o=�l#Tt���8��(a���������x�ʉi�-3r�32ˑ������ �M���[끭ۙb��'���{��)�~/��^���Փ���ߘU����v{�P��z�W?�-���(o�i���p�G�v���.
���Oɩ�$���Xkdy�� m9��P]���A�H/U�Y�?|����rwt���G���z�����Y�4����W4%��f�hN���1��I�%(وBP.d��A*q�>��_^�������R�72�یȨ�C�o���#;�9sece�W�B[�]S�g�>²�XI�~�93�B��$���?���1����ע[�U�kyl}I���MM�	�w���-���)��?o�w|V�ڲ����L��Mu��qx���F�1��𪡝߯��Ti0��
2����������W��G��^{����H��i�6���(a�9Rpǝ���86֠��{�����7�=��X�W$��
h`�x��U���Xn�XI�����������!t$`�ڻ\���$��ٸ�tn>	 ��ab��"=���v�u����k�z�vj����CJ�����ԈҨ,����n��܆����+�������IɻX8�|�G>�a��~��!�m%��W�e�s���]���І@��I�f�kgQ��f��B ��ؘ�÷�o�]���tJ���iP�q���[�ǡ�2
��@���?*m.�*�@a����:�q��vi}�'��M�l!S�rݥ�|��������~�a}�0��o�O!�"�%]Z� ���>%�ļv�%���������o|q����o�,�"�P�@������1J��W��iR��V�_i��P%�I@s���d�p�s��0��v�}0���2�Ɲ����rz�V�����+�oߞj�z,T�d0�HS�����l�D*�F��)tx�҅B�����ʽ\S����?U��R��);̾�_88a�I/�/�qN�מ,V�V<����-7ՙ�/���Q�$��,[���6�fߜ�i.��ٲ\�5a�R[9�/�}�%��I~�6�w��Ki٩�8���JS�4ṹ|�.���=��y=@�W{RF+�	'y[�$_?壦�!*o��s����)�,�&'����=������A��[=��Ҫ���/G��.7.��76v���'j��
�>�����	�dm.��j��M���(�I���P�S���Y洼����'����}�U�C�F;	u��%�قl����0%d�\����8�2�O��z��>�U���]��e����.�{hm��z�������Co�Ͼ��;@�B�������A��['���2�\&֐J����]�����+�v� I������6�<��< '�d���O]=���C����A��5�e~��/�J�}�>]���}��M�(K��	���$��Қ�m�d{��ߩ�J3�Ϫk����\����ZR��ru�I����)��%�������I��=�eZ��}m�+�s����r\�1��׈u=�!G�ҕuj��TC�h��A����3|O���T�ݑ�#zP�2rT�{�;��_d����a��Mثg����کdb}�U3C"����� ���9bn��6Z{(���_3�݇��'����|)P�6�Ư�@��h2�������?�"������D����Z��KM�]�Y�E^�o����إ�XA�V:%�����n��np�Om}ή[�įq�y&1V�˄^$��B�Pmx2a}�#hV;�C�9M�Țd�t�J�0r�"�Ꙟ����������&� yM���r�����L��~��ϒ���U�;?X[C��25�hu`N��=���!��q�� ����$_���ƈ�}�c����Ƙ�X��ɥ�T�*�����u���ºu�p�z�6�9��S�% �l��D岙L��9���%�W��|�!�Ā���"&��&��O����G'|ŅWR�[�k�JP��_� �/v� ���I.�ʞ7�D�R�=#�����W�k[��89��;��e��W�b��#a�i�<������,!�6p���ӣ�.;���Ұs\߇���e��	H���F���uNtF��/�R�ִ��Q�u��h_�!���B�;=����vv�gLh�������N��x�8�T�����#S9�MR�w�e����nV����V�G��tYܫ�vp':9W���*W�-����U���y(	Җ��4�p�gX�Y��O�٣q{�;���6�U _���Wʓ�ZGۧtZ�(�x�#At� ]]�h5��z�ARe���C��]�O�5�8u��M�n����n�
�x�pΗ-Q��?�^w }���,���ZU�<j)XV	�2�y_�0�^s�	�Hr��H��Yˊ9�"�o=�W��"���=�ty ۴7�@���]�tσ��;W�^�f���P�6���J1aG[�H_+�����
)�z-�Qg��l�x{Xn�d>M��!�LpOw,A~�����懙�tWYKON������L��W�!�'�Tޟf_��-���p�J�H`If���_��̆���F4Jܱ������jzg����,���������X�0�X��Q7���Ǯkq����8ΐ|�_N���bjnD��Y�`���	�3Z;r^�e�R���Y�zҶ��۵��Ү���n� Q���<*��ob�a�C��������OѾI�2��&�:9@I���&�og��f/_��tcȞ~C�	ה����rQ���0a����U�eY�?��|g��5߾���)c޺AME�Q�6����gJ$gim=����%!:[#��q5;���4��b�Q9��i�R/�i�p�����{�y%>ȯ:��G�s���eҍ����HdƄ��yr�Lu���e
6�/���~�fa�4�z�P�'�Э�R��?��5�D��m�שJXj��	E�pvX���p�|�o�4f8+j$�(t����e/Q�Zz���a�ɶ:G5�3��e�H��	7V�o�Փi+L�?CC�-���ƻ�<����Q��<0|�w˂�9컅�L��LN�Lm�B(R��A��z0&`���1���gҮ���R	��/|g��L<n����@�;�L�;Y������M���~i�3#�b�-w%�jtf��v�GBnL1��8��uQE/�E,9X�[�8�i��i( 8�rb���j�бb*z����H����
�-_��Kb.Ch�f:Nc��w�֠�+��9���{u�=5��Јi�)������!n���(�2#:x����0�VL�<�Q2��� t�<N�䂫��/E��E d�O;E������2op�w0n��{�hy%D��u9؜�]]R+o�7`�_�9iu��g���Fhn��?J�?G5癅q��Å"�c����?!�#�oy>
yC�.�-A��S������ݜ�Yp��B�K�-�,�Ds,;���1<ƻ�?����+B���?G��!�c���a \�D�KQbj��L�d��4���%ϊ?�c�_�d�!��ll�(LJdL[�B���@��"h�9��n٣��!"*t��j6C�/���'��'��H��_*����5k�e��i@�����A
�<�U���D)�Y�\ ��wB+^��8��&�z]X�A����h�d
���� ��Z�{'hҖ�H�"-�? ��[s�
0��:�ӬW���Ĳ������U�"ގ�*}���OM������r���znu}/!r���sLe��{���� �9"#ˈM��W���W��-紅/���m+NnF�<N!Z����u��$�ߡ�n B��-� G:�ӗ��A�Y��U��v�r;(��هCB��>��'��0����(�|�0��q��c�x�r��7i�f�a�[~�ӽ�0��m� �
��_�R��+}:��U/2^�|ȉ�s�Mw[�K�1���	�q0l�)��p�&��ԹM�
�W=ǳ-�O�c`�2h��|1��9P��*\�fc��ec�95�h+��;��m�.�G�t��� �R�ʻ~�K����j�b��6�m�Jfh<�?��#t��ۢ��´ ϸ����[�e��h��΂�6Cz-+m�r8l�i�{�O�k�����$u���H8Ij-���{�w/��8}�z�NBŜs�(h�����t�Bt�ڑ�r��W.��|�g{��.J��^���̩����8c�C�E1�X���-�N9^��'��X�n�^έC�(�Q
18���N��f�dnS0��eC��P�_(vDi���z&&�S�)
�V�%e��8f,9�wdʐ`��������[զwF��\��,�"�c����G�)$�퇫\uO�������*�<_Z��FrxR�����OǱ
u��Ch�5���⺑�K#�ע1M�@��V��yT��
62Ί�2��<����+jT��Ͻ��Zt�����y����茬��6�ۙG���Ó?���3E�������$����m�H�C�\���)�=�O Z�<-��t��P+�6���D����ͩ��;M���p��J�9M���Q��|�q�(G�s�P4���
����O�Ϥ��.�CN�����H�r�!����dw{��cW�������`�`mi/��o�B5t/�Xl}l���04h0�����0�3���Ah$ƴ��P��I����}*�����J�U���3�Qݢ�܋�~.���uس�����VXo���{��y��F�Ogv�n�M�����L�C�M���哣�H���/�:�F��,l�� ������A3�OkKc�}/�8
5�/�g�> AFP(U�bkhs�Vh��Z������!����4:����
���_ը����&�C�U,��^x��e>��v�6:?����}��-رJP�L����Y���|�a�V_�>%�Qi~-A=�i�rF���I��a( 3�F��/3��z5[��-UT,�V}����ߴ~�Yb����q�$|�	�ﳰ��
窶�R����$ئ{~$E3��\\
m�w|� �R��c��>�_�������u<�S�5��� R]hX��o���S#��4�+�ӌ�La���s�#`Uq��n�[,Z���]*&�ڣ����q�z�0�2�J�/p0�Ia_�k��$P��G	*\�.x��-2�8�nʌL���|��<�,=s�FCO�X�~in<�����$ {�I��H���G��5���~Za��� ?�M������C�Y�+2�$YT���襐rm�m(�˔v�|��_ڶ6ʂ��aS?n�ضB5M�sS_-G�VX��Q%�?~�5g-� �<� ���XŇK'�.8��	(-����2@�����9�[�U�h�Q�[ұ|�v�O�>�?<�ey���|"E~T(�/��'KP%�&їB�"�}��Ϳ�e�D�)í���
O�G<�K�8���ZQ��jj��W�|�w�M�r%�!�d�' A�Г�R 4�,�X����X�u,��Q�=���b[5���8D9�4ZY�<�z(#�1f����.L�ޜ1tĩ�D���H0��M�^lx��2K����$������0��6�3	�w�N+�O��UbĮjc�w�x���A�0�k�x�ry��Sb/ �w�>�/�f`Q����c�������^���cd��r嶪�)����N�N�{��G!%�γ�#`�잊qb��7��i��Pe��0�kj�J����:,����,��w8Ј�6�b���n6��Ċ@�lV��C�E�_B��3�W1��T)���h�̌&�d�_5�E����p��#^�C���lv;�(�x� ��ֆ�^5aY����A��0�¤���M.N���_����G�$��$�C�"Rm����>��`}�1mX@����g!|-�9�%�����Ȓ5|��>D1���+.�pܳ��G\=7��,�'�׬����g���d�����s��Q��U?1�	�X�0��7S�`h���,�P�����sT
�]~�r�z���|ϥh(��[8L�T�H�A}̰����x�`��[8���B����?�ۅ-6��0I�E�X�6pY���� v��;�[ )��1L�M��|���&L�7k�*3u�\/E����J�1�w�E(dH����"�a�7�� .�4`��<���ո�d�}�2N��$����kZͫ�E���Ɣ���"^%�n�7m{mڨ#'�$���>�)v;0�[!��}8����x�i�Q�����)ȑ{�QB>6r�H�� ^?JPtzu�����Ƅ霢/�	��*S64��A	�e���|��s���X��:�|�~+�ie�>�_��r'�=�U�Ήn��/{ta:@y)���d�Is/-��n�7��Z}Û1JBl���-�L�u�'Ԣ�0�t��&�|�^1 ����t��u��#�T�U��0����c!�������f=�C`�T�]�9P���*�ֈ-�	S�V��^� �9����SK��b�φZ�ܾ�2��&JW��ގ1�1���5.����Ȥ
?F{��γf����}���M�yY�Ѓc9 �u���RY �jTe�w���B�A�+��j�0%02��R�RBM�'�����D�)�^܅��zr�.�[L�m3�_��Gw����C|����X'|%��@��P^NԌc�����r��8�X�(ZHq#v��//�k�!�\�<�&�������E�����Kw��d��;��21R`J�7B��]D`���n`�Nl,�!g��8�*S�'m�N	���$;=6��=F��?��#)�zUt�t��nݏ�F�o�����-�$�}���w~�*θ��;�n�N8;ʓ6(��ᥫ%��[D�Kx�Rg�馪Gywj]��0�ʂW�1�|(�fI�~���S��ʼa^4.T�x��I�B��#�!c�(�ARm���%#��D� ?=��6K�@D�t���|�d�h�����9R�9��.<)�UmQ����9�z8~�
z�����/7���� �V�_Xy�`��h�G������ V�eEܽK �q���G����QEO<#�]Z����i��5j�QsG�������+m���#Ƈp	��֥e]ZijǕ�g�;��>""q�%'��-���Faš���g�@�B7� ;��X��%���ø�9b��n����/j��M����Dػ�C��:V�����0��2+�r�i��-9����{ߍ�o*ɮI� U#c����l�	�5���S����$쏞�Hy=i�`˔���>ޣ�v��/���1����³�o3/q���yY��$l���X�	E��Ss�
�������K�W���8V99Ŝ�1����#L/��ⶉ(�΍@p�����٘�"����:̏w%�-�ri���K͂�W^H��-��P��e/�<˵��`+&'F�t�4Rr:"��c��C`�!�0q�Ee� B��r�Z��ύ�=�Tϧ頻� �t�����<�k���-�jY����4��PJ#]����'u$~*�A醊��%�:�j��G�i�����dh^m�ߴi��p��v?a1���������8*o~�B`���S�\S���^v��$�~����g2U9�c�J�iȄT%�m�;kӓ��(�f�|��[	BH74��Ƕ@�--	��7��:zy�,�Ћ����N�[�<�L)U��eI�	6��imN,�:Fف��c�Xإ�>���a~qyT_b��C� ��@��v$A)"����i4��G���duЧ�3�G�Y��ζ�?S��P ?R�ƺ�:�R�iǋ�����hqQTq������X��Xak���c$�/�e�F�n��1����Ym^TF�^вAx���w�$M�b�?ˈ1
�ҕ���b�;*�PT��	�����Te<<0+'H?Y"�xn�?�j���U�� S^Q�O<ߏy����Ժ�,����F^�Ϊ�Y�/=��6۷����� ��8�`�di!�n�����)�c l;�F��
a<��.]N���uІ�4�
y��mf)�W[��c7�� !��V�
�
<Tn�T�	���en2�$K=-(S�JQV��l�V��?4DF9`�0�����{���!.��\�o���+��Id��f����ůd�����K7�lr�l��{�ƒ��^G:'��r;H^�D$16Gڗ�T��!a, .���Y���g�ٺ���+$O�VԎ�T`f~�$N���ſ�v$�l���w�ɨ�<��	U	H/���tQ,!a�yn?> q%��vV���.��&�Ɨ�i�Cp����Hk�Pۙ�R:0�	7Ót���q$I����_��������-����8I`:��׻S�.���ސ���j��;����]��,t:E�.qO�8'�%2�7	TqJ�#�0D���8VU .B:v���f���\��D�{����@{��HI�#/��fΎ����v�W]#�J�R�@q�3|G۴{>(����x�8�������D��!��^��\�"D~G<��u�|�p���(�>/.'��7"|�)�M����-�}��}+<����a#�gkď���k7���ɊWG.�`2U�~Ć22���oo�����F�K�t
����ԉ� q߇������r_�?��R=m������u�e�٪��k��a���C\'!y/�i��΄���.5�l�ʧ�ųs�{��V�>/T�JA�8)TS�裱�c$���s�>2f�a�4P8����5�Nr���R�o�����2I]����v�_��i�[	�,д�0�Ut����Cc�����C%p�׭��fn��.d��2�}��<Q��i�k]����#ρ�u�M��b�W�(o�\:�>�}|?��tξ��Ss�sS>��;�~6m��ǅN�!EK``�u�-�	Y��
�"�b�Fs�Hs���.���q�r�DSm[�κ��=lu��ј�jة�i^=�7lA�S��jQ��g!8<X_&���[Xm#4�n�}T���/#�֣�?I�zV��'hs�|z�`H�t�60�z�r7��@	�J
 �3���:��l|~9�&�����ҥ뚥����v�/���ɕ�u�o���\��a�;o� �ԭ��Cѫp�M=I�-W}�n=�����F�8V��H��|��R�Rpf��n��`���;o=��]�*a�7���t5��ؙU$�;�|U�yG�"Qr6��*�4�}�3|�S={^�1�����I4�#-M�U�!���$?����w�I[���� ��1��?� �dM�p'&:զ���14�U2���4ך����yr},�}�>�O;m��TC몢� �y�3y迵)��~n���8I��{�b�}m�,�N�{W�Tc��>���/�3�YvC\|&�#(�Rg�G�+18�G�	3��5Ȥ[�[��Se.~'�2@YnO-�v��r�86��L��cпѠ�.�&(B�]���l�t�M�`/[� ����?����f�'��1N&�/!��!c|�
k��[V('�V�v�$��L/1|��м�4I���t��1��!��yo�\o�HMi[�(�ϸFyr~v6dxSؒ���O��I�4��]�/m��8��՜}h��M�}��M���e��!U.M�;��C(�=yn�MX������G�tn+(�T���F}�|lK߸��)�%c��g�Wf��N�,�7��M��e�t���!kD[�X��:�6��2�٤�`�?��O�-*��PKg�;��rDI�41XXci�St�gc|��NzJX���7��C"BiټZ�a3�����f>�a�o��h�������#���A�⅙ ��J�[
(����pW�F�,5��ء�[\�Vr��t;�&!����̰�'�a��.!M��g��E��{#q+�2��r�@۠�ĸ�lxuʮC� �
�k�����U���K�+��Aȝ:�Y���mq���3�0?��A�*E%zg ���ȣo���R�D�F�n����dM�[�6C[����IȌa�d�aV-���I��"��C�)F��׶)�Y����|ʹ1}�DY�i��\�9��+��ᜡ�;i�M�Vyi�ɓ�/$�ɒQ�b�G��b�����QNi�#���%?�!Ҏ�����L�	�ٸS
��>n���Ǽ$Fo���ZP��묧>�Ҷ~`f��eБ�d��j5��39r'/�΅F���X�;�M8�L3 �����L���26��<Z��L��#�P��_�w���9������Yp�(7Jx�_��h�R�L�ځd-mE��v�x�%h���E3	����QX��6-�6��"E
�F�l&�1��H�"p��4�: �i�D�u��.���Ń¡H�M�?���1<`�"�.���+�F���B��� �hPC�l����0�&�sM�w��z��:��R����p�	�l�C�ܗO�4 �9��E��q�N*�����ґ�&/v$n$- ����.'�=8�Su����Y�|8��]�`�M�����}�aY�r� � aM����!|0��]��g(�q:܊6�q��q�������Ad ���d�*)�h�@��Լ:e:_�SW�J���:�Gs��`�rNh�cJ�+�Z���f�+����L܎����C����ڜӡ��<�2�ג+��4��7�W6:�t�-�ev�'�-���o�%��z���t<� ����+%;�I�0��M�z�ZL0��������]��-how��U��t�oy���_)�«J(��c0�����&*W���&�̆��D�U��P�X:���#Lkb!���M�Oս�*�P��	o�b�����s�b5�pp��0{v�0���/O�%�e#
I�f��bP��>���o�ً0֛��`\o�5����D���3�la^��<j(k��Q�G;J<����K����Ȳ���E�"қ����ɏ&M�HC������ѫ8Z��@ �H�j%5k�?D5%>z����ա�,��Q��Dl�BؽR�F�󥋔���|�-� �|L��R��l��Y�"�=�#/|�X�o�	哽;� ��E�gB�p�-���#O�(Q8���@2��5]=Bk'�J�"sD4�:/ps(�]2K������/�!7�J��T'*�j�\Gf�4?�᤿tX]4lt��s'�\�8���7M��$d��ڏa��B�y�GÀi�A
,���u1۠"j�,�cf����Y�\yv����Kyy��9m%i��O]y�ܳص�ey� ���.v�f��s����׳���N"�s��D�$�=���'����Uݬ���it��I�w ������jn�!Cc�l{$�ۗY���>.�$��Ow��w�`��r)),e]�$C����{(u�_����2�4h�x�n������k�6�jV��������50��r}r�B�O���H����N!q��9�#�A�&�עw���%n��{	���2
O3Y������;Щ@Q8�m,PQb�,�?_QfEJL���3���)qN��_����>K��3x�t&>��KV���?cmKzw�7�Q��cp��R����(`�%4�9��?e�T���c>�Pi��$��|�'L`����{�YEP뒍���������BE���f w�\ʆ�$SP��� �,�A�#�&�B�Jp�N����MΎ����yC�i�������$a�L$�H�_�Wu��hQʑ��'pG~����o�}�!�v��S�΄GX��D~�w�U�/ox��VO�,�ܠ�u�l
P�2Q��H
;@a��>]�� ��#u���t�7�p�����9%xQw9�XG�ʢZu�nA�/-��ɂ.��A>��n�Ո;�s����g}�ص v�{�9P��'��.�c��F"�FX�2��hT��]���Ǽ�S�B�n��� �d�P�,�l��{M��\s��0=�Qc���(y˭��b �q��UX�;&=���3�*{[�`�	��c���>�v)V���V֬?�{���5����F��.UHL{�V%��&6N��p�4?E�>x�`�TM���q�\��:<����p�a᷏Q�χC�n��'8���,����O�Ym:!�רV��o�.�-ڂu5!�ſ/�(�R�R�F�'k�W�+zP��r����"Dt���<���ǃ�Q����s�*�C��{�]�%��F[�=r�W{��Ϟ�c	O.>�tp�q�Ū�l�w�/^H@�ύ�f��vϵx�dx���W��6�&#����H��U����� ���t�:�R�]�r�f��,!�"���N .��/�-����Y}�1?��l�f���`�yA�",}���!ƚe�il�qf���DS�J�� L�/j�aM�L�Q�Ȅ~k� /R�l+p���[}A��\7=�D^as��ף�W�߸&7��a��`�$c��lj������-���3��[Е�2��b3�wן�5I�g�{'iXU���j��/��w��'���
��t�(�B��=��\���I(W6q!���[ͬ�_�-�I%� ���+�[��;^6k�f����Ms�%��ԟ�W�u��e|�ڐ*�f�J��	�{��Π�;Q��v�
��a ����$<���)�2?�`A��pfݳ1�:q�`�p�B���������Y/a�P�OP4��A��L�\v��Ďs�<�h��{ȵL���n3ۭg����S����7�m :���!�ƈW�K�2�nщ�7N��M�T�*��ؘ�� �����ò��ņ��;1�t��N�mx7�@\Io�v�>H�M�_��u��P��ق�Mȶ:5�J�����4jZ� �l�>���;�[f�#3}2{+���� ��C<`����PC���eoA-���jiK����2=A�%C�P���Nj0)��#�7�5q�e�*�O՛s�vJv��a��c�p�7�'�#m�c��E�Ɣ�܉��U@Bo���ps��������E�0K�T6�����u{����/�f�gC��K;�W������`R��Q���Q�`����As��;M�!QK�NUKO��o�=�x���.7$g��3�� Н˃83S���6�co�r���Z���C㲐!fA�ݭ�������:##>4��#�4��"'��Z�yKl���ܴ�y+"!�3������h5L���Z	�sZl�1�*����-IX����񎼲�:��r+� ��F��=c�ۋ��֋o!b�#�!�U���c��B|��,"�b��1ëE� q���7�ޭ<F�-`������
�'�=��,�Vi�*E�fP�QH&�%�1�%6�
&3=j�;.llq�*m��}{P~�����6����}S�<`�[i�N��g�����0�Ze��9b���W�0U^��%,c�6}-�~Tn'�������W��>���R�Mۣi,�ǩ���VF������@��i��947t��	�aw�ٰ�#�a�q��8 ĊV�is���xi/*>��XcPL �m��4聆��!$w�C����ExO��,�[g}}�3F[����C)fuR��`��x��O	�&�ۡ!��?ZMn�J��&-0�쪰�.*5�/�	���� ���%r<������ԧJ��q�;�k�_O��%�s��q��.Ѕ�jT=<#�ʭ�����E�g�p��}��0A���7�ڑ(�6��]GD�%�Q0��t��o/���.-����c�ݤ�֭����Na�)~P�z���yN�-�G	����F�M�P�&TlD�����N��:��dA>oQ�e�2bJ������y৥�}��j�d���S��<F�B�̲���o�c��a��yB�&+85�4٪l~��=~�#�W#��H	Y+ߵ�
)�4�tĜu���x�h�0�݄>�j�eZų��ǋ�k�h[�:5��`)������՗��k��Q��ڒ��|:C]@����#�"V�ʌ2FɈm���.��qJB7��~Cl䎸�d��؈�у㼭���T��l�����]�'	q_(͛H�є'��\q���_P���YZT�����?ds�om�F��O".bp�=���^-�L}�n,�]A!B��'�!f�`�~���O���D�Na,�π(� N(7�3q�t����(��{{hIc����)�; <��2皁+�7͸G��o��7��I?ڄ��#��oӧ�s5�v|�-i�*�+�)����}lD�0�1�&�2J�^�����h���z�8G�πc��X�H�9v��c�e�D��.���i�຀�R6*,�A~ ��.�1���pb�U#2�|￉��3Ս�Z��+�,����H���j��t�b&�?�f&(�{;/�yi�.|�#;"���3��󩣢���2��a�l^Є���v!b�QN���z�igV�L��5���O��';�6���.j�^t�\0X���~ۈ�kI\�i.��{%���r���-) ��`6��Qcg0���J�*A�T����p(�:9t��a�KL�*I�-l`&6��6��U�W�P����yE�� -��+I�M�����Y�vB%}ֵM�K��2K�WBMX�3m�׼S��k����n���[C�k%�:��X����M�������j�-[:�sGbt<����𪖚�cx=˅y�,0��Wq�؀�'/�Yd�?|�YIa��Ϋix��1W���>w<Y6����7� jM�?�Z�&�y����8���6��Vg��?�G����͜�X�ٳ�8��f	�JB��S@�W�e8�C��勆�y>�Nn-�c4lP�����S���rQ��@x\�V�)�]�?�/�D�M<%}ڸ���P���~Ɉ.R�^pc<���~{��^��J�0�������.�[�-3P���*t�I������`x��pg?W�V��),����1��A��X�v�|W��}�m	�ۤe=����⏷_#\�@%�G� HX�X�)�1���L͏K�<�)a����Q��R� �%c���;��M����+��	þ%`��J��of28�WS�pOW��n�
nu�`n���:`�K���j9���{K)��n������(��h��,Wv��5͹��1nr��Vo�a���Vj9�Y�ƈ�	|�YJ�}��Y�+5R�f��q��y��괶*o�EO�<�P����TV_�n3��u?$IN��
%VC�񟄤�vfj����ŎH��DR��LQE��Y�E�ʠ^[�D�ʅ=}�N8敜���>��Xi�Ǐ�������������p��^Q��ݿeiR̘RW@�G�녇"�&����:Qe)��j�ro�6��;�W��9/�A�bÀȪ��D]�����Qf ��)��|ſq^Vu����Ml�_�S�ǫ����h#�p�A;�]f��K�@���T"���KY��!��{젵��"ݎ8l��"�&�lcݺ����qÅ#*F�g/bBJ�� ����b��w( �X`��b���w��º�5�S_�b�IfP��βv\�{�&��5���~�f���{������"�W�rU����D.���h�*ꅵP��1xsT��	\��@�PIe���ym4F\��#���x:�޶< K��Dp�
,k�5�{(��/��M�Mz�\����0'�gh��jP͛���$N�Su6ST�$�Z�~�E���Gm_�;_���IΤ��M%�x<PV2�� U����2�5Ӝ�7Pc�
;�����'E�D����^��)��VI<�j?y�i>�^��H����|!y4�k-�F����Ú��X���UT�f
oeZ���#���ֈ�m��@̰��S��^��W�S;t|Su'�ꇲz�'��5�mˤ� ЀX�nլ3����������E�$/����~�VUQ�| N���盍��wH샷��������4��;��%�s�`if����O���:����O���;�}r�N��c�����#u�,S�釹19�z�M�H����:|B�.}�4x{���h����|�[үk:���͉=��K�d�=T���}��c��MϮI��PD��͆�}�������0W���/��� 蕴��T��Ա���.,�M���	�0�����"�(��}�Q���!f�ո��JA�<2wl��՚��9�N�}��i�����;�F���#t�pP ���C�O�ne��_'Y����_x�K����e����`���_�щ���`�:H��}�̍���\F�nl�U}�n�7Kq"�fq�s)n_���_��IU�)��nև�!� ��v^fr��0[�)9�u"�}��pm��L�6h��b+�$��]��"bEN#K��1�6ˑ�����TݨrP�=@�T�מ,�T۫b*/ı�je�9�a!�as9FB��(�oa��x��٤����f��Ҧ+�j�ư�v�BZ��G����2:.��f|���Q^���m�X�j�l�M��J0AL�}�lv�'��f(�9��{h������s&ai<�!��m��U�m�;�W-}�<&� |��/O>A�	�U�\���Ǳ���S!���S���w��Q�=��`��{�O�"���Qs�c7�
��7�cc�F	3�M@-D�,���DA��Z��'�6�6Se��A��w�[�R�m�320���p�D!�H��-(*f�p�*9_
��YF{�ŀN號#(+�2�P��ě�a�΢U1����/�`dB���y0�2�R�6o�2n>�\$߻/Eo{���{��f����+�c�W�:Y����Gq�NG�#��m�����2�&ڞ�k��wS�� �X�z�xO�ew�^a�Sm�>v��kʅ��3�5��Wx�:��%�o�RNh�����+����ǵ�����lg�i�p���K�cx�b+�����[+ξo�3�/���v9X�V�@���Ĺ�O{�հ�b���.�ʒ<�Nbh��G�M�>itk/t&u�=��sv�
�<�P���ر�'!����^Si����t%�]�p��
��H�����w�El�����ac@��g��]���c��Ә��,���l�2I���zwt����uƧ'�U~�8)V����A�hMH��T�����������&��Q����!TӕEk�	���\���ĕ�/?08v�I_���))��N{�h�G9�[P�n�#��O�s Ҥ��RcEq�k/t��a��>���\�E��j����*t~�հ��-3�|*�͡��Rv�	�b���Sd+
N���+��:�^�I8��$oES�Oˏ!�G�u����a�#ح個���p�ω�hinα�9`ݸP3�;��4~�_k����e�
��;g.,�e�(3�Y��N$��)���&�z��t[O����c�YF[�J��&҃T`�8ވ����[�%&���l���t��v��� 8���ͅ׭
�@��E�̇����绽<g� �z�c��ʐ�@ʏ�<��{��9U\������d|��Y�x��a�(g''�$��~+61 ��h���[W�g��+Z�د�6��Q����֖�~��Dgwk��=7�B�L�*C���۟=�,��b@(�4����LV\�J�{ZI>e#G��sw�j������w�&�PۢT���]�>����"�����)&���%��{2�����'_�K�Df&��J�Γ�A��-b_���[}
�	�8!��O}���${���f����v�")5��RЃ���n�kc��MK�WJr����Hax��ĉi����!מ�=��8��ѾQkX�i���LG��Q�Ԁx@Ti����^A���k�G�v���{��^������;h7�[�p�ߣ�I]���H��U�I�	�o����ә*,�bl�c��4��v����w
�{���s^���D�+-�?�Q�9���\F��RB&�v �}}E�6�1�����.zg�Jφw���=�C���!H6����x^�ܕ	�u(��X^1������S�,����DtF�ɝ<��[��	[��98�Da��ƛ �B�|�$�'����R�_�1�g���#�F0��yym,�h�uzj���0�/rI��@Ba3��TUrQK"Nl�����r�.V����������"Ä�4`���W!����f�6"�v�E��\�;�A�P��"��9 '�p/t�1|#�,�Z�]�&̫���J4(a��%;�;*��KJ�A= 	�%���W���
}蔧�I>�2��H�s�?�-���-��u_�2�Nm��J���-���$ԣYi�ݲ{sO��"��Vg��,�%��=8���V\`V����7�:�Ǉl���oF�;�w�I�%�H�j�zo��f`�qP�փl'� �����)����~�UѽL�z��]��#��c�e1��!�G��
�ܱ�X�CPۆ!���7l�p�����W=�IW �(�t˨óxtV���g�H�, �pk��K1���X �^�ձR��]>���j�/Iu�[���%'k-�����	eq��M殪��t�8U��ܳZВhv7�1OaA���X���1����3"��U��qx�Ĝѿ?(���k�]$_���܋J��lk��0#�K��4@�ə�ᆌA[b���Rt$m�� ���[u��w4�=60�1,���ʱރ�8�l�q�3���^ګ[��m�\#��tem˯����:u;�7g b�,����q�Zᚳ�fi�l���i���`��4�3�sb��z�'e��]���b��(:�y<'�e}$S��N:uSqU�?�xSSx���B��*��o���V���?6*X�5��EnǇ�<�/-N��z�EZ���'�v��s�J���o��Z��f��:$%�קF!/&mM	"6�_���8r"�4S�9v���;��?�W�ޙ�Z�sz���#27ύ�����{�q��ˢmI��z�I�T+�Phoy?r?���8����u'Gfj�MN��uT/�#�f���l��H� �t~��BF&��ɑ-�l�1�"�1�'�f�z$��D�P�p�3J����%��/��5n�C���}����@�M���	�X��{F�*�V�E���mļ=�[/�WL��!��>�6�W�����5ч��Ri,�@�3�]��0��@��`|Y�,����&�|��Y��h2�4.��u���(7�AGz�x�6��O������J4�Ljgq+ �I,�9�����x$0�i���b��a?�gƊhȔZ�!��8qq埙��Y6�siz����.��)��~��=�_y:r�Pe��}s��Sq;ʝſ�����<������sK���5j�!���q��;�ێ=�__����l�PO�Z���ǉ��>l{���D��� ��v� ����;ڸL�E
�Q}:�ݟث�%Q���>i �/���JZb�?#g��3KL�<
��� �fζ���q�K�8Xk�����^^�L��9c���ǹ�~��t���o3��&g��@�baB���D	��}ڟmv��G����5�a�j��͊�����wAnW^u���H�������ޓ9
��6��v#0�^�"0����ͩ���z��ڃ6}��W���oz��޲WbП�����5!9�.�ꙝ��x��Y3�Q����&� LA��Vg��T���]|�r3LC��W|�t���Tr���;�nKx��z�Y�v �f�3�2a5-[���Z��S4����V�^�]tK�*�Z��M�~V�Ƹ���l۠Z����3�:~7\�I"�uwx'U�}S��3�4EM�h�n�*�6�%y%��t{^����s�L�Q��1�-��6��]�1U,���X��T���D��P.iq�-�ڃ�1�$�r�Hk��8�~ח���g���4޿��ޕ�	������m�9D͕Q��R#1��h�ɧL;�/tf(6��χ4�^�IӅ�����n�d���4Z�U�Uc�b2��0�����%��۠Hx�႒[��g*L��&a���93�Gy�iT7�]ݪ�m{��������)k�?M�I�%�슬�����2��[E�������bz�n��(��t(|���K��x �S�`�)�{�ٚ���p��(% �[�Y�Fu��dzgqc�SK.��U8��Aq(J���No�ć��:
�x�?3�ܮ9��1�G����L���Ep�Ψ�d���a�l�՝�����VllKC�\X��h\2�D����$g1S���	���R���Uۈ4Y�g��k���V��x𿎿F�{����q&�=m�G�����sF@�����	�و:l�\ʲ#	<6D��Ps�`��#�����b6�o�t����ʯ=WV	S����L+�[��@�B��tؤ:�'7��d��W}�t�l��v'�#|�R�8�ü�i�NkJn]������kz��q�h�[a^��@�.6EAt_��V����Zq|�\$
�|��G�%<5�=��:�Dy����ᵠ�(�r��Ē���v��4�U���f��aҎ�����CYZ�E�U�x�5�J��P��=?f. �ɞ�s�������q�������
�Z�����>A���}�������mm̖��tW�,��4l ���)�x��u��ڭB���(���kO�B�*9��zy����MY���W�+p���;tQ�} Y������A�s��UޖL[����U($�{�EC�Zx��.u�ܵ~��>��:�����G�N]��L��]��HA�SI�p҃ggy�a!�� ��P���ā0 :���	/gX��5#+��=s�"n�v����rp�o������/wLF�|:%�պ��w\��bHڼX�i�znϳ�����$�*���0�j�wZ���^�Z�]U?J�i������@�%ԁ����mX�r�oąeF�v����7B����e�9���m��@
�x�������M~�u(m��~/�;�a<^h¾@��[\�,�l����h	=u���|&4�������0Nd�b��x%~�����c<��^?�7>����K|�%�Ń�w������ʏYӕ��4��� ���p�ZX�o�n/a-�+�r
�#
��N�Sy��x�־Ш������a�F@?����æg�n��t����88I������Ȥ/d�y �;-G�y�{\o��^$�{���zX���.�I�	k�͝}Kw��`,0��X����6�����l"/e��^i��6)�0���ۄK��R�ё�{;0�d.��Ҵ��2���`Y;&#/���
�B�
��r�_ų(W�Q`�����yS�.��~���D�˙��)]�/�����ċ����@���!,��c��FQ`�%�)g�����a�����4�Z�:9"�$�H�Ơ�v�a�|�\��8C&ޅݞ5���Q
�%��0�^+�"Z����^�'��ݑ_]��&�����.H�5̀.!�_��U�x�m$Ȣ�w��~s�6�]�;��b�N��^����s�~/ɇ�IZ�3ZIu����l*������J,Q��R���4����m�
����?�ӭ�5݅@�g��+?Q��S�1��1g�R(��s0�#��
���!K�o�u&pY_���6n]fk��c�7���T܃k�6�xMhi�z(���ٜ�fA�hDr#�d���^Ձ�2���M���n7�Or����E�]|�cA��P6���R�9j�FQ�;�m�����}���x��_� ��L�F����鐭�Q˻H����m���������a)���z7�Q�)�Ƚb_����B�j�j�e�_���q��_�[�ZYw�8��9"�#S� ��daN�W�h�
�ۜ$M]�PX��$��8 �,99+Mv�B��Liv.���f�F,�_m<B���P��]��FXOKu���ُ'O]��Y�
�:S~���&�:�܂�B�YE�'����tFH�sS/�GH4���4ڪhmEL�H�[CJ�t�X4P;�p������q��{�R�ܙnLG�N�m��rUb�Q�ȍ�eZ��vG	\��D9���	%�J1r�w[�����D׊ǡN2!�Nǹ�����@�T�R���^ِ��y�?[c��#L��� 'NTU��&"̎t���a���q���{����:Jٳ;d6��:�P?/%��AoL�}\�����>��_o.�ZM3rm�dh�ϳT�����*�hQB�m�c�X;����#�x�M��
������+I�ωϯp3/��)R�m�d:��@��-j5�U	�J��%��Ce�1ų���n�V��V$T��d�.�̲1���!Guw!6p�\5	M��⩛Xۺ�h�P��'��$�c�Щ͘���R�\�1\g��|W�<F��bB�V�3Gf?����יAD���խP
H/��*�b��3�w� ��Ћƌ�ZNh�/�7,/�C��o{f[�e�;��AJ��#c)n��R���Cb��e�ʩf��gű)�Ӵ$0݃�*Ij�V���焲S�J��$��7r�?�O��46�i���
��J��}��.!E�RA>�;m�J��1��Gk����L���� n'o��s%6!]h][����"'a�����ޝ2{�x��,5t3Jo����`1�抽Ĺ�+�1G_`Ӣn��L�f��#w��E\t��7[��\b�f�*'��'��[
BZj��>��Ż��T����I�\&�B�T�._ymN���Y}`)���8�2ն��;1�i��:n���Ll�␞�kH��5K�K���4��#)/$eI�^�C�����O^�F%2�?����F<q�nm�u�pC�N��2[<F�3'|<�P[1Q�qp�@�?8(k(SV�)��x��~��Gv������Ou1�0�:]�΅���~�/����	O)
�d&��,p2����d��%Fށ����h�?ւ=���B�� Q&o��(6E�],�
�E����x���Mٷ��K��vꖧ2���*�t�YE�j˶:��� ���(�K#;�� �\v��Ŀ'PC�Ąy.V�ݰ
�t5�~f���/��Y*3-p��KE$�����ҡ{���MW��iI1����I����}U,���4��Z�q���?	i�Ź��o�?k�*���XFKD�)��Y���X�@Tf1�& �WK:���/�u�>�j�-W;-�|�	I�N�G�b�	g��kpg�p�7����6@;B�@M�ו�!�H�
�ɭǚ�^m#�p�|ӻ�oX?D���(��!�����ݜ�\榮i�y{��oR^E�]�6�T�w���t�ΰųئO+1R1x������Dzg��}�w�DĴ��9��2���49�̏� ��ܜ�
΂�����:����<�"�^^	�B{��g��UJՠ#���֞�T��f�%�ľ4�m��v����=I����	��E�`�q�%��o�r�g�Q�#����
�ԉ��a��$/��o?���E� r�K��+�\4��x�l�V2����QnH�Ѫ<A�Y�K�Քw�^�Ĺ�.ҕVV��������8Ǘ�R�d;�����u;�G�S4�6-��Bu����Պ���=�z���K`��E��^%���'u.�b2��LEI�Υ4M���?�����z��S�}�7߮vՐ��Oj��J�]�"�Δ:1���ҵ�&"Mw�����sX���q0O1�V����Ԋ6��7��s����m=����!�#Op�[���	��C��=A�����w�������yj��9;w�8�G_���N"j�o��A�(�����ĺ�T����� ujtia���O�`n��+ �;�%އ����PԽ�TsNOwH�Ye�9�͕��@��Q�U������X�d]"/��:-�oM+�b�Rǜ%C���{�!�]������k��"��
��� Pߨ�����'��}qKUkw���,D�ϳ�F�.u�����]�pH'�K^A's��`Āl]��>�O ����%��$
�ޘ��~������v�rw�tź�I-2��"���$��\-�J�*N��ۻ�1���f�P��&H�n�������l8z���dM�ˠ⯪L�)�v�YaW�O�a&Bå�1����C8�� �:��M�gҠ$��z_�sh�S52�_j霺�~�Pot�+�u�%�қ��8�ٙ4Q�P������3�i0���.�N���FG ��p�T�\)K��v �h�::j�N�->��jM4\1,r*�/�r��P�Ǟ�D"[A��z;��9&���7��j��w�=Y����T�ʲ���z�[R�g���2亹$�\P�O�i��,n��|�K�~A�j�^+�,Z�>b6:S�����v�}�V�s/jY�������K�L*y�z�H+;'ui�%5g(�s���(uFNTD��6��H��F��~d���wL�-��+�"���>}���g@�;�o�x�F��}�My(�o�CE!��#�Ib� �#|kL�G�,�O�x%��U�h�e���hx�]�@�_�7[H�m�t,����i����o:Nw?��R��@���	�;j�	���[ߠ��x�t�7C|@����
�i���TY2p-����5,�/�b{��~S�]a���V��O {oe���rS�Q����ܼ ,�TS������k?��:�N���?�ش�I�	�_[l�U����0V(To��uٌ~u�֔^��K�=�¹�w|����V�duG�#.n�Z�lo�9� �Y��Q�"*����<R�N����'L%����
G*�g0�Y��s��Bi�(��j�r�Ls�R8`��P�NrDؿ �}5e�P[�wԋ��ϔC�z��H5���b��h�j:Rٙt�6@�'�u���A�I����=��V�ҹ\f%P
7���|�#��%���V�A�-��]��/a���7Dx� 8���=.�KD�ǁM*g�3�~�v�
g&��h�ot�SUn�x��u�-Ig���|�I��)F�g@tY|w��q��'�,x�x)ӡ�ԬM��
��G{�3���cD�Q�E�w�]ٓ2�y�����[=����Zy��A��佂)1�5�A����ؖN���L��@e73a�>)x�D�Z��B�V���2�,������̀�>c��Td[�tλ5�����i-S�,��<����R(�l���l2V ut:�������Mbz����?f��<��E�b`��	�ZGB�c@t�em�C��8��}�'"W��:
XID6�;^:� Q�Q!��0[2D$�j��7':T��%��s���(x�Q���ƄAPP_4܍^�}L� �sz�RkL2�P�gM��zoR�D�h�(9�����_�$���`k���E	}r���L�����0���vZ�'u�>��Oヾ,W�7�◊]�͡*�'���B��9�2��+]�IJ��ɲ����6��}��Î�������`)����r:-$?l������F>���*j͞�P�������C��`��YSJ��.����'����891��N> �h�?m���8n�̕�_�U��aI%�7�W�
c7`�2']�l�q�R\	�6�=lP��U�2y���KS/��=�.��~>����s�	�j"�gpud��;�;��џ��t�-�=��+��q�m���C>����껽�4�p'7�m�,�ۥT����(�p��>I$s~j�CN� ��0�j^l��A"g,�3��b;��-�?T[% ��m�S�hu�U���2M�o�G�|��|�fiA}�c?a8�m�~~W�S|� <��k�C2�����+��1!t�C��F�e��֣����-�$�뉋�:��<j�V�! #�����\����ԍsp���at���0A�}Zp�B&�CKby������+�W�cm�VSgCyU��:G��[�'d���bUv��a��}R�k�A��wT�h��ljcʻ�P0�����5�'�p/����E� =AA��� <�f�D�A�e��;^�roi{4��fK�p'	�BX/��)��(0b]~2���P�vm�B��H�Z�bӈ��m��U�Z�m�j^C�vx����5����� ^�ݵ����
Wo���FjuBd /����r.��Z,Dhh�'R��/�;"���r�t0Q����q `$aV�S��t"�j߁���B��W�{�˲�Ϧ�S��uJ�3�&f0Ȯ�r;�x/�i������G=*���`*h�����\jS�!sI��S��Z&�gص�tx���H�V>2�"�!���48�W^~!*�`p�<�*�FC�0��q�]���+��?f�)Z�%m��8~��Y��X4$'�>fH4�L�*;玠��$y����>'�bo�k���IʑUW�t�t�#��b�i�8Z�0��a=��J���C��~2T��x��A����[�Po��;ɬ����$݌��G	UuGϼ���r�TH>�֫��^�=� �Q�lL�#�P*�����
����Z�7�9V���<$+�^����ź���rV���G*�a��}��	��OD�����,,]�:^�����hF��1x� �)`@��`����)bׇc0��"��|��θ�����G#�A;?|x��5~,n:�D7�r�tu-~�J�8���1�9ˇ �J��g�#��M�չ�T�Ȱx�1��"n\?;�S�E�T�A�SUTя2�A�/7� Ȯ?�L�V �*����J���x�N���Z8�y��m����C��u]�T�`19��T'-\׍�G%���SrVw�P�!��dE�T`�H[�?�&idu4ޑ�Vb���� ��l��R�n�T��ՠ��k�͢�_�' ;�!7@jv���k|�������/�q��2���N�f�V�;C�bꈜl#�k��Ç#�k�s՗��,�5��07�
m�ѥ����(��񋿿�|Ǝ��I��9<u���{L8@�m�5��U`�ڠ��V��ay�A�&��M�k-|�ܘ,�n-��,�����7�~J�_�@�6D͈�Aq������;�V1_y�D'�������R�TM;�����N���z�B�*	�)�fZ]|��
��P馣ܸ�����C��x�ݚ�z=���\?$�l�ayC{?Sq��pB��QL�fi��U�3Y�n\��L{EUe�|G�ҏB�Hµ��j8����d'C�љ��y�э������8����1��diB��!����6�'��O���@
���7����O;&-x`#�$���L9��k8S{����n����U&}i�]a�{���� r���q��<H�Tf%b�:��M�IĔ~�2��y&G�.�/�,���R��� ���$��zX���[���bS&�U�R�����9Q�^6o���k��������R��F�_9{���+��Y3P�`���g�-?��j�s7�Ͽ�$�WS�I.yڗ`6�u�m��i��]R���]�><{�𬟨�#�������㙅�j�z�c+�"�uA]=/G���$��F:��=u!�����Ԃ�hzW�z�<�޸��w5�~��	Xs$�+s��g 6ϙ�lys�'�<�D~�^@զ2�UT��C
�<j�z4A>G-�?/S�����ơ�S�zJ��/I�%�gH,u�Q���0B�څ�̐C���tT��R��.XFTŪHD��I\
A��({��K��Y�.F�ϲ'�>���)��^�����F�.���4AK�bO�1P��Nc�*Ú�����]W��]9�>2ɮ�����z��LW�*���hr�9��G��[¢�J�[�b�	��E����$��eO�jB��=�(hCIjI&�T( �b5���	o	�q~�4�s�v�^��Z3Kku@���J�JĕK]MI*��_�k�R�P�(�u��I�#���
S�I�E��=�B:�sc.h=jz�#[��K5�:�h�O�{.���;��Nk��>X��2���Y��Q@&-Z�ڥ[�58+^6Ǘ'��CWW���a��NyuA��$Q��Q�k~�#xۀ^� �&�7x���c�D��\��R��g�B�����Bn��$����jO�i"�O�����:�Dt�sU[2��/�Ӈ��KNm�	؜
�6�y�?���t���Lj{u��g�eg��ޖ� M��$�������_����m��VמFr�W���ҙ$�`kܲ�
/�\瘌�mY�Eiy��݌����B=������T͸gq��@ǘ���չ�U�<�-�������k�Lh}�.;���`��.��@#�0;�<�3!��B|a����Ԃ{�������[�G��Zg1�IZ�������aR���FA⌟ަ:9h�N+�d��I�M�p�&6(�y�	�Z4l=��^�9�5���p�Ԑb�cǕ�q��߫"0'�&2�'�v� �0i6���8�2���}G{����{��t�~FP�G�=�%{�碊~��@��w�����Ѽ�i�PBTne]�q}piey��`󕚐3����(�aJ^�k�/�����v6v��pϨȸ����Ѓq��΄Y#
-�5����Tzk�Y���ec�bV\���C���w)q�£/Œ:1��N����s0�|�&$m�(9�*ZW��R)�$!��Ǧ���]��q��űP\T5��'Sm�̆3�
��<���Ppt�!����M4[����e>��v��J��4jd]}�Ҏ���x|s+#��Iџ�f.�����g&R�|7�;�B�'h���±�eN{�}q�h�#V�<?b��ZXKy`[�<�e5��ڕ��{+;ԉw�[Hu��<���#�VǙ�g��%l7��tu��@�ʱ��aƕA ��������_oBQ��ۭ����GF������D'0p�J��>�eV�:Y�̭�.f'	�d,�q���gjf����X��-�
�AՋXp�>D���p��klup�9�}ӟ<{�: �7��^���3C�q�����f,�i��V�~0�0̜&ɮ�FDazӓ?������$;�@�n#h㘂NN�����ܧ9�g�G�
�$�k.����ֶ���u�M���ޠm���t���j�b���g6�c�߸�{|=��|���d��=���R�u����#βb��۳�U)U��NFѣ6%��#d�`��"�\{��!m�#�7����_Ǹ��/ ��8�A���ƌ�f�G8��#u?@�Ҥ�U�6[��<��v!,xh�m]�8X{����S�ٌS�Cz���%��}�B�B��t�̽P�1}���j.n�ӈ�u��#���ǳ	�}ş�<�[�Y��I�@��ɩ�o�3LLJ=]Rq��},���@Q��X�SB�	�<|ߐe���T��H]���'y�wwbY�����B�3�P�V�+��:� �@���&�#�QژEk]����cb��X��1�cl�JC�_�1Q��S�e��#���f��i�W~-	/	�\Xk����[y��$h�E��&��ܒW�\�����`��z�'l_�����D5�uׅPX�c���CÕ&ؗL�/���3$�Uh����a�3!�>m�
RF��	r"�e^�A�:'�϶�j��8����e��N��D''���n�15�Ϝ�I��׈�[��z;3�oOrW-�J�-�< �n���X�[��M���y
��xPi㯷�]!Fj$�I+�����yEb�z� TAZ7�'Y'	sD="�:��ǥzPU�б�^����.���x Z`�;x#e��B��'F:jP9��:���j
�>bN7^s��I�m�n�����=�ۭb��Ul�XN�U������Ÿ��<Py�iܚ�d% �\��-<���G+$ኡ[x��f�!����P��"�K��U0
6
��GR�`E�� ��~;N"lc�N�	����-���d�`&y#�p�'����P��bfw�Gj�K�� X�N?�I�6w0���tY��AAd�dK�f��@=�vI�և���7�ܭi�௒�1�tO�5�7Y���=��f]]9���^�V�H��GÈP�� j���^� f�tH�NN��*�k�K<�]��3��X;��*J�Z
ݙ���W#U�,:�zX;z;C�h?9�Z���x׏ܦ��Z���P-���sgO9n��-�%��Q����(w�¶V�k/�X(�`��4?��8Q�w���䍪�J��e�}�\�l����0O��aϭҒ��.ҿ?ף�d强Lkv�F�����b��	�i����;�!�Ȩ��Q"� /kgC������bn9.yT��ͯ�=V�E'{J��h��b=�?W�6�)�Ga���X��w���>���L���#���H��v�*������d(@,
e��w��N�)9Q�r�0e��A���^��qMf�G��*�)L��g��s>�MP1�EE��ӻ�#+�Ƒn�A�`�#�i#���9S� X�3��_$��0}?�}�Bu}S�,@@�qs;��~��������&Ѫ��*��ޚ����׼��,���°_}���Ae��5�E��Ɍ?݌�=(	4�g�r��J&��1WɿG���V���r+y�~�&��6��@?�.�麽�Zc��>C10r`a9დD怜�}K��3�D0�+�n�p�<������X"�(&v�[��ҥ��z9�l:�
Xһ�"�.v�<8X��e��R`���;~3��yK�YM�ɾJ^�� W;p���qj at���R^���Ǵ:��NP����gCt�wt��~�x[f?ĆD	�')Nu4��>Qm���*��4Ϫ�mx�I�8���n`�x��`*|�F)�c&�fD]�S\4M?Ih��h���oocU��̣�|e@��#�'�z0߻���;��gp�7=��Q��2���ںk��u}�������#�;6O���n���i=H��Ӈ�\G�c�	n<*�%���.?߹Z$�y��>�� �T0"��t�b�s���*c�V�5F�r䄤iȆ�vfU���+gK�ӟ��%��� v��˖x�ӸW>]i@<��3��"�
b�`��:z�-aRH ���%X���0Ŀ���Z�ɛ_�~P
�\���,pvi|J���ny����tHz㕺�l4<X;R��h�z�$��Z���Pq�$�6;��>S�-VV�K��S�Q�R�KDj���W����p��#�q�,9��3s�Fծ&^���/ ��5|�a�F�V�f������K��3�9��
y³qK���=����o;B׌�w������ɏ�x�Ϣ�~���|�u=\�hu���O�"�}�2.��n��j������_�j�N���eEI�vTC��Q{��M�}�84���
�pg0��e�������:�G��#�l��D\f�E�;�q_�I��ڪ!c�>�j��p�XMM�(��G�2�v��'J�X���Q�	�e.o�9�)��6�� ��7d� �έ��]���J�8�?�%(/�7�֋�������Lx����!�Rf���R���=�KLе��=J��@A�Y�\OL�-��# ��cʧ�G��d	կ���k�bO��,�r�a��T��'�8�#m����Z���(��G��Z�^"�Hh)��"}P�Nq:$�Y��9X��Ծ}D	BZ�x�r>�IA�~%Y�`���w�7b� [&k$�+�qY�����N�N���\���"}`�$!�,��8�
��&���]�AZ�����4�����ED36Ulȫ��˼ƣ�UΏ��	�W�!�y�!!�hj�W��\kxeyC���Ө����r6z�.�2�u�.yW �>N��$B�z[��i��q;O;M�]���i5rhIej\�
����-�xm}���{�^q&�id�4�	�>�!��&�D:5�J��d��~��<QD"�؝�M]�/�J�F\`Fx:�e��g�@�y�l��=��}�<��>�p��(�d(���
pO�rM�ȁ���R�5F���oV�ӱ�]���fҩ��Q�2�������ޗ��I��Mȣ*'C�F9���,�9~-��H�dy�=����e���c����Rhh����xy�e甇�x�ro䃥�TX���;�B�N�G����x
l�Hg�N��~�V��`�CA��ijə#�A��ٴ; ��/>0V�	��o�f��R��f�U F�쎠ȴQ�a^w��$��n^e<��G��ƽT*�gL��@�ŘZ��k��ʧ��^�]�U="�)_�>�O�����-[5�6₮Xn��f���µ��ޡ���!p=�(y�H�[T
�R��ϔ�`��K��'���G�CX�@���Oǔ!?�r4�$*�(�
ˑ�>~Q�$��Y������q:'C_�<]+/����"鯎_��]dOs�TC�$��=�2Q��4!��P1��&L!�;�y	���9<��Qi��j7+�Q�����5�}�w�t���5�� �UCΔS36(t0���𵬥�L)E�T�L	���"��qΐ�y'�=3Z��7�.'I8,��1�5�����uV�5�1b��蠡P��ܺ�ћ�u�u_�LW^�Q���]�c[��`������Q�R��`d(�IeZ�3�jDJ�S����B���%�afz1:�&�,&V�f� �\�Y߽��u�l�%P���$�O�3+���,���
�om<���lS����� Ob̈�D�Y����S����Gª�$���~���1){7��[@���S |�S�$�C{��q�,����q����?�6B�˴��"�>�)x�B���m%.�C��k���:R��~�Y�cG$�o**Њ�hF�p�bT��:YFĒ��c��{W=��( U(�.U9qMx��WZ�"q�}X���2*n.��~��̋9��a��DZ������~A�
�#L`|�:?IHb��\E�H��U��{��(M���Yw����&��_.�p�Q�1�SMۃf+�O/�VNΦ�����|�\� �D�<������|��5��=+���s��*���,����#���o�"���p���TS�O��o?˅r��F"�IW4r/cJ���-�~rϧF(0)@g�;9úx��d�� �Ut%-�f��'z��?4�`�O��da�"�x��i�ãQ��T/w������"���8�u�����^s��t�����~M�C �[��k��H�,�hiL<�����~߳#��MlF�$�H�|�k�	er�:;/ �j� [2��K8��['�+����n2�+�|�I��>"���l�S�!�����+B�IvPuy��I��j���-B��%g��.k��H��r�ݙ��1���G�3RJ#��2F �

qL �w����h����܀
��z�-C]ku��F���� 4��U��]e��Aki�#�8�:�Iq˺��B5h�*�|[�F'���ޞ-~K��@�M�=�:�9�ҵ�/��Ր�kc���.�� ��Y�&U�B��O�	�)͎���>�a��siue�O�˖�^'��H�&�A�H�I}���)��ϫ����m D}.�a��T������i��a�vR&#��o�y��i�pv����h���kIw�(k��eS^ǹ���E�'^�)u��Tx�\�z~b�5G�+X7�!�CP@�7=\M���?�j0c`e+�V%}�e�c>�5��}B�������f�~�9̢Ώ�7(�E%_&3�/�5�yW��8��>T69�ҍA2xi�ַ�)'%=X:�6ZT�|�G�l�S�KF8.����h)�N��	�-����r��dWS���SD�T�|H�0g2f=��,��FЧZ�q������Q�	֖t�������]����9�Jx}Q�J= @�,ܪ�j,uí�.:%�lC@SãGX�]1Qc�"�>�U��@�Fb�~U�̚�>v(��ٕL���H�z���_m��t�,����n֪���C��������bq�Ř�<�
�Q�����$P�swpިER��7���_Z�!% ���X�`N_�����p5"֭i�,Kn�W���BP�y��i��~l�"�T�ﴷ�$� �'B���N�	�# �.ES]�eW���d�2�I�1�s�=�5lƗB�M�r.{�����$���yU�̩5���m\����I+�=_lF{x$kP�^E��E����Q�>7vSp�	cd�~�W!1�s\�r�>��<`? � ��>�"?y)vۡR<�k|�"S�mB��J����eݪ�1l������1z}��t��\�Wk˚H��O#��sz�%���&���%:N��Ta�u`GP���Xj�t��������z����lw�Ä����>�����ٸ�11}\OG?Ӥ7�g�lP]��EE�p��}�5��+�s�f"��w����8�t��]��}8��v�W��� �gmg$�<�}�g]�tL����A~8�'՜�X�I9�IzG"�@�T��Mrݍ퐛�M���6��+�gU��W�/2k����`����i�}|ȝdB%6�UKe+rgB`i�,��
�]
kIJ�������炃V����U����`l➌�h�v�b��OɆ %��܌����7�,_`�4���$���mg��V�Pv��_X���Q�L~����Y>�oo �k�iZ�)��^
�^l�P2)�W��҄H�<Ʉ��*�ZF;���isK��J������L+V�'�}��˨O0M�jV��t�}9�����t��P##�|���#D�n���E�pu��/QB�7ۺn���^,���6)�	�(��cy�S,kE�Tޗ�R�	❖5(�j��8Ĳ��w�Ҵ� �8���7�snEq��Oj����ޏqN��u�K��LdMl1%	�	r2�����t�lc����$�I0T�e��K��l��(��Z���0���t��|b�֕A��_(�˻�ې�����
7������b�拮H�
?�Z�Z���
�s�Be	+Y�_�j4��X�g�������da��1���x��ht+��x�y�Y���%J׻Ca�,%�'Qk.B$aqX���vLVw$/*$4 �NCē��>� ʵ�Y�)ϙ�״6l��S��v@Y�r�v�[z+D��eb�m�����4&E.�������0�
[؅�Mc��yi�y�H����?֞<��hd6���s}�_�YQ� a���O��4�G-.�dۇև�C;�*��ǝ����7�l���!�\&��	���.և]˜��N�+��Ӓ��&��k�ci��$<�A�pA+|l�!�4�;?�J-�hL�h�e��B����[����%����_�*|]� J��a2GwPCzZLn�0��ݥ���	�K��V��eh��syΥ3X&�Zs9�f$޴�r3)��%���Pjk��DT�������K�_Ԙ�1l��S�N�g�D|C(>�`�*(>�K�#0;e��s�����Z�w�׳DH1���U��ȃV��rL��0���4}�tܿة�Q��+��I�e��Q�����Ԣ3�e05��u=K!O2©<HT�|�^,)֕�PR��[��+��h�4�:�vU�&@,��\]FO�i5�x�3���9�v�p�hsz�=��nY6&���z��� �S ��{�:����B�B�ۊ!Rt���6�ǂ�<% ����v���������e���4v���Gg
����^��v�m��V6�P<��[ķY�h�H���
�#�C�L�d1�n�w���CS#h��(��<\�h�=-5Vg���8ˉ������$<[Mr�$�Y�����;��ɑk�b(��<�X�T����6���ϟ�1n���vW��f���F�|����a�� s� �(Ņɩ�Tb�_׍���,E2-*r�xș������-nc\.wh�mצ������>�'	�����Ĳw؀�r2_���nA�bp��+��xP���X?r��F��O������e�J8�|T)������vpa�v�+d&F�ob\�5���8v�\�cq�+>C�^c�e�%Y�	��I�ȡ�84��>}�l�Gi"y��D)Ǐ�5
6vV�:�
C� TX�w����mjH�	T�9U�5��Æ�j����*����)S�����J��,�#ݸ����uWeE0:�IˋӀ$=$F�b���noGXc)���gb�W�2s�T0oY�;�ح��>59�z�g:������@g��Z�?/��:�8���\�|B=p����!�~�:<YYjӘ�b|�{��L�5����k��'s�d��{3�$*��{��#�f��f=	 ��,4��zw�0���'�'���5?tIV)#p-D��й�x�B5$����>`]E�*�m(��r6kG���Ǒ�����yCE�KsC�o�'l~�Ш�u�p�G�;��?��ȥ��ض�lĝP�z& �YH<H����׬�?� ։xt|�˻x�R?=�?�<�H�e	-"1���A��&-��B�YṰ�w!Osm�g��N�h�Y"��4�g�� :6�~��:�(*K��w��F�I�r��SPEA<����Z���A�d;w������	K�8��VT�0��_%gM�Ϩ8cCS��٥�Wѥ���C�y�O�WV��q�Se��c"��
�p$�Hmţ�U�Sc|� ��F�.����Y�뤮f$�}��HrIoT���|�O��ͅ��_X�6���b�ޮ���"m��{�MrZ��`���"u�2
9��X>�"$"�q��F$iV|�,sn�5>��E�"�n������X��f��d蓒�;/�^��z��B���1��{Aj�=�t����n���M� ^В�� �����i05G�%'�N��~2�4O�ލe�v�~wJƕ�O_x����$ �7�1p��6m@� ]$h:��$��8�C;$?SC"�j��)Z��x9���2�3����|�]�6���Y6�� ���w�����܂o>h�~.��F�)AY[��%�o�Ww/��)��)(�P�>Ç�+,f/ H;�WmXꔗ������
�?�K�����(�����T�բ��-����fd�)[�Αu��6(�P�V+R�'� �>.��Y��Q�m{k,A��i�B���i;�S�(&��j�9��1MZ��2� 0{W	mh��iD�C�!ﵙ�R��&�nv>m��gr�<���� �"�<����S�[�&��rKV�?��2��	����0��}E�H��5�W��=g��/����DP95����w�C�G�
B���6Iq({}юċ�oZ��}n~��؁ݕ$�>icJ�ַ��!q5j80UQ�p^�8u��W��n*#�<},��h#]��S? 1�O�v�I� ��֖����A
�T�d����h=����Q)�\{u���-Gx�;��켕w&	���U��~�_4g���@��b��AD<��2��y��ྖ0��3	.�~,��zV7J:E��ǩ9�0̔���v&ЄO��l&�b����*�%+`,�����m]��`�u���-l��x��-a/�����&�����9F@��luSF��y,�8%^�	�IvPMw��B��V�E3���,"G���\� �|JH��%��k1�p��b{��)�nۊ^ҀH�t�}�t��Õā��t'�dF!M��z���{�s��tm.�%���w�IY��Ɲ��|Q;��w��9���.��=�O1�1 LD~��l�}jk���s�gR�Y�H�	�J����o�r��$��]���r�4^m�f jFm� �����/�kaxR�/ܛ�ZJV��-5Lue�J*���_�,�&�zv!��<������ ��x�!��n��� ~��d������mk*����)��,��j�J�i�^n�oVd��
�)���eD�2���gT4a�S�Ÿ�����|a@~�E�����(��s�Tp:�n3���������>���`�vվlh��P�V.��S0Du@[�m�^��o����e��ݎ!�H���~��D�oV�IW+��,��T�IQa�ء�?�v�?4�Vx�i��[�E�����[i�6��%f�՜~g�,�1�����Ω�I���6�]ڦ�/�r�3�ei Z Lt�4�+�>��^4��q��|W�a$��N�dO�m`�5cc
%�ު#)T#
��W��aW�*u����c�X$SD�;D�����-����vE��ъ��ZH=����!l���j{�g�^l��4e��=EF�ݗ(@��8�Γ/C��T��x�
�ˎF�#��G(УQ���旺���kM�7��"�� f�Ӷu��ah@�ہy>��(ruh��-R���.���KeK�.�ՊMcE+�ɣ�+5L=/:�'��ָj����)�q�*%4�7T�7.I
u���ײh����]ܠ�~s�HǺ�pb�]z���P�y��=@�I��(I��\�H��vK;�1+�����������
�]�w�2}���o�S���:w���g_%[�/�I<�C�Y����}k�ˈ��;S��[���2��^���=�i�:*L�?H$-��s,�0A�9 �U��A��J0"�r��۸����rVl[�zGo����J�$��)��V���)���a)�ك���"��Ƴ
`��q[����G:{�+��jg>N�w�V��ޱ�5'�{D򘀚k��H���j�Ww#:h*O�-���q]��˃Y�t.��JAeǾ�&rdi��0)����	����@?�����U����&;a2n��p@���0����+�7��-Æu��J.2�����@v����$��t��<�z�U����}J��FL�.��6?�+IZ\�+��`�;�,8�ģGS�K��TJw������r˦zE���uԤ��GD��$@��A�Qw���(��'D�,�E1)<	0�\� :AD����9�����}�%������'J���Hc��'�WS{�cq�k�_��"��yQ�T�{��"MZ��8
���Q���FF�|J�Gcc��̷�&�)W1^�5(��i���#��A��Զ?7L
�Ͼ-�	0�1��<�z��U7O��NY����3�M�/�P�_��G����;]����n��hϥ>%��'���i��Ф�(00���nf֢o�\��FH{�<�Y�yd���O��j��,ʳ�7x(�<��I�Z��~���:\�5�{�yÛH��o��cZs~��Ff�3g4�?�3o�	����߲�b1��<�XS���Pڪ��S�ף��,�a6����	��]�o����&D<7�r1# �A��j"�����&�U_>�F�3p�zMD[�?l���άa��u>x�R�N�8T<�����:E��_$�ۖv���J��SI���XU�������+����x��`.��Xf�#�����j?Uq��|������)��y����|F�㾇G��%�R���ߙ����q�UFI�_5$����D���P!�hvFq��D[t��?>D��_|Y�(���i��&�W��:�$���$����zx4�q>v�C���,OĀ|P��::�?�q��`�~1h��|[g�b���=>	x.O1�*D>C���DQ�.
"3T�T��l�oZ�v��4���d�	=���.�����&_ąF_���	�\pI�����6���ͽL��tG��KpH������C�7R~c��~;�K�si$\JE���R�Td�6�"�s�W���Gg�U�t��K"X��{[�Sr�-����G�4n�I�	NJj����hC�gqu���$2��C�Eť$k�A�DR����z>�θ_�j)�L����ǩ��أ[�}v�f�9Bt��T8ٷn*D�2�/��m��Uz��%7JV��`b�ty��^��kUtt�q�o� S��9!G����Z>��ۜ����ս�I�����lI���6�co��BR8�8�g�������ǏK4[y� �R�2�k	h��Ba��w�
H
�f���m��^���pmM����Z1'P���L��e�M�3B�MY,�{Ŧ�)yc�P�5��\Љ�n+�����p�D�/���/��>���|D�k�'|� /�a �V�/^���7Ck���)%N��G%3ӽ���{=�����C���D��Ũ��R��� ���`��m��yћ��5�s:TC	o�Y6Z���P�:Hc���7E |�(�zt�� 缂d�[�9�I����?������o�oA�
�����g� ���N#ZD�.�9m�FgRV�7���ʴ�T�g���3I`Su��|=#d+��>%C���)���' ����HH��Kdj�T�W����[��(߉r��:��"c���ҿ�U�1$(O�a�˃�G���n���A���'V魮=Gy`�����SB�a���<�]���+����K|�U?iᄪ��.��M�[<�y�w4-�=A��h��AΜ<��mV#�d���["��v��B��<�\9J�Qw�B�B�/\�͚�@��SNn�2^����j��B��w��HЄ{�uq��i�G�߼�,킯V�*=�KQ�fg"r��1�#w3�j�d�<-]׵2��5��/|�%���l��S��s\�����5���q�FI�V۝�OW���-�C�-Q��nWp���LH)5*�9�dQ�i8���'@r�&I�>{W�Y8f��J�����{��ܼ�-vU����AN:R�-Y?y�Փ��N�וK�N��uz�����%� �V6�mȫ:bG�PO1��5p�ߗ;̪�׀o�j����h_h�\�-��O��
��F`m��{f�������E�}�(ݢ�5
T�"�>��)�݂iD'L�]��9tO	�� i���z��ϙ�x�����wK=��K�DϹ[?���w8c��ި���� �z�Á-���K�3��
�|����Ȗl����X~�L� ɢm�ܯ�qAp�I=OX� =2,�jd~�+��{�K�no�����i�%[l������˝�Nє��na϶`�1���S5Q�L6��+[X�v��%�[В���0����HM�o�s�3��i<c� n!����׉(`��[�~����|����M�N1g���RY�R⊡>�s#h2�$(�'����f\�zfu��9��ݚ}��58�8�>"�����́��x��W���y��PLÝٙ�BKРaNШ�#/���q�����:�`h���g(�Ե�	�e֥)vc��@0z�2E$	�{��x#�<��y�N��0_%�f��Bd���@���P�Մ�S"��"�1/X��N5~L���X*�*�]�'��>#+��Ba����e�;��m���N���k$T��	V��F�b�;�β<�]@����AwN
�����Q��2�#eu�e4+�0]������訁 � -NΠ��ŀz���EY�=��t�b!adu���T���}�C�1���΅K��d�PH�����3Oá?5l�2!_����l����kA��Lp���F�do�D��n9��>6$�8���1m�m}����&�\�d����@�V����>ʃL�tt�*��g�������Y��Mr�"������^���@�M=����;��n��Z��J0�!U�ꇯ.g¦-Q�2�m5:U�(�U*L$@Y�[v�վ�|6̋�X��V(�
���P��;�q���[��ݐy�%Lt�9�#�u�����5Xm��W2�c�����I�o�L��*���о��͔@2��R����9lWKc6إX��<o�]cLu�2� i�+�˩l�4��/5w��[����x�""���336T�8��7מ�8�Jx!Ϻ���̓ԨX�Zꊔ$LOc��f�#=�(wX#�~Q�Yz��+U���1Y�;512�3��G��6 T�2��ג��$�k��E�/�,:�1����7�)|�۴�KMz�#ݭ@W��3*���%A����䀤ޅ�v (*�D�qVJ�Y70�O��|3�w���,��C�q)���ϐl��$�c�9�����a/�r���P�Us�}Fؒ伃�}��݃(��ل�}NJ�g�%��}H���*��=:e"�CH�x�KeI|����皿�H���h,��WL���*x|7��9?��a�熡�l;�у��m�"������c$�.���E��ɒ�R�M��h^�'�����yݿ ��4b���g��l����.s�~�g�ݴȴO=B`����i� ��Hc�g롍"̎˟�3I��`�"��Fqm�1 �b�#�(��`�����\�jfH�� �}�-�%]�`�;�~eRr~\벟���2�C<RMLG�{����QN}����n�Q�y������Y���P1Q��s-�C�tޞ�r� 5�r�$�е������z^��6
)�WF?#tA��"��� ,e�"��k����]�HA@�9e���8�i�L�R*�Z���e�SQ|�AX��U[ +��L*�z��t���d�]9٣1uz, �Hӵ�8L��`~k�4��.�]��${��f.�"��yl|�	�I�bhȴ,�0D��q�Wd��h�$4d�}�u":-!�Q��֙�>Y���x���ZP�hl\�l!L��K�-���Gi;�8�Q\��5#S���EP5]�rE�P���*�k^��E
-��$��`?��� ��ٸ8TMlӯv�b����7�L�"ʳI���>��T3fm��ҭ��V��ߡ.��M�JUa��86i�'wǿ4�4B`�a{��' �PfL�ec7�]%��m"��ϙ E��z$�~=�%Zm$�+ڰx��[�~�r�ό����P��;md���.i�!�1������w}�V�v2�`�M2I�/s17Io�h2ܵ�:�#�}�����y�}�fS�tB:
�O�m����c>1��m���=|���^��E���]�$��[��L�^�ۏi�	7{�o�)�I`-���B%𤌺F��ՙ%�Ж��k=7�hh��?���h̃�)�gO�q������{�#��+�����щT�?0��I�˴�#�����%^j�=��Ά�g<�v�9��zM�)��>�W5�G^����g��-��p=�
��V��Q����=`�L�+�P�e�b���4+ɧ8�����{��]O(�u��2ƅIAД���k���T��G��bO���c��{��C�;L�%�,S�H
������b�6_-7��"�G(1�pV��[���-ӏ��{<F����)6;^Z�F[3�v�ײLY��1���-��܁z��ôܹEa�~��\��!�H�P�� �#O�4�kD�n����X�۔��T�a.������otŚ�)y*J�ᙽ�/�,����L�[?H3@[_�- ��j�A�A�����I3P�/�8�W���s/��#���78l�,��*܄Ƌ���
�ye�/i�F@p�'E=(��~��ޥ�����U��9�S�<�$�^��Ǜ�j�͘y�H4�Tᴮ�k�A����c�`ӡ�A^�_8��V06_����k� =��}�#2ߊ�;���ߠ�@��-�n��edv4MV�A:N^���I��XE>��^f�E��F��� ��}�W�|�������"�V��-��<?qS=�	�YaW�{FJ���*SP�$�I�Z�o����43 �Ѧ�R�H@�r��2��� �eF��q�&�_���6�-�W4J^�ޅ��O5��(QIY������8����k�qhA���(N<3U�G|���%�6�S��#����� �0h쥣���Fԝ �юLX��o*/���A�_<�Yz�I�q`�G �Q�`���)Nn?"��iO$=�xT�������9����VK�02�����$�p�5�����D1�'K�?���}��yU�񏃟h)���
��o!�3u7�Є`-u<���!��b]QI8����+d�w�$'Oteu�W#m�:�xVMe�&�Cx��U�tjD%�C�8`���;�c|2�����n�ne�}v�1fm_u�#��$���$�K��n#��0v���O�L��W�j�ו�	LX�_/B8|	��{��w=�����ݒ�X���[`!��9]��Ƞ7Kt��b�,�.hg
�[�$.O�h�Cr�s��}��Q��J��r����<lY�Z�G|;�_o����h�b�\r����X`��c2˓E�����J�`¶ѹ�����{��ӭ�eQ���A((��<��m��z�����,���0��A�A�ߟ��j<����C�]��W�\�������Z�[[������8�����j��}bc$q}�uM��\����=�f�m� �������p�{�0[L���!���}~��ھ�,�<�,5O�X��d����̾��J�����d�.�a�0=���s�uz�����NI=w���%�#�90��?O�RN��U��Ub�2���ʦ�:/�`V7����]�%SIR>#.�K���ԙ]2CB���ެ��S�5�? �j��P�[��B�4���nR�0<��/b�&�������3=���t��Ȏ
u�D���j�`�eD�!�q�>����$~�QG�VcR6��Bd!|3L82�n���L��0W0�8������T�N�ʿ0����3�*{������G��Lt�ˢ����iĿE�T,P�ڬ3 ʹX�$�l1��AM��6h��EȔ,��c%�D��ͣ2�C�����φ��_)���)yf����&��j������� ����\�cK\�1�0�@��
���0f$�m�x��F%�V'?k	G�s<{ -���fG� `2>-Ry��VM��/�yE�n��vk3��E͜�CG�-��`^�:�$d��$t�)J������}�I�֢ěL��4��읫�cm�M0�_L�l���|�3����d�RTB��_����_>||��~vv�[CX+�T�F|��E�\��ȷ��4U��X	�8����|�3�b��r���i�3�/��w(}^���73�}{GKK 7���g/虒J�ʣ�����h��5��?
�ym1NV*�ٲ�Rw\6�`�Q�G���S��J��(a˶�gÜ`6��|�`[��H�A"�Xې�L{��mp��x�v��ek�)�J�Ő�pZA�+D
�4iK��umx�`П��kb����T%� ���p%v�@��{�dS��t�Þ�
�:�Ob�m�� D�ׇ��S���ć�hG�5W?���� ķ~o��rɲ�Eb4~K�dR&Pc�iT�Pp^��;WH�F�G���\�=Ckئt�Hv������CJ�2F�rGK�X�Ъ�ձ�G����`�Z���:�	�y�� W+%]���u��U[�A�5C����U��e����b�F�������2vȍ��z�]�L���=+��J�]��+����Y�r�%�w��<���ה
�L� ���ub���a��u�y$��q�=���F2V[�1⿒���@L�Z;�-�ᒀ"����C�(��rL�`�"�Ux�ڟ��E�Y��r��p~��m�r*��������I�g�Ԧ���jQ��f���$���Щ�=��0=��\�D�xt"�T��m�LJun�l��Mn
`+V{��{jQ�oT�/�OO]��J�)�j	-"uwr ˢ�]Bl#�u(i����'tnO�J�u�������X�~�� �M��)�5��h���XP���dm�_
�]t������ڝ�B�LXL��w��E���s���#P.=���ހ��l�����侇�Ь�����*= �o���X?�v��q7��P�� �ƚfx[Ȣ\��A0��� w�)�����M��^
�D�F��m*��x�x�K�7+��&=�/�$����t��Ɛ�s�}��^gr�Z)�5ք�� &��ɬ��y�Џ2���Z�$�S�����>p���dw�}b��݋U�q��,�� �t4��sW�fE�ऺ!�|��һ�O���NyzT �'fj
�X\S�;[V7��&��^��X��L̵a��r���h}0��hr[��3q0
���k!��{����ix>!n�'��p[���l�e-�;k�l�"j�oQ.�-)3�/�u_�oHE:d�~����t��
O�_UwR���?о��@��ޭ�mLDXs��uЭ�=	��3;z�m}��<1���ϛ�Z���	��dS&u�у1\`�)�I'}��F�8��݌��U�0���nN\9W� zT�^W���t0tV&1u[ã@��x�N��ǂ=6�a���_��R��I_���,�qۄ�Ն%�4�@K\ t������&[�a�h��<�v���8u�(�2{����Oݙͥ�G����&����bc��� ^��CΈ�!i�Ne���v�,��*3Pn^�ۋ8r���nm� ���
rZuM�(Ր�v�f����7�h�D�f/G� |�<+������%��*asp!s�d�ޙe�̐�7������xu��Ha���騬G�\"d����(�Pe�0l���J������6?�L��S~"#sɸ9:���o��V��h�����B�r�o�ْ���r�`�e���4��iL1~ʑ��B���k���N�t(ж�(+/6_�� ����(&��-$3?����yȊ�8/�"Î$��*��#��������9�UE]A��[?�8�	����WLL���]miwS����0/DU><,�Vl��/	��v�Fց�n���~�LSJaZ�)�����GS��K��ɟk�;����{{IxVy�@���{~������Z�M�줅��ED���fu�u�E�d	�t�7������ܪ9kHޑ*�YӀ�vb�{l5n`���Ka7Vn&��2fL�&JŞ���/盓�� Zzz�{SE˞&�aAI��E����q�^�h��~1lk�4�N��]�v�iUf���F�{]S��3��bB�?-W���U�ڤ)�%Y�����A���Z����J���S}^�X_�;��3��wx�u�k�4���_d�9&�$�OC��������\t��1������5n	Ժi���մ-C $z>��08��Sh��_���5Gy�Q�ܫD���B�z^PtB�~j��P`a�37��uѾю/�*��ۡh�oh��I�\�7?]6��L�W>�tgޙ�i �M���<3��bH�Ӎ�� <M�� �)��oq�k6�O׎�XoW�pj�g?H�˯ԉxM�Ŧg����Tہ}A"_Wx��]S@���yt��-���q�؞$���n��;'Ot���\�y���"�9R��L1W>����T���]���ʇ��X�j�y��2ϧ.v[-+&��8=���Qy���g���0�7,`���j�*UfY�H��,���R-�4z&�K�F�o����y�{S�d�P�$�3x�h�,��� �x����o��Rx��r�8��_��+�h>���њ�A��#����u�T����⽡�A|]�^��1��Qo�I�D�p��o΍�.���.��L�=�K�s��R���.*>������7�:�굘��iɤw$�в�7t�u�����Y-��N �rH�p��:�!gɞ�Hi&���;5N8l{%�'�ದ����۩�M��� �M����k[)_���������Jm�/@�t��L5���D��p<���'Q�\���C|�L
��鱲@K��I6�͹�2�Z9e���q+�sߎ�
�R�Pi&Yq�ZA���b�s�����e��������;�3S��OVQϯ���9�j�a�j���"�L,X�R{�-<<	.��IW���nK[� �M,��i�R?&���M��#��o��Ezf����#�(�(�[�Af����0���6�o��]:Ɖ�惰��,�V=��r�vgS�|�J(SJОh�Ғ�&��U�D�Ҩ_���8��˪6��̆�ׯ\kv	c���o����uC���)l����4J
T-��Lه糏���v\���0�P?�:/p�=0���HVR!�y}��D���}�0���i2��4@�a��Q�ز�t`�Jibsk3�-b������uAU���V���@�WGp��c��'��Z�`T�t���݄JZ�ω{/���ŮZ���/���o��1 }�Є���x� u_{{�{��B�c�.쫬�k��	s�ٸ&OPZ��-
$W^�m�������W�H�J���=T7��~v�x�L]Ii��"o�
hC�#�\
�.�>'3g��H�W��ń
n3�̸s)G+(ӧ�ăo��`�,��/p�$�g�j�=�f+:�(~<�,[�Q�������+�����<G��+d�7��;
s'��(��(�CͶ�9�Xէ-���k�O=Բ�>�۔B����D�O.�xF��}��7}�j�@'G=���	܎↣X�cgώ���#5gI�jN�[�u�|� �Q���J2	ԝ=���p����ק7"R�/]�#��Lp�T��(����%�,��2پ����p��;�ߞ�0�6�7�!����k�#܂� 7�o�N�AYZ:n��v:���pWj�e���,[+�"WXgھ��`� &�`5ϱM~�M9�*o)�w�T,,�5$�y�&u6�`��M�gn��:mnd���o�#<X����_��i	l�{%�T���&9sl4Ձ�T	 ����]ص]Tͮ��
��0~�}	��z�T�@Ab�=طc�cN��D���F�N1�(���bK� U�S|`e"���#++��o��w����"����iᔭV>�b��T.3>�3��&�!h2��4X�ů����c�����V��f^���`����,R�Ҩ��� �� ��*�ɟvP�6�����
Q�.����T2ĩ��?����q��7�0�;�s�Sxw*�u�1�q����|)�
�G,f� #Zb���١�4���ͥ�L��/�N��e�����[���<�:���;��_=��Cu�0����$:y�+�%k���G4?��Y�d�ɋ3z���V$�$-.<�kNt��l����[O���]�Kƌ�������g/�.D` q�r�̭�5��6��N�{}5fD>l+İZ��f���ج��"AM)2����_�R�A�ik�s|�T��we�A����E��~�/�e���e�}[b���N��=�H$Q��N��$I�׌�|˵�V��m}Sw��z��(�2����' ~Y�BPӰ6�8�%7�N�-�f�UR��L��YH�UB���%�x����v�N�딑��J�L]�5@��%ƣm )vt��2���8k�ޒ=�������������[�х������uc�&5�A(VE0�^����H�z��"�ֆjW��#��3�:��E+O�A�T��ZRgU<��OH6[�j1�SW�g��o��V�pu���Ƀ/V�����Ѽa��,�N�H2)P'Ł�$�4��P2���:q�B�)�����پ�|��g��^U�Ti�I��u(���H��[�z�D ��\Ĕ'�4X��r��Eχʼv� �m�ln<aچ��U��8�]F/I�Q����f5NZ�U��T���t�}��.�12z֮���4�/o�\�/n�xN����Jɕ­�����ZΣ�����:7�/ܼ��q��V�HCs`Ԫ4�����Ҟ�M���K�!V�|�<����WSK4�sxx.D�B!��C��//�s�:�w��㨣1?
�����٦�1�eH��QjV���6bT�'��Sk*�]��H`j��bϤ��_�%�]�����z���Wx����د�\��X�PH�s��"
���1�p	~��#⾊� �9��W��i'���\3�kU�CK��j�f�g9+���H�ϔΓI��{�$F�4���9�f��E'���	�k.���]���|���t3Q;��Wv?���������_3A�� j�wi<��>y���ż�4ք@<�6�Ʌ���Q.o����W҂- �<��h�bZڧ�(f��3���I�+2ɣ�!�F��@�+����l��w��&���@9d�#Q�٣�n �fǃg���x����b�Ϸ��&[�6U�>�YCH����J� 1�i�5��"Tp &��}M���!0�2$c+��%�W[� �%7�.��us��
ξ�m�W�Z?zLroq�N�C6���]f�6�x�T�Ѭ�bC=�^_~c�x�]�)ogb��P�F��V�ƺ�l�g��ԊB�B0ԜD�X{
��!�D��G��1,����a�V	(b�l��N>�B{U��v#�������i� ƫ���i?�Yf4��E��A�o��󌓃lQ�3�^TP�_��G����H�eQ���A��T�v��P���� �p�T/��
���;�S64r,?�>wA0���Z��%m�\̉î�>{�p�vi`�2]xV1�@��J{S�.]�`�}�����)G5�,y�� �iԷ
��!Sv�i��s���FH�:�/!���8�|��S�=��0��݉�`����N�g-$�7/��ϵn�G���kb�j�0����X�Q�;Gp��I�o�	�q
<{WJALY�o��#׷�ඁo��	�Y��\!֒����v8���M۱�HK��S�i���Ki^Ò6�Q���ǻ��eu\4{��.60%m��u�!�tW�7��ʎ[gq<$�l-~7"�*�ߢ��Y��X瑽�,]a��v�&�|U�|��u�.n����!t�v�5.'c��vPӇ��Kػ3r�r����R��P�O���xY��e��P�ؕ B�,��A��d��oP	���zG�Ĺ���!����d�Zc�F8���U�!����o�(�Azu�b�K��F����Di�<��3x�9��n��C@Ͽ��.|̐��8�o!��Dy���[��pu�)8�YT�?�+���	1���9����L��u��$�./g٧5��$*���P���APo<�P��s�?�'D=��!ڠF*Q�Z8*�hG �:�\K�ǑdE1�,u�%/�f��#'�-��q����<cFL��H�I���J�͚9�Q��4��NR�m?��$E����	�Ԓ��~RW�M��E�?Jo�H��!��4����W�CM]]��c)18�_{�-��X�p$EN,X6��Ȁ"�l���Eg��3s����u�,�`0*o@��g$�l�h���9�����t&���"���{�%���`����`�$, xs��c�(Ř�{��${�e,sd����_g:����#��^���?�Bݯ�� U���3N�o�b=��w'��YN\��3�Ǩ�:,C%���GU�x�s�z�LE*���G>h���伝|Z��u��7XBFPpң�.(��H���-q����Sc����Y~b!ߢ������mKa��{L����vO )�C@��+�6��ܱ�]�/�ˢw���V���+j=Md�+��Mg����@�Y������Ī{�y�3���@��L'%_��z2�RD�ޙ��-��(R.�*|��ڼ�����v�JF7�
7V�>*��r*���-lh�C��u�do��]9U�Jm��IH� �iIB�J�������������M�]Ɠ{�+`I��6ʻ�+_����h)u�PK$����G(�;�m�t*$�Z�������^�pf�К h�/����h��l�����Ǉ�񧐛��H�W�M:�.z
*��Ʉu*��t�&x%�ȕ��l ��m��`TÈ�����'񉎉�q�ipyU�Kj�Q��[�;r��,��������G����������J��d&=MM<�T�Z�y[�I����d�5+y }U�e��[������2
lxB�B�G}/��d����T�P֩��|t���V5��Ҫ��<˹���T�sQ�@n��m�DKt@��vl3�f��	Ϝv�l�������+J~^A,4$��R��d��1�0�>�o��G� \,fVS�M��2=m�Q�*�P"���Zn�����7�������w��F�]q،{���%ި�Ba�r���d@z�@镸=M���n�U]̫�~��&�	o�Y#��].���
��:�_��]����pK,z���q�T0��Q��S���gL��ݏ�xת��U�)� gTdS�#9>Qj�����h������� ڄ�a�ε�����;]��{q[1A�g9��������_2�
HȀ���k`�
_��`}��`ֆb��s�*���ɓ�@�����q�Uo�g��oÖ[a�Q�A6���F{���XȎ�)XƂ)�>ѫT��i���{,�P��@G�Nf�|
<h���-�
'�d�k���=i�wSv.�a��۱!!8�a�DL��pQ�]����{z ����v���u3�٠+��#;��=�nn|���޶��q��
8yYP<�M��J	��t�f���Fع[t���0�������xVvk�^sA^�ӑa+[~�(������H�3��{Q��,��j��d��n,c`�� /��Zӭ���@��<�+��Imz{�?�vN>��@Q�n$5�Yzho�d��֥0��:���o��O:����	����-R�CX�4���e/dTٻ5�چ���ݢ����8'��6�k3�c�����%�|
�)�����-�݅�f}�"�MH�#�m���[���$�u
@�F�k�p]ye�M���Yݕ#�[-��&��G��%��1�J�{��6��+YG"��\+��3�v�[)�r>@������ Y���o��턂:xW��d8s+�|����4|������T�$�ľ%��|��mC& � D�㓓OF��u��P��� ?��q��>gE���x��s$k`��rO��g���^��z�&͗n)ed:2'�_D��G�2)�"�~߇� "mO�S@��Qo$�=�!_]�,��6��K^?�)�po��x�R�?Yy��2i~A��@p��� ����n�	m.�(���Ȧ|p�a=�e*�?ZC�1zcH�լw���㥌�]-EZC+{�U���h}�#�
�/�i�?/wZ�]�aަ�G|_��p�����s��X M��ֶZ#x�}����e�
�{
�X� �SW@��}I��Z��]�"�lg���·�@��8�l��N�C�<>�	���Y��_<���'�3!uar]L�am�űo�M�7�_�13KKʐg.%���&H���v� ��+33	�S������j̶���2r�|�o���)h�:]k��1�-����
M�HS�i�������N�QL���s�R�ട���9t�繿�*�u:Q}�G�B�	�z\���#嗻��+�:�ݰ�os��?z��m
��k'Yʳ�b9��4����%����u[D|������c�����S����މ��e�7��?�YzG�	e
D/k��IF��ީW�ш}<���:�De��%�lĕ6p��<��D~1�)[`:n�s^�Ӓm��x�cv��[�7*$6��� k��ѐ�h�S5�0�נ�֐x��^���F�z����Sw����s��σFڑ��E��x�>?cC��VSo�%�	X!���Nu��ӆ��+N��Ė��b{A��a�4K�`T�g��}�}]�����/\�+J'+�s|u�Q��٫+�'�~�B�7P9�wӪ9"t*�� w�����'�%RTY����0F�Uڻ��׽>㲛�6�����T�:����n Ջ�l��3MZ���+�Abe�6h"��<�#�)~R����h�YM
\�$f4uJ��;/O2������xg	䁟�q-�\ڤ=!��Z0q���Q�Hs�� ���H*�@_'�l\�r����u��W�a)��[����X.��K��C�G�{���a��~�<�{���ټ���~ /R#8:�Lݹ���%GUW����[e!K^@�"�>tQ�����k��[�/��;i�3�K�?��+�E(����W���= �c�,��A�=���5٣t�e˩r�2���\�q���5=�G"��R������KW!|�$��Xc��*��\���T/~z��U��:��}ˤ�1�WjkjX�d���@��Gt�%��q���}��1D!jI+�W���U`j��Q,���!�,�$.�ӫ�@��%GT0��sx��%�S�V SǑjr����!DxCc/��(�hF����*]�O�����m���C�Գ�%K[���g�6W.]I<>���t+y��R��秂"n�������|V�3
W����>7aZJ0���| Z�H�ކWOG�WӏCt���i�IfR}XGw���V�@�g����%Gss���pOy9���ƍ|Lm�`��V-2��ˑ�[��u�8�Q��3$D�|��Z�k��=D"#.A�Go�w~���:u��n-�V�T��B�׳"x�л�.r|Յ#�7�h)ˈjE:s4 s���|��d	�}W�|&�3=(C���W�h��<<�����@
�3�L��}u��;�/��|}��_���_Ϋb�yX���DQ��ǲeuTW�,�븉�0�8�j�J�F<|�M�]v4��t2�RT!'4#�K��ݔ��P��u��ڽL7��՞wӻ*a/�;
}e�)�t`� ��.l7%r-�1��geP?����r�^ L�H���N-0�Z���Y04�u���U�4�U���Ef�O>�W���'�5��ŀ=oEJ��	�	0���z����,��>T�*��H(�'���g��ۺԇ�n��$�+@��qL�>�)7C/���P9��P󈅒�����P�0�ѓ\Q�nz�����$8�zY,A䱏���#�Lo#xAA:'4\����8�2Sy����'����9A��U�¾s�Lo��/?1�>Տj3y��Yx�E��C��5���7ȟ���9�V�p'��b=��b_gog��8�=1�"b��p�r��#Ɵ���2�V��R�3I���,>�En�$���N\f'1_�Pa�&��mՆ4PA�}_�k4b�� W|�n����e�L��
ޖԱS���UEw�\nf�K��?��W��Q.����HJ��u��`c|߰H�%��Z�YW�U�y�O�HX��)\mՈ���G93R n�Ȫ��M>�Yp(/�ƙ���PQ?���IjE����s�E;\)��Zw$
K��4�B�W?J�m��C��!�+y*�Φ�}+�$��W�K�����^������i�g�y�Y�x�S���M��iT�u��j��ב���������������_^�8��j��R*�oUq}��i�G�����L
��|3�L��:Ms-0��d9)�[<�;���S�j	\�p���p13�+-����[�����*c ��y��Ԉ��,$9�G���M�|����l�C��EA���xʠ��6��
9�N|�#�(ie��]�T7��T>ǻ�#��鋙�H\t8fR�p�8���Y�k��7+�����/���!H��4jPdb{��3%%+�Q}1��V��=7MC�|�)�E��3��N��wo9!��
V"�O=�á�0��ǟ�g��5s��K�o�J:�÷:�T�:���4'��8��;t�(C�Tkj��5~!
�B1����?�rb��h�6b�#�5@�DH�3U��G���B۴��j��zM��"tDFܬ�����V0IO�%��3��ܥ�HA �Hث��q�n:]�+ae�_,���_zA&�<8:��|R ��9?��􄐨�OX.�c��:��;��.��fP3B0��5��-�#�F\���~�=7�����RC��ԑ�B#��I���c!����f� ��	����c��&a�	h!�N|p�o��]z����J�Es��Vs+BT��6$ߵQ��>��w��{�T%�xd]T|V�9��j�������3�q/_���0��B��Y*�@V�>ş�[f���%4,o{�X�xۍKȌRh��L-ϵH�l�+㸰m*�kq=}��0)�Bz�?	�����6�e�0�~(Ь�	h�Δ�{��.B��ɠ���QVm���g�� |e	�ߛ�cp�JI�e����]�S>�:g���u$��sD�A�����Ʉ��]��z�S#����D@e~p�+��t����]�f����w�w��W9P.��]��'�����)r]��u3�EVZ��z�S��p~���u\h���>�yL�\�V&Y��6����O�����`�t�?8n݀Jk�Ф{�npr�����'sX��Y�t�"v����7�lq%��&����g�J� ��Љ�⺖� ����
��w������1��}U�,B��ȃ*S���?r���%�7�����c�*ϩ��?9��&�ݰF��e�[b��p緄�6h�]��%��7(μ���b�.;B�	 ��C������\8&ң_�g�_����D��I-(��)�˜�k'!Q����h�yΒ\�n���e&|�OE?�T����k�Áe����U���M��)��J����@����qά@L������M+H��(?\:⵼��<�Wm3=:[/?@w�$��ਁ�Cƹc�#�g�����.��ô@����o1����ʳ�\>�j��b��������H�����u.u�W8y�{M�YI��C%�8��qZ{���l�!H�r�t	{�5Z}�m!8`pk��o��4�ϒ��{V�U7�ФЮ�<_uyX��� �A�3���P,�:�� a�k]�ݧ�֮8L�o��m�"'V�`�)_�1G�.�]��V�6����w�ys�7�Z��2v���1�Q��A�as���Ùs�+s���m�N����L� �ժ�4(iw3Ĭ,��Ko�d[�E��s��kڤk��:�9˯��"��M��5�+P����q��;L��)}J*	��?_� �C���CV�r ���|~���Y:� I��S�vc*U�SޟJ�C����i��Ճ�6ѧ&Rܽ+уO�=a���3�-a�����W�U���Y�����:����(}k5-�Ed
�+��Mb�����lۉ�G��;���KpւN�����9���y��W�t�tp��BQ�Ȩ+�_��sJ/�.�W�܁�iz�����G*����x ���ƧhS�?}��o�}5Ǳl͞C���_/������R4���v.���ɏ7�}���f��(:qR�v�g�u(�d���Z�x\9�� ��!�-k���;������8@���+�d�5�h��/G$���N��R�g��ҿ���V*2J	��͘jK�a��Ʒ�%+�A��cХ���q���MR�)���֑�@�<�q:�	<�%�A�4�jĎ!��^G�s:_��DS�\ǻٝA�דF7�U���aש�<�jP!���Ub�� ˞� �?C
�8.m͂��k(�/�x�Z��=>�у�F�,-�N)�q���4�l�:�6�X;B�q�_����5��)���u6f�0K�DH�C[�D�1�lMSB�YWcW�N�p�)~GS3��[)¯[��gJ9A�벭��!*�r@F����3h��lz}FL.��V��J����L��Ai�f���z$��Ϩ���%j�	����~T��{Z�&�`>�T�o�|��7SC��t�x��e%5�ePƺ��	�]�((�e�t��Rg���Y�,�JWz)��\Uإs
�Y������[��C�'O5�����'K{��`���[�Yj���`�L�74C����R'W��y�1�C^�����3���&:���KP#g�����>++�!R��ڝ�F1��������kh8���v���	�4�^`&�G��`�s�Gn+Vj����(Q7#P8�6�c7<k�̅if���f$��ˠ�����5���?�]l��+Gů	ٻ-w�ɷ�w�p�"�@�F�@��y'��K��W�3��T)��Y��6X�t:씐h��_A�$�-�)ү���o�N�2	v��z�������h�$i*@��;�m_H{;���X�U�(��/��kϩ������=o�S1z\Hk=>N�S��n����"����?��x�Xi�Z@�_d+v���M�2��o��ވs�y2OB��a$��i�o�Oo�/���dO��w�c��T�!^c��r�k\�	xd	�N����o ]_V�"�,�[�i'�I	��V����usA@�0:1{8�8�W�x�k(;�9�g
��j��1����q��	�_���8�eq��\��V�q7�s�1xM���
�E�HZ���J�"D2����A�&ߤ����:2��^��Tj��)C���j��e�(OW���R��!)�R���a�N~�Ѽ��b�F�q:����l�D�� �-A��i�|8�>�FpŹV<��`a;�������$�r1yo�
u�w_��3�T\E�\���6����͑n1K�(��l��+^��l�8���E	���5L'�f<F3����5u��3�����+0��14\����@�v!E�l�)����8���^��_d o�M�d~XjV�⺗U�.��w	 !��S���W,��gfuS���K�:�APۡ�@�?���u�T��\�mo��43�լnX��8�����`�gi)Q�����z�94�c�z!-�O����>�7�ֶ�RaO��/�����Xm���
b콴��~-�	(�d>+W���K r�G�V����w�Ad�l��G�����~���7�D�D%Hi��.ߘ�G�C"���8��wT-E�F\[�IV�Tr����~����:1&�B$�����z������82��]3���?��LL�g�\Dp�1��yKy�!dD��>�:SG�{�2��h�LPSo���R
��pN�kǟ���sJ&Za8�8�ۊ2����l�Hj��ڸ*�,��?�G�/E]�-o 	dR�*d����O��:۶�\L~h(Ө���l�wB������w�ႋ���$B��*<�K���ʄ��d��:!���qa�r��u���}�+\����mR*\J�B,rK�λ�K�s��P�[�L~�- $��9�Ր��h���M[\��b�C�%��V�����Tޓ%3�ybv�����8a[T��R��I�(�R�TVhQe�i��)p�$EE�zq� �s$sHcƱ���ǻ��b�D^�C�J�'��H����վ�Q�?]�|Nv۩��Cٝ^5Q�U
��iǨ>��Gؐ\�e�`5Ԧ�\��F�B�D@��i�E�4���sM�ո����ـ'��Vj?�*\l����1�Sa�k�g*����'$֦�?��;z�(��x���=���u�)s-�c�RG��:�v��r�b���*+v�0���m'�<�C���	�*8��<V��I��W%G\vI�O�����n��l�[j`~g�hZ_�G���9Sk|d0dr�^��p�üI.N0mο:|��4��	_&~Ɓ�{�v���/X
���֨7��(J+���д�%�o���8 O�bĊ}�ro�c��	����a-�h�Մ��R��@?5�3�}��;���{ᴅ���J�;� ܄y��4K=��H�?�<�P�~y���vZ	V/�!F�`:>ⷃ��3l����<�s5V��p��ŽJ��S������#xI�k]J��ϻ�l�xgd�yI�����|�\W:m�"`Q�	pn���]�k��!0�
��mq��8�DA�|�d������T>�׌���
���=��b�����f���iҏ���S�p�A������A�(r*���sF�a�X#��#T�����T�ӓɵ!G�@���D+��u<���<}�V�T۬%Y���f���-���?<%�v��Ó;wB3E�I�ݡ���i2=��kUƘ�/
pP6�����(���W0�`,�s��aN_!=E���l��^���V���k�C����3���$E�{�%�S���|�1�$==�${��OH�EܢSv4��,��Uc%���������u��T�����3�����ffK�[|G�oQ
\�Tt�<���.
gDѱ8����1�4'�p��_�+*Ç�K�L�?<埥�W�����P����0���8��)��IW-L�����P["���ۏ�ҳ��C�U~�ߏ��	I��y���4f��Y�`��"�T�ø�0����Q���O���ß>��?p��*�#+�A�
C�������=:�&�"Q��	ȈX4FH��Q0��,�U��hׯe4<OG
�����,1s��>S?T�ᚹDb�U�fC�yG��}K1���E�qviP�R*�ǖF�iO�9/$~�A�%�Z� 6�YO���a�ӹ8���oU0��n�KX#��	���t��>�De����� �T�� ��+B4̩���q�lh�ǅ��'��g�o0���M9A;Q���3�/����9>н��&ϩ�;�>�YM���2��M>��]7	���c̷].�x�_�Js� X�%���Y�ᓂ��]���/����FA>M<$-���ؤ���H����B��ka�D7

z�g˷�Y�FD�<�c\�q5X��TP�盼ތ���>o����M��Z���8e�@�^��}��L���#���a|41i��X},�d$wӽ�j�۫��#��p�gf"����CT���i�yNК�NU-��qI)Ҋz�����'UNоW0����v,ɨ?$x@&�.o'I-���k�4��9i9?_L$352�K�>Yu�G\�=b����Q�D�$��c@�CǀD?W�|Z56D
�ZQ+y{��2C Hd�����Y���՚Ck����+ayo�C7<�r�n���z�|�T3��Pݗ����Uʕ�7�	��&G��I������o��Pl0>����L����J~��������R�?�t����3@��_�m���$�y�Z�L,���{��}0p)�Ir贩�ȠF�����2j^~��D)Z7�Q=���k�%���	�tv��@�S��N���2�K9����eG�V��.r��X�7�p3������W[m	� ?������H7����(	��+��$WT���q�@��y�q6�s�t�X�`����x��D��Ad�}����(��v����a�VB��b��Ћ�KTɺ��\/�c�Z���8ź/`^l��zQ�/e0��7�%�vWG]CԤa;�p�E����^n {י�k�!f��96^� =*���2�L��Ù~�3���H��SM�o�0$w��L�Ut�.8��\=%�o��6U�:ȟϴ�\��)�Wq5C*L5<H���z��r�J�Fe{�P#We�zR'K[	���rє79���&YX�-Ͳ��D�ӌ��ݶ&��
b���.�,Ve�Zr�����u4^�3�C	6��̕�3ѣ�r�Ϧ_��9�sSȣq�̕�fe�rB�D2�1Y�u�T���=ӧ�Pl`?����qH$���S���{��n;heGZ�Wt��#B_K�R� e���_��U��rQ�;�LDI#I�N�����kh' c���(W���tnx�'+�p����C��sL��I������2�hx�N����3�$�ԜIS�Uu�7M�ʭ'���A�a�8s�_6�s��@܆Ѽ�xr
i�Jq�c�����j�9ӷ��K��2��A;��⷗$��x:�B�j&L�^��O�v����q�)��4�GS��ż��u@��d-)1�).n!�������yQ��f��c�|b�xNT��a�Y9��nZ_����6�ӌ����NaW�[TP:Y�
{��K�H��Ȥ
ks��^h�9 ��]y�F>����Z^�$ �R�b"���23C���&����G��Z"|�"�߯�;�3,T�5t�,��ר'�&籫1A��$"N:9�k;�4-^u�z=^3�sL�V{`��� ��p��t����9Ts�s6Uz���K����U��?��$b;z�	˰<�b��x)�f��X���ܳ4A훿T���7�Qj���S�cI�X7G��?'?���
�؀�1�x�T@�$�U翾 e�����"wKz����7��t@���f��q�H��X�}G�VqyP�f��p������I�HĴ� Ōz���ke=�gQܥZp�-1I�Ӱ�#PW�����"1�e>;Ӝ�ylIj̓X1c�q�玟��g�*���B���R�)��JS���s*Ya����p-n�z�&�������p>�KL'.�^�NϨ��/U����\Z�U�'����>�
��)��~$�'���������r����B�u��)�O�}?���J$�$������/gW��)�ۗI�����	,
����s�m�¯�Aj�hۤ�ԯ�T����rT��8�e�wR+>hR��;�{�Lim���J������zR����/�zRk�O�U�?��rI]�R�
�L��NC�>�V���}@A؈i�1	E{��/͑��D��B�g@��5Ql�Է�8}����XG�����]�`���Sp��vg8V��#YHV~�K2*~_��;d �8j[Xo^b�7Gt؅B�ӽ�=�����tk�L�@f�|ޭPr��.��%I�u)� �k%\&"�����E�1�ă�Z���~�m"�@m��w�.��ꋇ��ڇ�Ǆ�К�u*]V[�SK�,�0�x��p��`��M����%!L��[����4���a��oKQ����i�P��	��9�-t7k�B�ZH]�ît�vl��i6�TO��
k��D�J��e�)��� ~�x�K��U�ь�9Q���a,�����j-M�+LbvSJ�m��^\��E�3��`��Ⱦ�
,��Y����,L=ˍJ�6������m����b�5/���C;�Wm�x�꟨���j���y��Yk�G#�Bm�Ł?A?�|�5�q� �7tz��5
E^�w���	c<�fQI�]�bvŚ����F0��S�a�4
�����4Ŕ��Y���a�>ƈ���VXi8�;ؑm��-F	x	VT,m�P8O��@jw:&Ր.Њ��7!��rCpY�--Ǳo�\�~�F��!��s��� UƁ��ƶi*}c�p=�K�w<�@�.��� 1x)�M���)q��X�����>�����eo'(34H��ڢ�l���������]�U�K]��?��pd�)������x���x�����W{07��C{4K̭~��6�MbAsQ�S	�M�n�E3���Cxi5���z��G���'�V|�5i"8]ID퍕�U(�һ���BE[ޢ�N�V��7̣u:�@ޠ��ޡ��%΍�űԭs��q�_��.e*[W/�O�[�e�nK��N>_��>��F�^�g_`�Us2����ګ!V����TA9��'k��q����R�^7�w�𿇵k��β�=�ݸx�|냮�����BSn����d���%8-qw�.o3��'��T闓����`AI���!����jXŪ4�g=I%�_�f�ʮO֠��4{�u��@�-)�y~���s��\�1��o"��@\�R{���,K���nd�3�uXJ���22��nh_{��g�`�W�^ɥH�9VD��
zBx���m#�ִYt��eQ��lu+:��㯗��W�I� ���`Y���k�g���fHvjg�@��􍵢a�c4�N,�5|u��敔��ޭ���_U�̧k~&`l�'�kh��@��K� ��J�Y������ۄ���"ns�+�=�#t�ݝ��:3���v�d�F
��7P���xN�����.�V#OH;�/�TG��Oa�J��ݩ��Ձ���Eћ��\r2��c7�$��!,�"�w��h��N��"���8��_�B��̫�ڊ�B�2�4ɅY�t]��na�a-���. �q���a[��S�W����j�l��Y�S�4��P@\�-��9��n>9d r����'"���WЏ�`�K~��g�hA�<p�g�I/�k�z�C�p��G��܂a'S���������7�>Bc���C��+�/�����x3���Y+fZ5��M�B+8j3�Z������Z\U���.K7֎ǅ�ιX�E����":,�B�U�0&�GSj����J���0_;�w����K����U/|�7�X=e=A@VW�2L��b]"~Uh��t6��$��\�p���L	ٓ��M�ZW��P�6����eRJ��-{�d�m�ߍ���Gg^�����G�T�����f�9�/�*u�{�"@ႏs���"id.�S��Pܞ���rY�YK�&I~����9�49���I%�q�����2
X�yC��i9ξ��Z���L=���%�Y��l���J�똤����������I�g���EC���?KF���C�t5$�� &rk�6R� ���gF�=r����[oɮ���Ala��]ؽK�szбN��T�D6=/)��v[���"6�z~0[�#E�/�M�	Ƀ��H����x
-�qsv=Ðu5c��:�b��dL��x�G��o�6�se��K�j+��s��i�O�i N��LL�-��C@�]ytG�`i�n)����+	�9AN��<l|OdW�as�i�#h���4�Y��:�Y#��j�V���9E�	ƺ��ґC��%N��$�zUW%��Z&ng�/��d17�&�IxS��Y[����I�	]h��͑��G�q�{����"o/~[!� 6�o���G�oZ�����Hrp��Y��5����#}����&sǄ���� ���j���yZ�p��Σ�v�� ��# �*�K&ꭼ�:����v(Zh�4e_��۞�%����zt-��[8�_�SF������8o��!>.
���T� Ԣp��q!�idIkëʼ��	�C`� Rƫ��(޹�f���7�dh��`_sf�^AV��q��Cl��>L�F����]��N#�d�բy��Q���!4��^@����t*�����'W��&%�x�-���׫*��=@t����:���5�&R��&��M������9��MUΫ��2+��wY�M�.`&��r�կ��^��	L�悕����XB�tw��㞏+]W�;�\���d�J+hX��v��@��2$G���W5ON����*�A��BĔ"�Rg���)�o���j}����|�a�)�N�(��UU���1LtQ-��q�Z/V�Fz>�� 4����Bw�L���xL����hm$���k��;b�����}I�����6K� �>��=����Dua��u��R(��x���Ս��d(�d��!R:�T�?�/��	��Ɗ��c��j���IR�o���;M$��xm�"�Ӟ)	3;;�Yy�2�r�)��hW�i�ry�Z�2���H^�U���Mx�T��>4A�\�D[�nC,�'8�Rm�I'�J�щ�k''+Ji�](� ��\���vՄ���LJ�@�z=e����|�O��֒4�, ]� P�����{Pr���_B9��l1�a�� @gL�I���s%�H���o�પZz����o�*;Jk\:vC���|31s���\�gs�3��r�8J�Ec�f޻����b}ŏD���^�^^w@���3n��7?���#t�ڿ䪌u�XH�T�P�\���?�+ٻw1{ *�_qW����aI|��*�g���B�J�Ӯ"���1���q��V%<�{=,��t��_�"��k���lD:vw�^F\�2 yኰyQ2�\��xf�<�F���6#��;��ؐȍ�a3?����Zs{>�1%8�!Fi*��7��V��o�%�� ��&�V�)JhK#�R���&�$o�	��|ƅ�CՌ���lc4�b��r�]^��Mػ��A������<����s���y��!��i��]9 ������fw�E��14�����ǟ����S��>Ե�ϕ~��"�4,(�^��k���.������P�.KM�����Ę	鐅��/J�6���j ���aW�*���d����SKQ���l��ZY�xn)_\j���f h�VC��#�s�����]�G*&�C�Y$p�w�bv���,dj��o�B���a5�!}F[����X��ї��+����iy�b�} A���bOD��4	�%aS�-9uth��	�rEr?Sg�[��);�j��U&�����O/:b�:ǈ.%	D�w���{���Y���� ����؛��V`ޗ����#��<�6��T3�)�em����%��OR���qs�S�#��k*�H�9o��(� я�����랱=e��t�,s�$����=��`�)ʱ�"���G�ɕ��,��`�&�mO�&jM��u��4�b��^�5�����f���"�G%t�82
�[���XH.&<I�����־���yU�m؄x�@���Yޥ\���v�Q����T�J&FiPS���{pZ����%A�4>A}��q�HOFV1���#t�m��^��=r���PX�!\6*؀y�,,��h�a�y�np�����]��.�p%*��Hk�[�A}��޼n��1�S��F?�:�NEQ7?u��։
�������Ω��*��R�]�|m�*�˩:%o�;�KG�a}0#N�{K�Hяɟh���^S�Ib��哟vv�@	�ij��u��Ya	��T1��{�������]h����+@�����FC���#-I�rWN��=e���)o-v�=B9�_Z�����T��D���6i)7�m^��8��B�	�,��x4�mOQ�V6=Ñ�[ۨ�E�4�P$�\�L#턿(�6S�%+����{k��cc$È7B�^S��v��`M�6sq#��]�U�CS���Iŉ�<qH)���#�1��.u�G]:�1�?�Q��|fWM�@[$@I���j2�>4)�D��H�y�"�P���z�/W�9�������|�҇Eu@�}�/�z����)1���0�Y�_&
��k��*�}�ߍݕ�١ [ݺ��>"v=򹭧wM�blOs���9D���M0���T_]B V'�fhs/�c_"�%�O�SO�k��̰X�U�����>�G��$�o�W脬����߉A8h+��Դ֋��\gפ�#M�DX]��yt:a��M�����sS���Ea=	������H�F�j�d�v"z
�����ʫ?Z��Q`e:Gc�eu���5�?�ڦp:�]���yTu�k�ϟ�o�A[U��V���k�r��\����n�� l��mg��_8jv�8��΢xX0.9��U/,S��;�E�W��WZ�&�F�tu��R����:{��;�֫,�,��=�׵�}6����H�C��7"�x�oF�C������k��eCCN���/2���\�!����{'N�#�;0\��Ax�,���P����Ă���UY��%�u�ȑ��[�+�������f8�(u��.g� R_��>	=��]�R���ǔ��R~Vn��VE��Q�<_�9�\��FV�ю��2���h���'��pE}z��G$�,V�>� ����ʮ9N�SR�������fO�w���}��;]����#_A�nq0��
�n~ӢL�D�A�
� �.Y���ۺ��7�H[g��������A�`�ν�J��rF�{�X9j�"��FO㾫�_WG��YmTs����x�Z�EXc�Q]��#���/�f�D_Tj�<�6	���5_���V/�����w0����:�$��Qo�z���\�f�+�}BkS�4�3	{���7ta�9J��|Ɔ}�ÌT��2���vG C�ޓ��m*p��x��ؕf��k<��4WJ\i��+h�����Ҷ3�-5��#5�1�����8I��PU��!��W-��E���6��URf���K�:�fQ.�`_"� V�N`����B�5����;��D詂6�}�Ԗ8�bb�m*����	��m)Vm��Vp�m��K����M"T޽l�-�p&M�zd@Ac�M���W�J$�8��Oy���沴���aԥ@��zN��X?7�����AӦ�t�A���<�=��)�f)=�}��ܾU��� �NŸ��累i�}Qs����������(;�fZ���V��ѭ�/KS2�w#�P��>݀%�0�y/��1��m?d?���aǡ�Bsl��3_+�m���)�����}%E�j����$�*D�5`�LYz'W?�x�|�S�/�#��]�Q`� Q��R�<p�s�b���/k���]jLH���Ua�T��2�{#�jT�"��d�Ϊ5�J��ц�� C��!�N
�6�����rIT(�y�*��ge_�u|�th%J ��DZؾMO��y�/�q.J�k�+��W�Ϯ�s[&����%�v��S����g����H�꥙�aT@�I{6|rq-��n��r�O���E6-��@^�s17|��{T^^,��9U7����X��1��µ�1���Fa��)Uc�%7ޚB��v�Uh�wn�g�Y�a "�� *P�g�Y`N��5��kI-rФVg��c��I��׃��
6����p=�F��~�7S~���$���/Y�-t���G^#"Ծ��nN�Fx #���8�`��~�<�)��O_|'���OT���b�q�
��2M'��?]�R����e���(�O�H��`x���fȆ��0u��"g�t�����{t�!�rj��5t��\���������������H��vJ�G��%%�冥x�>�s�zS;G�d8�6�t����	xo3e�����^>^���A��2-_��G��l:2�.�Dw7� ��AVQc��=<`iD��L�ؖ2�އ�G���2bh��)��/�Q�H	O"ݻ2Ŧ��1JƠ���|ĵ́{Z�#�)R�ȊytmZ2G]��+�D�j�RV��l�0���h�&�]ڤEV�å\�T�R����Q���(~nn.&+�O�g�0��յ�	��� q�罜b��8[U��aՇ"m�4��er)���S*>e�l��ɶch �R�g�ҧ���>���O�5tb�2�IQg�">h��$���Eq�D�ҧ�ᵡdC���yew%�gG���!Ys��[ǢF�8!�̧�Т��8(�S$FnY��i�kPY���Ŋ�{���6��֏���C�dueuE�����ґ��|\�q@�.���*�DۣZ�"��WӅ������Z�Rk)��Hl&O�;����CC  ֭�|���X��
�&:Km�a������dB׈6�/=&�>��/G�� �}P�w����m0�ֶۮ��-��I��M��X/���g�X`S(y��9�Q�����%�ؾ>0UZH�|>H��*�2��Ⱇ7 �Ce�N�Qg7�j���-�jw��Q�K���Vz\H:����-�^��V��r���Ԑ��Ō�����8��ڒ���S%���:����4Ft��Ď�͇i�Qߞ$O�6�ÕRa֚�,ǵ��1�ݏd���v�"B����]6���L�7T=��s0�:PaQ2dypb8'=Ϙs9��R7��B���m�+�w�i^6�|�]�uZ(Rr^�_�����[��W��˲��;�}{��L�� *����E��_�Q31/��n�ԭ��A鱎ӭU�4ǽ?I��!���/17j�ݲ"~F5R����g��y�M��7�cF��s���p��֔�"O�1q^�O�Ki�~�j��l����p#�Y��wg5gv+�1�]�S�c��)�IJ�݉.j4Mr;�/t�վ�fZ��e��o]ج��f��^�F:
ȍ�J�����5ЂU���e�%j���#3/�<�e�E��D6�;��������
)��@� l`��-���Tm�q>�2j옄��D�C�St�=}��V+�撝 �Ƽ���E�ld�����3c��k��X�:�_���ؓ ����c��~�-'ՆT*?n!�S	�ć�Mخ���**�̛���>h���q��/�aA�>�V�,�nCT3�6ɹu�0>�'*��!���b�����������|,X��e'aeK���7�1�EC�������'��o� �Ώ�q7
*"q��e��Gg�/�������Y$���cdF�G���~$���|�+�`��%:��,�~nb�~L�h���g�㹭/�͞��N�U�^�F6���.e�jN�=*O
-"D���b�`��og4ŕY��g��"?4|��[!���iw�)�.�_���������D�GŠ�	*S7�r��"���q�=�^}�� Z`O3������q��/b��!�1�l��=DU�%�t��!����!<��·`��G��pvi]=�Z9}ɱ���| Ė���5R�C�Y�j��R�R����cO��Y����ڡ��JU��W����r�������^�Z�`�m�����R�I�~���
6���§���H�����LYt�	Rc+�`3SSz@iQc�n�v�0g�\B�<"��fn9�j٤����!�I�I`g�I?���{l�&`��}�b�K��ԋx7�=����p��r���i�q8��c3�}�79=�ت"�P���D�0L��
D��港T_���Y�����^�����$B&Z�&x��Ix8ni�[r�n��٢Ԟ��V;�a��xC�o6;�&�آ�u��S3�\*O��};�%�q'�#��#��	bQ;R���ɱˡ�J&�1��ݯ}���e����r��Ĕ��e�O��>�:��SJ�G&	�PY�(�<�2��x}����v�E`��Wry�&f��]E����m��;�~1"td0����1YK��Wo4)��JP���-e�7�'�S�H{kCSK>W{��c�w����T�A_�씙�U��G�2oδx3�s��Hݣ �k�~0���� %�:���[՛˅�z��>e��+rh�BKQ�Q��w�mzv��wS䙰H�*^�.��֑��0�E�{'+��I#�'���	����)����H%Ǌ���F��:	�a�Z��b'�?��;VQ\R��r�pQ�ar��HXk z�cc�_�֒":�n줼��@����>6��P���S�X��l=Q�`��U��.����`�g�yI��Sgt�h�떹+*0��Y����Z���[,��)���b��l������:�܆����%_�fmv�A/���Cp�UA?����Ձ�[��p��B!Q�Z!l��8W9Fp��1����v2�t�)"mC�֡R��;�R'�to��E�ǶSSa�d8~{d��$H�w��"Ng(H��_$jKtla����z[�}̱M��	�CPo�Mzʵ�;������پ�������ѿ8ۦ�
�y���π.G��d���@��\��xG�ʗ6c�j����!(�$�oƌ����c}H*eB�����4�|��L'�J���o�$�	.�g?j4��>
�~�6���w]�|�|��+��g�w�-n�RW�����6X��]������1������}�e��	o8clQy���{���)ʅ6��CZuӦ��b?�I}�A?�m\Fø���O��B˜��p��Y!�]%kzS��}�qc{��uF�����t`����KS��Q�i���ړ?i׫A��te��R?=�|a�8z��Ȟ���Y�#�p�|;�)��Щ��M�ܕ����#�[x�����W��p�:���b]f��<�Ч�� ��fGυ�Y����x�I8W������qU(mj�]�!��Ӯ�x�OrT�K�$��6�C�gȻ�["X���U�~fJp�ᙲ@y+*,�F�'u+��ҷ�W//iP��SO���@����@H�(� \��5�Րs�T�3׹�0�گ�oM�a��d^ct�]��ʗV!#Z7N�S�Xʇ�	�#x�^[����כ�^+bfA�Հj�j�[j2���jt^�˱�~E���F�]ߍ�l�eZk:a��U�+n&� Xz��2�rc�.cD̰��v�ƺ ����`~
d��	7��Ht���ID�C8@�^-��9���J��fM��6N69S�K�I�\F��| 3�BJ�(G�b��7�/	�|'� �@�Q��a�o$��5d#iu(��	i2��粿�Xb�R�C6/�,q�ζ��#4�`�U�ׅK�]x�C�	��H��%�EEJD.�w75�{#�1��mh�(�egyE-�a?�ť�����v���=�0��-��~��zrU�����S����SV�J��v����7�o=`�[ל�h��ڏ|%8�ęT�����RCE,�8rH.���^D%=6o}TV.�ŀP�@���
�{7���� h� rn���w%TN�A�)�I.��9zPU��0Aɟs�2�c<������M�ci��ȋ+�OY#�����@7�����,�=��j0�r燰k��|�4E��5���b���Y��J:����)�3v��rQ��[*���f�Җ��5O[&��W�M�r��J���~E�{�t	㵚0v�j��r?I$��X_�ܜ.��}vk��G�)K�,1,_@����|%�_V�����Y.���s���77�u���{�+�oڒC�v*����!N�����dK�	�0��]ʾ��J���P]�=�t�!r>T�Ï��i&���e禛�͚���ӧ�Rl0x`X_��ՆaB�Y���XM�I�*R�Uw��}�&����mp̔�ͣ�-kH͡rW�������%��5�?�Nn���A�2��Qp��� $,W���F�A�ɮY `;�M��/ӭ�!m��q)CZ�X$Ui�c��6;ͷ������*�ª�6�,m���5����4 G�k~���������=FOV�C�h^�Lx�G"�(5yј�q����G�j�(�ёR�$���N�gE���Ą��z�rbr_�����+��g��&<B�S����-�|��e[,p�m+Ǐ�|����O��r�������F#� *�ӧ�M9c���`����r�J}����BP@�#����K�()D=[�&k�8;`j)� C���f�d�3\_�t�˰۟ sz����W,1;ǭڌ����L/5�V5Kˎ��*������9L߹��	�JE��1�u!R�p�X8��m��9��s;�4�'H��P�T��G¸���g�՝#����|�%����)�$K^tf �K��<~j��d稢���bj�	,�"���%��ް���B���1�S�퉌]r�+��0�#��m�]�l�f��?��k�)��wr[�p�r��;r!s� �	`QFÅ'����K�kZ�ô?rb;6%w�l��n��#�*����c��+=�Vm�)Se�vǆƋ��/J��@�UOm�AL�9A�������tE<�~��	=�a�=/�/��0zu0�>
ot��+��6I#2�{���ӌ2s��2���mO1�;)��T�!���ǃ�F�G�݅
CF�E�o}1���ׁ6����g��+/^�S��to��i҄�}���Gw������9�����tf�����fL����4Y@R���rܦY�|$�Vr�B��c���ld_%b�gV`D�G� #�@�N*7T�4��#��?��WptJ)���x�֕$k�0�:���h�]TMӜ�a1�ͪ�f��c\�=�'�O)�@QN�^0��x�y��$U����x&�}1�f���D��A��&��+��W�|�n�0h�kQ/ay��\lv-�cVJ��X�y9�� .S�0�Ìp<0<�ܙn��pV!Y^��u�'2�y�ig9a5B��7c�����i��(�o�Hzr5{&J��0���.��DӃ(�Hx$�Eq>��{��v��!���K�Y�w�(�݂�)��ڨ���'I	Z�Ҩ�Z�GPqf��Bf��ϐc�N��&�H�@�p`�B�X��Ν�?�Y��d��K��/�*5��5��J�18z�'�H�P�˪�{�y�Ku���8�B�[�����cn�Z�,��ר��GN�<=hv?�Wgq_Pg��jN�8�棶�vG�>ײO��v�OZ�v����Pv�oPXk���ߴrC�J�qp�-eJi�J�������޵��9{ s�>��H��Ϥ�!h����ߓ%�r�z�b������(6�90��*3p�r�I�׽?I'J\�:�X��Y]N��H��.��bSu*$	��HM�nC`@���>|���N�(w<:�N�O��9W�%��5(��曢鰍Hys����AL�%Y�mP�l/����[�Y"�|�v�s����&��b��m�b&�U��$�?g{�{�>��#�claN�P�K����΢e��JCip������0a��IbI�ǡ��k�4\�஥�4*�-g�Y�*|OR5��5_��z}�K���A��Bq��(��!K���߄ ~�����7ǲ�x�!�U��F�sE��KJHS���|�cp��j�jf]�aQ�(�OM��>u�!����,؇�
�,�~���F���K�g�ֽ��g;�'��1�#]���Y
&�1�32RT��v�Q�@�5=��>T]�|����S��{�r����b���X4m����m�SӱP��)g�sJ%�!��z���u�zm��νx!�2�`��K$���g�R�v2V��Hj0�sD$]C9�#���?�@z����#m修>*��D�����ͳ��u�7���8֣�	� �؏+�����t��m�9�n%㕠�0�Z�Ux�r���!������$�@���� �P,i�߀�6�*�2-�M���z��(aA]bbȦ��W�ڙ]�Œ�s[��T߰F��m��'�5��#'��'�<>ًη�`�'�ǵ!d,c�A�/X�,�UI�Y2�����7lWI(0	�~��F�E�����P�����kJ:���,��95���E[��(�F1R�Y���c�p�NԭH9�Ӊ�C�������=J��E�,3/���*���gj�#&�fr\Ȋ<R��Y|3�q���[�D�q��k�ۄ���l<����G،�I�6�ųVZ��[��n��|�~��A��@^~�>�a��$U�6�1�Wf�QWj���F.Br���\�HS���󃃓�{�߃������=�o����&NC]���᭦|k�k~2�����r���Q��Qx2FN����$��?�ߙ<fKq�u��n�j���,q��]���[lI����x�b���0;%5ՙ�Y:�\�ᾧ�Aԗ�lܚ!��R���C��J�0H�R�h�<�{�������Eq��
c��h'(v0�'��a��9S>2y*<�Bag���h!��Q�"�ƐM[�J���Kx�����Z�t��4�7g���<��w������L& ,~w �R��7�t��=7���>���|�i�]-��&�#�����L����O�:6�4�N!��(��`����x�r���>!�
�ť�p�0�6D�XO��l��ϗ�3�ݖD�h�u��?@��؇��P�~�����O-"��W��*؎���v�N3a\�V�.2�ܒ�d��VU�| ���[�1#����I�צ ]���%�'`ΐ8l��=�`_ߞ�|�NH�����Wad����þ�u�G�4��q�tɟ+�x��s=,��UԬ�fO��Tw;���T��h~yM]d��*WOX��4����`�w������l[36]�ra�"�E� ��R���E�RYJf��nS|���<�L�C�#7t  �S$|OJ,M�59��Mo��"�#v�ʢ���r�{��M��q�	7�<�񺣶��׸F���1B�]9�e&t�аG�J�Sg�|�8���iR��h�.�d�+x���=>�<[�-�<8�����s�(1�7�d+~R7����Vc��P�$ ne&D����m�ੂ�\S�v�ԉT�K+��t��#F�-]'��4O3虫���Ԧ]n2����n�/T�^%luڬ9(,22@ۤ0r�?��o{:��!>?e1�����H�����������p_�R��Z�t��3+�`G9^&./	�5=������n�{ xI&e'@�o�6�kO��S��J�,I<{ �6�K�G�a��*#��=T[�Ǻ0���o���o�&��.��|��H�JώfϏ@��s�����X�c;�л�KL�|�%�M�쌂�t�!^,)�=��&�K�`��)3�;�ҋ,�u�V�%�;��'�c4���P�&�����p�ǺL�h����i�Ii�#���~�ȩ������|����J��6��fvz�vR�F�7,^�j��Rò�$��7ҡ#re��'J���T�Qn������RD�
V׏yF)$�Z�	"��b��s[�u_�k�ԔT%R�	�Q�x����p,˰�v��݂�,G|.?��^���g���T+B� ���`�)��͎�|fu�
4jL�A��*�2tSۣa"���ۯ��V�C�у�����{�.�����}7����uMἻ"��Ge.�f��3����D'�=T2T���g�%�~>�Qf�z�^1��M�{��B��҉�Q�*�� ��o�F"7�N����Ԍ�{Wo!�-���0����o@�j��>*А~�)�S��	tQ�0�*Ln�w��|�@fs� �)�\�3u�V�H�7�����ᰖi��%��)��k�5��uC�.�r����/�?�O��=
�Ddq �n^���g�pN���Q#G���c(D�~ q���/9;^@��_�2�^c��ӊF ��*��_����\ �ڙF�.� ^=9�f�j�X�۟��Un��(Zϋk�y�cs�S��σ���9���+6}|��/x}[�'�G݂	C�B���Z^�ISy�b���s;��&��bڽ�ٟ�Ͷ�a;�Up�;W�:�4�i0 � �8B������/yz��7�z��n��UG���˺|	�4��)2#Jl�h¼���\xO���p�1\�N[����,l�����z�`�T4��/��bwyE�~���f���'4��*�P��56���K���:ZILq}�\i_��c������U�������9DA�Jח�F7_����C����Q�A"�D�~��������k���/���1x+�
fؿ��̟�r��O����N>����>-�%�]���#�y`?2O�����u�Z@���Yœ;0�+T��Y���HIa�s1��^���,Fwcyh�wdNr�G���S��F�m܉�]��W6����a�j�[�Zk�\z|k{)	��ᑵ�}2� �N40�����K�7�����>l���0(�zt_m��'t�	��`�`�b6�U��?��k�B��
_E��Eݴ_ r�01^E�<���c�+o�`���#m���1����m���-�2����g�1��1��W��d�M���?��X�H�Ͽ.�P~D���5z �T�J��F�x*��x����==�h�S2s"�ܜ8tz5�o �o@��!i�֒٪u_����Q?�`�~�W�TY���绅������0T>��?پ���IAa�"HV=�Ƣ�l���2��\��n1���Ǝ`��~iʹA���׶E^h����?�6/Y����p�]��#"���N�qf�G���6�,+�'}=���%і}fO�b��Z��)x���X���@/2Ŵ�v��c5�E�`�]hh�1���ۚm��x��-���������v�^���h�� �B+g�҇#r�G��Nc*�N�`YP	���Q�r6����t:-.)����N r�Y�E�+�O��q���
樠	�ېJq���%`%��� �~D�v?�￻�S�t>XH�_�M������"���v}�MS�#O���yMD||n�,E��H��B��><.NP^� ��lK�¡���ZFP�g���fQ�[4=N������m1«�K����~.��)��W2�u��]!�8��3%��xu��laT���=�hx�Ƞ��~
��̉@��1�P$A�xU-d�>.r%���G��u`�;�p�0X!���i ������ްb�;�= n��پ�x�)w�Zh���ְ�\�Ez���?����=?�!{n�Q�����
� ����Y�s�1$�X���`c��C4s��L�'y�y�fZ<W_.�s�8�B��'�]���嗲p�ܑ��8{bU����O)y{�臺(�<���ȓ�W����R}������$ןj/�(���$����w��z����ȀD?�զ,��Ʊ�m6�B܁����y� ��6�Z~�,徦�D���J��X�#�,�Y�|����[G��U0��N�-k�ro�.�{�n*SB�TbͦBb{����#�f ��~.j�����!MF	�.�ׯO��~��Ɇ�8��Y1To���=�#���7k���˼�!��xsx0Y���Ǒ�+�puŵd�ՀZjL��Y|k/*,�~~R��&����1R�X��\��[�h�w����灇G�6���C�H�l�J@�]�LG8��to��YZ)[g��2UC����i:d�\0%�w皰��YL��w����Ts����j���Ifo�D�r+�q�L"\n�ȟ�jS��F��;2�bqՅ�x4���c+$����X�@^���V&e�f���_$�cb��Zi��¯�d�CPf�^��i��R�d��0�x��M����E�O�Ci�ZE^5�*��icȈ�&�u�}�4��F��Y��I�����П;n�KE�x�$������u�/mн�
B"2��]�<���(�}��s[�).��w�p�TD3�n�=Dy{+M�I���ĭ��j	������N��i�9D�_x��]���z^�9��A����+��G���Ɍi!c}y8W���JnKֶG��;��yf#���N]����7
R$����9����,͠� ��c��l�����RH��t��p�,�H��\+�qC�-\I<���Tu�rd{r0���T0?%�|(�� E��
�nc�?À�9ּ�4#]qk5�t�¾�װ�S�͎��i� 1sV�z����3&�"�T>�sOb\���K��z�Arv�ƍ������6��"(}��c�V��F�$�rH)����s��!�с?E�RUD6cՆ�r�Ӌ���t׉�������X��FT�3�a6�$-�)���-����ɓ��C��!p��D�aj��i�A�Úh��Q9n���>�lwG���%�������(����NclY�v5�}�#���UV�4�.�0���W� �iFk�a���.�?����������`�"�`����ϲ�$��@'��4��� ��bo�s�)%L���4^u��~����
WEgO�{�f�\����1����a�Ƃ���σU��ᗅ/��c%53�\"(JwXT���u��W��_$�K߲7=�P�w�H!�j?vl��S�B��_Hn��'�i+hL���i��=$���H90[e��NhP��m��g9�~#�o���Td):�����u�I�O��e�8��O���C�lfg�8��l�w��"���ҧ��	~F�S�j�"��|8�+�1C틤;�ʉ���y�z���O�:"�Y���� ��-���0ۿ�C(�T�e����4Q�\O�ZU�8�r�@ۀ}�ý+�~o|�"L=�`���`�b���)�Ū2�u���A�������O�?K���~̭���0�*�J�/\����IOsEP�YM�R����]�G�>B�[���fOu$l8�`��B���X��Y�cj�bj_Y��7��V�g�p�m�ܫ{ӃjK��x"���f��j���1�[ڧ�]�H�ɾ����mѝ�G{�8�����8��\"�0��mPk�𙋗��z�����C;��s-���'?�O�a����u�8�=k%�B��u4<J�������o�Q*�{-�� +s	��|ݎe *����͎l��y�3����0���E�Ac:���.�V2E�eiE.ɶ�q���\�����M��
J݅�W��v@�F�QM�0$�뭎�F���=��Z�\�[�[�U�� /�ً����i=b�SJȣ�w	
Qꉬ�V�OS���"N��,sw�\ב�P�}��l�
�'�o�uZw,F�hSM�����fI����+ ! 3; �r�%��е�~ܚ�7BX�驶y鴄{�X�� k1Yf>�d8	$�����ے�#�G��gg����k�
u���t%��υ`�����F�H��x�.��DQqf[O�
g��QG����)6;�Jڝ������ҭ
{���C�с���g�Б�Ĭ�{�aK�p�}0�&r���j�8�!�����٘�� ��$I�d��N7l\櫠��6-eG�%�?=1ȶ��!�cAz��v���8���5q������+��Tk�7Ս�d����^�B�顖:�+���z�~��s��Xc�R@J�Cb��Mv��*�~��
�!�}u�M��N��K]���# L�5l��SȰӯ�!;5��j�N��:�$F�����R#p�ݙ[� �z�������6�`��F#;a �t4g��<���	e���u'�H[��̔���0�9}����|�����L��m��)��2(r��v��:��w��kS ��X���Ҩ 9CO�K�C�8�-������!Pz����"�TL�Y�e�?*��&4��`��6,��%��5���Ў>��;�^E���E6��	T-{���ط3���Y�e�V���zG5���Z�ىy͕�8�W1-�� a��a_<�P({�u���47;��cڳ����J���F�ę��Bv����w�A�@�������js�ZW�oK7��b�L;�<Ǵ���"�ڨ�hkIYɋ^C~ST~A!�R����nD @v��b9�*���pa״�ú�˼�{ih%e��������ȋ�2��b������U�O�Ӂ)q��2�����-܊�L�IJ���;��]FhT� 9SǊr'`	s����n���\�a�݅�d�5����x�um5 ��~��d)>=b˳�UG�_.p%�P(����R!�?��2�V*z����]Z�yo!��53dͪR�F�v������,OM�7>��;bq��eg�6��H���_��4�o�8��Ԅ��G8��C��vL\�����#tq��i� {�����i-p�>v����b���Yq���H{KtN;P�2m����lM��p��JV��)s$W>��	�P���B_%�w��zD�XI�	��u=b�^�M��T�����Q�t�j��)VX<�h_��U�~�9�+�&\��F���/B�Hk^1k嫪�(�B���!��K[	i���C��ǂ�!���M�]��W�l��������9������H�yh�"$�ݰ��(>�����>D� My�P� �	�Lj놄�~3GֈP;��e�w�'��*��J�W�1����&��+����F�e�r�Z��a���1��XT�̋Kw�6�0��.ōکi�����G<'�1��+��>�����7F��W�ϊ��!P�Yg�5K$�=�Q�Gl� 0r���.�jqT:���qSq��r�򀛚	I�W�#!*/�����	0�_~�(��3dT��+��q�X�6x~��v���q�;�7�xN��ܙ�;H,Ӳh��%���V_j<]ת~���0�;B�A'|�_�hg�%qE��(1����>����{=ǉx�]#�s�b?�*T|兪N�
l�	Z��33e&y��]A��LX��R��O �@q���x��n��;5O>�ΩO�U�@�zA��bD�J�ZJ��ܗ�\��uwM�(���5���jiX���uTA�h�<`�1��r�,5Y2��5��9���Oꥐų�-�t�7�v'�D`���W��Rl@�H%6���'�}ޭd[}U�^ͯkBs� IԾ|`���жE�1�odU���Y���憴��b�g�f{�'�Z���zw(/g����T���@�S��m��a{�A-&83/(���3��1=�r���^�N�[�DBЅZ�6��v�k�B��g�+���U߱��@� �f1:g����∘��G{EbH�>m3L�"z8��Q��)I����uU��L�n{w�هO�����)O,b/O����Ri�0ØU�I`�G�Ҿ����ȡ�Ϝ8U�>�(�_y0q���B�2~N��i�=�}j�0�8R�\����>�C�v�UB܂�P ��Y&_}��(+B2Ң�=��lw��몇��M����_s �G�d�_�Y���s��+0kFM��~|��˱�W�s�X�^�{�Ea�z�z�X�����t�-G��ƀe��ڇ�c��w����J�>���O��Y���]�g4��⼢e|��j�?���?�?�+-�o�+4U�4}���J}a�L��j1����l���U�T��� �㘎 �%kv�jS/����8��"L�'���T=�ϾjO~nҚ��!��$�,&����m�6	�ғ�� 4�e�)tP؃�q}��4�%����|����ؕ�^���/���Sᔱ�4��p��Y�?G\S���0O'\�z��|Μ�����I�K��mad�����9:����a�+�:��Z5t	�����s�k�=�+"<�������0�;r�{̮K��j����|��bS*��.#;��n�f�n�0��("F��D��X�����/�(%�=�^w�r|�l�|���ȸ#�:fE7E�M��Y��]Q�T� A	��0K/Q�C�o����n�����_����}�B�+v���u��9]�.���G��8��o��\<d�]ڮ���'�ѓD#K-��,1��9��!��-^�`B��2K&	��)d���vKz���S�¨�l�J��j��*�\��+����F��ߵ�W�Q�X{�j}|��_�?�d)�}.�Lp0�YXF�_�t$x���
4!P����n�:��ī�Vf��,��	��I��O��U�x�Ok� �4P��f9:�s��[�ّ;ѕ��hV
uG�]Q��S�@n
F�<��p�]�Xp|G:ǔ�<
k=N�)�=�R�`8W����=!I����jbx�&%A~��D+�4�`uR����rh���د'׸�7@,�\S���1��*���ٓ��(���)4�H>z�M8cq�pZ�ク���x\����P9j�J���^��ű���6m	��`_Żh0o�����﹌������y�G����W����(������ߑ��\oO���D*����v�- �4��tG/ǐAo��*B"E���(J��\����X�J@�e9�w��kB	Ib��.�@C<+0��E���L�� Y