��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��CN�M��rY���k�d��%�����]1�d	a?���u�P�e�q{�;&nĲR�OL�D��M��:O!����߸���:�6���R���{=I�9`�DW��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�I��U���B��<s���f\�-d�o꜓��
5����u�9���_=�����C8���M'�py�tT���)9���q��V4T$��G�CW���5�` Ă־�7�}L�P��$�����8��
&����w÷��AXR������3t�c#��@>���:Ј=1� ��|���U#�tjH�k}�Ҝ�s^��H�.�îƆ��}	
�ZD5�2�xd�����bv��֡�g���؉����=�<	_E$D�NLTi�@�涜~GX����e]�1����C�1�>ﹴ����#�n�v!�Z14�遅t,�S��sH::�g��AjR�p{�lH$V� ����o�>a��Z��nH��'^8o�<�����^�B�i�9f��'O�uV�h� cN^ƜC��Q�-�[c�.�j4Vg�šB�B)���+�-���؇��J�Z��(�g�t� ��Ѭ3�b8B���e����gS�4\O�c���Oz�$M*�����<}��W��c/�8ɐ7���Y�ۭf=|đŷq�D+�/��vA+�պ+Y�>nd���|б���������F�%�dYl,�u����d0QG��s��`�,��� 'E9�8���,D9���3^�Pp�G~j�'�H�� n��_��w>��r�i��V@�b�d�sǐ>&Ѡu���:���N�V���E��6mz$Y�e���S�M�<n�-��"�����vǠ�vi��"��iP!L.Q�ܖXmz�x�\c%#��h��/h<k�eM����\�G��RR�Ut/X9m�`@O�u�uG�<��mJEo準��E܃-� ֲ�pL?�kQ��|�3�ƴv<T�Y�ܱڽg��%�� �5��Y�)��W�|����+��[�w���)Z|l���}fy��G��d�81��������E�t�{:���<֘���|�yQ���Ɛ���{�['�f�1�|·��h�����5���߀aZs���qF��!U���7��K91��&�+w� ����;tx�u(�z��݁H�8fK�kx87�;�YFߔ:zs����b�^��
 U]Ol&)���&�JHATv�Y��A��{l.�ln��z�d�����۩��|��Wײ��R���D}'��w$x�frد��%ow�@�iԕӶ�LM���VS���p��ܮ���6>6g��K	m���ɔ�L�q�ߥ�����8G*��)j�U��oLɔ#�!�f1/��R4qO�u�����R#-�iM9�n=��ZZ�N���㬺��J`���S=L1]����/�K����+E��͖}5����z�$�g�9�h���Z\]��g9��~t�J��s��؉51���
�l�xW���s�W��MM۵B8�Ɯ�X��^INTmL�ԟ�;2��i��Q�Z��<[$Qz�&��۸���]c�i�W��-��\���>�O�!"��\���y%w��c��d�6����-8��R���b���l�JYT$��L��~n!��	$l���
w=����=�x����pߺ�G�a{����=ɝ����� 1w��K��t�Q�oXSn/J%�=b(� V7By%F�E�SE}�<��?�Dq�M�N\��f��W~x�uj��-�U�!��	;�� j����y[V9٤�o\��-�C����t�iqJ�Eu�8�O=�ƶ���h�?U K.G��9�	Q2ι��x��w����0�#<W�	8���|W&R���Ob����u/�L�T1��GwEdQ1nXh�#PMN�:�"�2�"�ԭq�RI�n]�MP���մ�&���$����r�i���z�1����J�	q&��p\�.H�.���/����_��i�%���[E����PS��ZZl���7R�&�;	��+a6�u�U��enY����c��HW�/v6��U����,�b���#,(y��J�߸����7%R��h$��SUx$t��S��^��0^��������T��4��./����KQ͘��T�5���'/x��l��t;l��5Ȳ|R�t�s\(i��J�q��=��JQ1�h߫(�, �b�J�<6�G��g�c��1�]y�Y�ao��/�?��(���YOj�t�9<�0�l�k	�����c�ĔM��Auan��!ӑ�����p�3�M�*9��s\%���f]��I�#?�Q���<O7��0�j�:$<���J�������T�%�d�P���o�P�����O] ~2�z[���N����y]T��b��[f?��FlB<vFzVá���o1�#]�0�8j��dl8���-�"�aԝ ��'�A���cwT?�����S�p���ǛW{�eN�"G��b�0�Ug�� �;K���;������@{A�-Pa��-HŪ�_d�F�nd{{�e�[2�ݾ�����n��3���[
E)��%qĺ�d�/X��ȅ��j4<G�2H
�� Li�黊�I�2 ���B㎄��AA��I`)��]k��Z�����E��ͻ���h������"�E���6���V\��F��F�y���৑ F��vo����a��}�,��1���Kl ���K�����fv��f5� N *[)�ި)-�.h<�s���E�l���T��EWf�`	D{t�ʴ�݋MX7����
�o�6���Rτ6��\�}h����c9�g��q|Q��.��ND�?f�"�x{��%w�9�\��K������GA�C��a�l)���h�JG^������]��wo�Οv�"u�I�����'�T[1��J��i���<=�����gw+D�ŖfU����M
ۈ#�Y���r�b���e�x���w,}׭�p<5�T�P����y~��2&�~�o=b}u jآ�ڻZ �UVO`�1��l��y2�F� H�:��
]�ߡҟs:j�#â�;�T1�	��yQ�>c�&�{��K�Ы�Ŕr,4�
fs8����5Wi `9��_���;���2ġ��Ɂ�c�t��q�듒mXa��lW�C�,T~����0b��d~�ϐ����*#�1-ŧ�]!VlJf"�Pev6So~V`9\rJ���";�����	���`>�Y-���:�!^�".:��x�,|���-Y��G-,�z�Yp���|7GI��_��Ɠ��i�$����0i�J8ʀ�}Ή{9��.k�m`�&��] qx�H�S��]E_hI��	)I1Uq<����A��T�� s#�����~��Lp�e�צw�x�n�F$|$bmA��YcĤ���_FhhɊ�t������_W-�v��	���E�ш���[W�:-B^�~gu
���,Y���W�\x��vab��k�JL���k��������S�
�[t.�1F��+���
{L�u��_2Q��Ŷ��T+������xs�r���C�E�ZIB=�螅
�h�F*g�`ґj�v^}��Ϛ,Ov���]K�L����'41ic��1h������Ac�S���2J�C�O�h��2v����T�j@e9��Q̴l��bp�������]����e�0�a�~�4�܉]#���㒥+�i������c�M ��߿Z�-wn��A�}�F��P���ҩ���3__���8肴,ҒIKP��x��Αz<�cq�ח���Yw^({Q��bDWI�~� ��|{`'�-��`}wZ:���epo���8Xd�I�oI�Dp�
����?zr�����9�A6@�( ��Q_1��?t�D2��Rʹ2�j���������!���W"B)������z�sM&��B.�Bf�%�rC�W+'n�g�i������'�т���>S_ɮ;?(��xƸOj�3^3� �dܔI�/@i|g͑���ihtJ�6=��lY��Ӕ?���/�:�RK���]��Q����:�T~{ �?XO��,Ct�-A�׈.����e\ZD���>jPPܿ`���Y���Z��J��X^�*q6�W�v�37��c&hC�w8%�{�L�U~���bs'2��n8�;�ߕ���o�������|�5��\�i4y�e�Bc�s����)w��Q	�(�J�@�j�� #�;f5���q6�Y�V>q�B��i�&��s�z\E\E�wNeh�^ݠ#�����i�s>����Wձ7#/O�?"��(����gֵ���Dς���2<����<r��"_��Iddk�!����+�)�>�(��TWx�ȑ���W���7��G�:J��*�'&S�xR�I(K���u!l�D�Tp�9�"{$ބzF��^�pJ$�)B.;t)f��Ã*s-g	{:�X�@ĕ�ψJo�Kc W{�\�p�kHE�o��� yCx��mQ\E+�
����s�'�eKg`d�z�[k�V��+�)��a��:k�rn�n�.�n��a��Y����3����9��MM�k���"~筋T��: %i�'���o�-����:D���gZ��:e��s��;D!��T��X㳇��6�չ�g�_�d�^?�t� ��5�,�a?�q�'�� Mh��8�[7�����6�M52�M���{�h��,��2�*u���Zm�| �˃0�;U.l��[MK�{���fϋ�� ��G�F�O)��
�xc
����ѹ&�M)��&��Y�V�e��x�;�'�D��Z��-3�"-�ґ?aa��ڑ�8����.,/�K�����7�4�:�ܦ׵���n'�)����=�yLc���H}#m�GJ�+�Ih��'#�/Z�)� u_�"��ra}���#V���G�F�V��I����d���g��BKt�����rL�A�%uܚ��P�?�4�S0	ԍܬ�|�,Qz����T���Ro�n. T�("�i��H��:����oo���:��Y��ܠ7�0�?�oY�֧T�s�+/��o#�R�x����Xh���0�� 2�ܫOI����<�7�TӎS����֕���H؏2���i��2�n��>O��u���Tw���Ճ�y���(�����Acc~$��Fpr�J]O�1|p� f��C%sI��m-
0S���|��^��cql��/�D/@��d��ٿc�>��G#���*H��~��Q�v=CX�g�� |��D�: w^_	я����)H(��4�sxu�=H	��:�ooc'w�]^�!fo��^q��Txu�[��r +�Qjr������Y4�Y�i� KyW^n�p��ñ$E$Q������Qa���3�`�L���Y��_Q�.^�#�޼��8��3��=,���F�A�����>	�M��\�>�y�>dT�9��%w\R�#��OvD���ԧ�G��	y�P��h���Q(����z�0�dF��S��B�8{a
�$���X��6ɲ�s���Z��ՅGkE��ld��S9|���+��Ԙ�T�vNƑHN�h#��T�[Es�o~E�K�H�����];pR�~o5Ώ?��!�ձlX����yۏ�G�lD�A�o�M�U�*�Qx뺳�x�0��xdE�&�=q
��,�%�ضA�nu����t?u��E�KlH3ќ�a�4���b�v1&໔ۡ-��ȅ�ձϡ��{'ry͠B���%��ձa�R "�D\5�fld�A��4���8��ȓ[VPn��V],�
�,�͖���Sw��Mv�]��P����Lw#5��U���j�?�Δ�+���T+�+9�|�t ��m��&��:jː�g>_�񳖯]q{D�H����P���S�cn�Cp�E���[�B],r(��P0[&iIgZ^HR��I��a�;�}w]>c�%Ըt0ݹi�I_��#�p��*]���6�i����/�z��~���v����y���xڔ��#��'+z�	�Rt��]�¤k��r���� ��q%b�E��l�YaDQ��5 =O��Qm�9�1M��AZ�ӵ�i�d�������_�,����nz��"�|�D'�g�nM��}�'�˜ ��%;G�� �s ��<���K��D���0�����Bj(cr�3!ɑ
?O*t��Ef<<؜����'C �"�����>�A�tp�&'n��A�m�����d)��壮����;-\E͠�1�:i����E��E�w.;�;.Y܈�Ę���b��TJm# TW�)�^��zt	�f1��=��v�͘��4�����,���P�*!p����#if��������2!��M�&��W!媔o$O)��ow)��l��z�þ5h�вѕ�̛R�_�&��|���SM7ӵ1��%j8^�>�f@��I���n��� pN�mg�u���(��=��m&4
���ʢW��':����*u/�Y��9r+-��Tہ�����?X���|(t�i�ہ�Ok����
9�Mf��PC����e ��_�p��D��
����M����oj�{��Wo�������|�� V�g	G������N��$$�5~|X�JT�>�N�V-����&p]͝(N��M����?�G?F,�,7�s��[��B��վ.����I��� �Ӯb�b�r#�ޢ[9�>�nE,��U��`�����L�7xA�v�S̼E�?/���3�h�W��R���S�O
����o�.f$��T^n��,�1���U���ڳ���0�³ɯ��Ui�\ӹF��cڭY�x�fO��A���6�8o��Ϥ���Rj{��бS /�^�w�����T�3�pp�i�0E���D��45(�.洕�t�kw�lg�O|e�^,���Y$�!:��/Rn��wϜ�
��KZ�K2��)۪D���>����I*�V�c�\�\��b�(��1�cY�B|ynbǢ���1��#�K��a�b�&l$��I�{ьCM������*�7D�sRA���	hܜ��AcI��juzr\=si�9Xu	��k�kM ����v�	�p���4�KFRA��}%Տ�@�Oy���,�c�Qd195=�dE��@;
�9%�kfT�-��/���Γ��4Yr��Y���9���k�g9���S��HX�����?��4�@�w��r.����C.-�f��t�
!fY@�1�u%�vD�~G��m����ःдj𢈶��6�|��A��A�]�Q́�-���b�k���)�e��Mm�k #�g��b��<�YRXrʯ>�C��R��*'i����v.	�*���)�$�כ�!_�l�c��<�4CI|O�z.�z���RT�w��T�������2��g��Su^4!8x����wDi�oK��{��~��}�쒬Vwtլ��?��\�2ʡ��\���9f�8���S7�5`��,��ȴ[���u���`W�~�L�	b��PyȖO9�2��|yY�KB���$����o��\^�xGC�����w�wyZ��w�t�{���;�kfE�`�T�`�}^
�لB�����}��-y�����G��O�1�Vtҭ��E*lw��-Ș�g0�k{��@#�lr���FE`%^E�<��&��):�F�M	��u����a�ߔ���I�M���g��cr�'�mF�r�f|Y��x[����`B��m+*~�Y�3�?:9�\��h>��j�E�0�U1ک���X�~ٓ6'�sNp����'��[dֺd�{0+��L�V�;<LH��'��.��e���W�G��oNv�T�T��e���>���索L���|4[_��)lӹ��MeLCMl�F�Q:}���@RW�� �f��ƌ�:E���7��V���{�����ʿ��s�	�΁��-�9$hjeޠx���}���^�.+p�~��d%�텰���W���<e��7z�Bf�O+~ٹ�g�ݏ��T���慠ȕǍ�f̯%�� 
ϙc:�K,p�hnUV+�;�y�=I�����h3�%��̑tqh�q��2�s�!
A�w���a ��;���)�u���gQ�_����6N����{���@����-+!�.��sP���b�闆t6����&��d������I:�X��`̟�?]k���	�Y�4�Y2[���0B6-�I�:�Y�b��od�RƹЈ�R`}G�Cճ�tgx�l/����@ց����xR���d�kfQ߅�*���H�`j�ܚuCe�@�/�K�-KY��-א]\���ۼ�9�9�ʊ2~���n��1�m���ڼ�����������g�P�Y��LHZ������F�y,���uP�f0 2n��! �,�x��d�ORc
���vcE�8s[��M��$�s!�v��%�:��D������a�-���볯�8q�ȶ��(�W�X*UR3���հgϢ��GO.�5[���:e�ߪ�{Pf��SL�[I�i<e+?�r�7����a/����C �9*�p�Ϻ[��4{�VN{���P��ҙ�UY5��_�h T�n9B!ˤP��么~얯o�`)���nj3���yf�yn��� ,[��+F8\�'���L�\BMa
��M;��Pitõ��򐰿�#l)��=�ecȫMPP/{Ż/�s�?ԃ4(y�5"���sOw�<@VG��>�ܟ�a�2X�&6ߛ`�o5Ҍ)�a�R,8�m).!���WJ�j��YzNUS�i`�6��G��l��,�פ:�ք+�w�:fh�����nq��ܬ��jU6x(�&���)�8(��O�J�2�(� IdhSɎA�+M�n�s���(~�CQ�^Vt�Cٺ9ML�2����2Y�<@���l����Y�1Z*=�`5�jݐ�n���'��!�bIë>����,����X�{\t���,A����ͼNH2����Q}m�`����/]��=�< �3��J�Sk]yV� R� /"�r��Op�j_���TJQ�b<���<"w�}��K��%���7��Z��nBZ�&�st2V.ܹ�e�$���F�vz�|o�4�'59H,j�&%�]���h��FZ�#�X��À������p�Uf?j���.õ.�Mec�듿��M�~���6����SUEf�,Ʉ�O(��Q�+�B��g�����=U�< F�:�#"��_��H(��/�N�<�D<y��5Mq6�\X4c���\@�=�����0��U5ůU�w�OB�rj�wʦ��{~���v-��Jǣ>����n��R�s6Xu���1w��o�L4{�4�'g��DH6�R�%��wQ�99!4���`����߽���V���*�3���ĥ�V <Z����G3�ݱ+�"\Km��Zن�|@��$4`�3���Hv�8���S.T��uL��ɠ�_�P�<�!dJ�ٯF'����-����%ςs^X�B�A�W���Ī��� 4G_��(Q[���+��j	�f˜��ib�@5^Zw��Z T�`�,��[&��!��P�2�7Mꆶd���#��?�+�ǰy��2fۦ���Ք¨��u;�'�b8khg���D�����&�!,|�	�Y��>�����:�>;eY<�mc0�h�'`�O�� Ӿ���F�\͕�/�t�Γ���7�?�t��[����E���Cok�^����G�$�d"�oš�D,v���>���©Ӓ7��k�TP�`bD)��x��&̇Uz,B�v�עr�C ���S����}��Cs��-�r��ԯ��cS��DA�,w�wQT/�5ȅw#����Ln���ݙ}Tv���$������x�V?@͈\XN��΅IYa��Wf�^z�NFA�[�6ϦG�KG�P���08�+붪��vVdwMt1�̈́WL)0�"jx~2��SYn�8��&�3S�cm�)�[���N�$�	.b#;N;@PZ`��9���z����n3$
�����Y��x}�][��]�_�r���
��3Kx�t���>$ �L�e���-�.]�Z�{$��Z%��Y)-�˾�\@h�?(@�������F<nU,Ę{6!�&�f�ML�,Ω1~�3_�%��C�pb��Мy	�Y���o�+fCG7X'މ�&���r�9KW�������T\��R�Vp" ���)P�I����FI�]����
�X`�0L51鮥�~��Z�����s�#M��K�pك��9��%J��9T��Z�h��v��X貵���c��ݡ�9>D [Y���^���Z|Q�(5�ń�����H�+z�|w��-�mH<�et���� |�H��#z#ᷮ�<+�A�#X��g�
��EF����V����S]��k���EMn�l���N�X�ݴ7�'Ff�~��(��bM���L�0қ}g�Y�_N{D:��e.�6I�Sh����Y�x҈����bǻF7��j�켉Q�������P:Z�.�Z��ؒF�#�Z_�~n�3�����+�U�s��aM:��X�G�Wz��Ş��+	��������o_� �����e2��o�:�zz/5,�x�n.uٛ�ϭ����t��D�O�7��W##���A!79��Xd��tiވ��S\Q�}���^ӯ��$X٠��k�;��:y�2�벶����������%2K����P��)�R�8���ڪg�D�G�`~���ی��e�6O�[�&f^�_�C��� <�UmHC���D�@���s�+Fl������l��-��ʵ��þ<�,ڨ1��Qͅ���	�P�4=db�$�*1�t�c�и!w݈{�es���^�3�7~�&��m�6��QbcH��[��'�7�Q#������)�:�R�[��j,�V�w{L���U�t��i��S�s�V^�M�L�1�l[tJ��Sj�3�k������T�ۨ��l��Lۛ�����p���%�F�Ƞ\�a=]g��.��p�C;
L?/+O��ZC����Sַ���H�̠��Pv{�f��6��g��}3;+G*�#���
�F���1V�K�˅␵Wi��xw��H�9���G$C�&��z�0��$��I㏈�A.`戟��h�CʤQE�'ӆ]'��S���(PC�/cԐEC�殠�F���0W�ܭ��J;b�������Unww.�;�Yε�ߠ�����,��>q[�䜍��NiL����nj�OQ[��z���u�cZg��f+�T,�M��(����Û^T�1�:�㯩�;n�/9�."StqZ����g�D>��~؏�<�l�;˙�é^(B��K���mi�-�����_�ᜆ��>8��e�.Cd�͗���b$�7��-o���:�!W�����$���J-J+x��Y�o�J��;whg��������|X�=h��|{��E� ��^z5C-$&�f���.��&:�wo�?���bM�KP.�@ S)� ����e�K^�܎�!r �xɬ��������$�R1r�Ti1��>y�*>�^�s%H���"�Pq��xf��*,�t�{�i ���px�wlG�_��
	p;#����u�7Tz%�$�Z!ۓ��+i��X_D*��r��Y�>��
0�A��M�kaP��S�ӗ�B6C._�#F	�C.LʫA�{���	���T,���׻U����/dj9�1W�v��]�+]5���DS��B��s��*vT��3�R�bR�ӡҼeo��P�����6�`��� w�w���Β&�lK���o��>�
��aj�/�����]z'���e�A��C��g�4��+���_����{h�a�:����֙b}��x��i����I� C'���G6S��h�o�גe	x�t�3���:J�{F�.��~X�����Ψ4X^'L�&������������|)�rl�pӀ�4`�b�����з-�gy�[�'=��
%�OzHS�L���E�!�X��Py9)�{V��Đ�j�B잢���F3$C4�$˅����?T��7�0� ���5�t��K������B�j���`f^ۜ����{Tu�s��Ʃ��8�Wa�@t�{~:ӝ��K��(p= 3����s8�i5�vU[��|ĵ�f\�ѝ89�J{�)X<q�G;h���n���ӊ�%ߘP9�TY���1/;�&�k���^�5���e���225�)I�4�B�,�� ���-LMU
HH�2\�#����`���V�E�{��f<��Fr0�\�ۗ���-�5M7��	*<�]��b�o�J�Y'�vXƺ|2�G���V�n��K�qx�E[@���K����H������G.+��A��D?ʎ�e���\#�
-�9�3	��_v�%d<�4�(�L�� ��:��%n���3�^�3,!�D�l����b�
�	�^m3���9rAC�Sp�e���_�}�� �JD	?3r��@��i�'w��`��ۮ~��SI�����H�vӃ5�G��dW���k@���u�H\cc��L�o`���K�b�՝��^O��4L�A2c�W��Y��g6_zU��D������'����5� ����'
���G|5�׀���Dr!(��@>Tz7����"�Ȥ�nUY.HXVh�H�|o���b�8�_X����H�ki��h�C�_�֙&�׏
U!���o.��@2iL���w�,�s�&^uťn`�ѻ�NBS��x��x"�(��fm[צ���D'�1�VZ���p�)��J�`Ta�d�U)��Q��]x�<�ݺ�@�J'3�u�F�-�	���4a���G�Cr��ޏ���-�X^"fĩ�믊��֍��J�{�ᦉ�M�u��������~'��xD����i�c�J���\��͓��ٺB	ɵ8q���̿�`x_�<�ҳ��1l��b�'�A�����3&�kySF�R����y�xS�Z�ȃ�h������W�����KZwo_�.����ɒ�
�s�ݾM218߹S��>�F���\Y��X6�|���}�xB�?X~|�@�z�#4(=����V{AKf�W�bD�"	��L/T�
�Ca�e�:еI�*	�$ݲ�ݪ��͕;��B��F����:��$�c�!�t�IX���R�=[&tļ�-�V��{&)�y��Kc�nQyސ�W,WHwbZ��-�ɰ>�u^Y����E�X^U�^�C�)QA��K<�=�	5��}�LnT�}�n񪿜�P_��IY���7\�=�jGM��n�����_�]~�1x������q<�{V������-�J�<=�(�Sh_jp�'���j��ƫ�ܞ���|���ûI�:�u���9�˖��8=�!~���e+?���yQ|H�[��lȌ�:��W�u��M�C��s\� :i��B�Ni���O����+,
��D���1����%�N �3�!�5"%�&շ����T��u�ZBԗ�dr�
�#"��|V�ol�R��ѩ�0����&��>lָ[o��o�<B�FN� ���m��J��������\�cQ�}���)�A�G!�Fh�P��^�URY��O�%S����q5�ח".�+���	R���no�"f��+��	Z*��Ú�|=�4"���c��8��n��w/��g^��A'8�5E�D��s����pw�P)0nEicHX#L�ɕ
�2�B����i�K���Ɓ����|  َV�")�F}
m����sϿ�#�)����}O9�W�����<��Dw g#@[A��ꎞ����d6�/ODK�%����/j%B���5�ݧ�A��!s���]`tn&$���"�;��caU�p�I%��4�Ŗ�!&x�M�H�2NX�k�>��봡	�:m�ç���^=��`����M�w�f�0�a��G�7D��a���1�4�ʨ0�c*L��t~Z]>K�,�~)ņ�TuǪ�#�hi*QYU�(��?�V�E�(y���$�A���Bl��B�V�n�m����4|l�3�)
z'5S.i�XA��(k���|Yb?iz���}c�P�Y���BI�o��L��S����ӕ�Y�<d�S��Q��g3������%��ZR~�R�]+����Z��8+N����w��#�T���.�����Um��1�Q)y0�&�4gp��dm���zk#�%��qT����2���O�i�|M@ ����r�i�q3`q,��Z�g,о}��ZV�y���1�5r�`��_2*{���6�>υ�Mw��	i*>�6l-E ��H�,]D�7\���4]�8�>�HBI���X��+ S�~m;@e�\$�HJ��1o�Z�+S��^^o_�#�%PbΒ�R7��g�A�&�^DX�ϡa1�d��@A���*z�����C9��/��f�Ph���x�rh��a�
IT]J��Ն�ɾ��-�0����'Ԉ)?d��J�D���ϱj;L��\B{]��ۂ� �Sӗ�{�11���1&�E?ߑrf݌\<H.���A�:���b����+o<s�0������!���qCEY�����3µ^�>��Uk�ٱ��Ǘ^�I�%�+���`wcN���hfX��Μ_Ӱ�Vzʃ��`z�6���b.��?�W�|rA!�4��Y�6�O�����4���h�=��%[�Am̩�h�j$q՟��
[�Em��)��dd�|���1BYe.�Y[�G~gߜ��Ig~r����A�+�u@�U(K�D�:Ͳ�J~˚��T�B�0j+����Vɣ��Z$�
�R�'��b�_�4��[�۝z�\>|�ڗ:�-�*��f3oJ�P���>�J�G���%pإfQ.H�t+#F�W�|0D\�6h`-���S� �JJ�;G�VV��زA���L�U�L粿ـ�}���<"���%�ȍws�s���ܽK�x�n];�ep/���̘��	�6�ƌ���t�Ѽ�����C�O�PN%QN���G����]���F���Nd��fd�*G,G{D�)<}���r��0�-;QoS�c�#��E�d"��Em`À�Ss*vm'$��?�d�xjC$|#b���Ą/+�O���`��~~6TZ[pV(�p�ĕ��&�״!�r�g�=pW#k�_2�`�W���:��l�9k����4�C{��O��̜����~��U�\ֺs g��s)!ä���ቔ����K����٫_��݁X�s��]gm���4L;���動)j�R�$�ݯ���tq��S"?�@���P-���6����+��F|n�k��4����G�s�R�$���X4h�����1�nWJV؛���$��Ij�u���j��2<i0r?���h���e?u�������� #�E�W թ�����^�$��O�?�\������n�z��
%��\���<�2z7d�!�+��>�R;��W��U(��l���Ĝ2�#?Ů�>?��E�s���	�a��*��f��Jog����2ՌX�Vt�Sf�j��,�� #��h8(�V'�� ޜ�L��[��*|@�;9���^8���i�7��ጴ��Xm#��;5:��h{�����<��
yD�qT@󺓸��)t�W��׹�2��-�a�R���1ܷM����e"22����5D���}�T��Z6l�K���H���X
9��(�����'��F�T�M׊%Nց�!�W�ԫKf���t���n�ݥ>��� ,��<h��' �ʒ �d}�s�N?�D�	P��|$��)�+a���?�|؄�
K6`�&��~���A��[��۽k�$m�A��3*H#]_z0T�d�:��g�~\�K���]b���wY�6ɒk�ƌ�}� 𒜎��]���U6��)Ť;N�������C4�d4�soid�I��	���)cHq?�X<u��c���N��j�~��0�F	�x��O�& ԘXG8�W�6�RF2X�L��!��+�1����&u� ��)E����%%!w")k�O����58��A�~��>P��|,����lm�B��)����J��[�"+$ s��U��AU'{߂54�}���$�k�Bޓs�&��eEm-=\����o�jZ)�E8(5��A��
 �A�f��@Y�sL��U��\�C�M�@��ڲ,#�`���!�ˉ2�#wěB����/��GϾe���
 *z_�?��^�l� 0��'�i����$R� x�@yC��ʱJ�A�Wd�{���Z�ڬ�����ay$��0�M�i<DbS�� ��Ӄ-F̋�9碕ٮ���/�����8�2=@zO��+A��	�+�13�5�j$��]�V���TC�]�w
���(���:��֏2U2�$��:k��Fc���
WB���h�-����v�A%��pq��`���ѐ	>�廓���!��ߙ�q@_�R\�<l���H�qr(�.Z+��QmZiD�����F27˴U�����z��^�E����>�!�]�-Et�tE�g����p�6G��P���w�[Ngυc}Zwk�8f�����a��c<��r�p?�>�`�E%w�3��&�}$�{����mQ��Ku,��Zڇ�lz�f-hj�Z�[xڎ8p��C�xm!����T�b
�OҢv��/���gg-�����[�y`D�	�z��wcl~P�6��Q�A]��6�C��O�6�2i�k�^9��c�$�2?���@0�QT܍ #
	�vԈ�29�X��8��ob�&����������mL��A��?!�?v��T�!�v�$�E�`�Nn:�}#��\�q���ڷR#�Y��A�CE���
<1A���J�Ai�{�
X<M�$z��V}�k�qL����Kf᠛�au7s��\jkI���F.�m�yO��w��j����P�h�E/W����G�knP��y�YU��a�LT�(���\?�4����{j��L8^�����������Ȭ�����S%��=�7�*���黄�`��Lcij���;L��4�0`�5�'�ڳt3���9M6&ȗQ���:\"��*�7�f���t/,[����2�	�\a��T�_;�%0_W�Zoa:6�>��v�9a����<�������t�p��BDw`�v{��C� )ij�4�X���?{�:�z����yo�E��2�1If38꣣��:������F6܋��2Xh�f��d�-�X�Ɗժw��3�Q��D����Q�Ö�ۧ15�,��_�.����0��x&���d���J'5�����?t>�a-��_��^16���T���b줤��o��%����^�q2]��@B.w��l@�I�� <���h2�]����`�V{���Od�V��F������)���Щ�H�1tT¯r��:�FM)����z'���
m�n�_'�u�ig���w7�q�l_ߴ�ڴ6��ƙ��h4h�v�.�&�&F	�߻ix�$S�zZ�����	�����d)�-xXE$�`�h��2�Q��轫,Y���=*eH��� >k���`��?<zg�e���OG9x.���*���/S�`pٮb���_��������[���k�i�����GU�h�����i��=Y�~n���v���+�\=��#0J�C�����W���ȅ�D����PI����іEBR	 �X)�j�T���nC����/�����0!��P��}���Ӑ+��`V��+�����n�fQ���� ���PY�l�Z(�[�}���k��rl�U���g�l^%Ә5���̧]�m6��L�Lځ�J�/�Ajt�,y~��e֑�	:L�	h�����M���g�Ÿ$-�/��!��r�T�F'��[��PT��x����/�t"�l5^�A�=�<���tȊ�;��LR1ϴV.�L�i�!�duj�����~U?�0>T�*O?fV�U��$@\���׍���a�]�C��s�hR&Ą$���L '��p���L����v��z@�Z"S�_6;Cz�
�,H�i��DX�]��>߿w�c�I���8���HE
��ߘc<4��p�O_ВT�j��26�Q}W��s��e�ISQ�4�P(1~�y%]gu�sh셶�r�=>�{��h �t'_|4�W�{#s5��z��&����x��pq��v�F}��#����"h^v�	 ���e���5)�4�óyw�ffNbd�kF+s]��'`�Yy��_��E�n��Da�2�1�`���K:�J���i*���g4�<�&��ҧxA2�k��jLo�Lj����0W�����
Rx2�����V�sȰ-g�����r� lU�\�E��3�l�h%��t�^ Sh!3: ����DU�r8��P��%u�<��f�=iϠ��v뭩jI�A��m[� �ʁ2�8bPґ�e�b��p���f�48!2�C��9��!S}�KⷼM��^�8��/`B}Ȕ�����QL�:��1@k���0�	;\�A��y����G4)���T^"(U]��PӁ��W{ �#��+���u�xF����ܥ|�w�n��,:}��?���>Ԧ�D?ވ+#^w�B�fz���Ig�Zݞ��]���,;�:FD��?�1e/(�`�(�@�̉�����B�m?
�j0�
́���U
����+[�@����0��
�T):��|~$��KB�e`<u�c�%��Uj���r�d��6��9p.ÑD
�Q�z^>�5���rig2��c��`���C�Gv�]Ÿ��1�i��{�a��N&�O�"T$�*�X��N��hs�895�skW����8�- -�0{�y�伬O8}�ڿ8t�GTQ��x�y9��M<-Ψ%�)!�l�Z q����f��h���P�37���l��)���6(�oq�^bQ����h$��q=Q����tR�c�%p�M�ۆ��1GF,ע|%�d�ϕ�mc������Ll���7��f^Ӈ���}�S�p��<�i>6�hs�bZ�K��Ɲ_i�����l�J~���@�-=�������L�c�������-!�h�Z������>�����/tY%/2����p�{�*���N��4|��G�V�Sk��4�����_[���6k�aP�g��_׼+C5Fe:�����7�O���U;k�\�v�C#&��<Ub���b�D�޽<������:�t!�� �Cs	v�[섦,�N��~������ ��0�G���s� �}��L��T@��H�~6����ɕ���OgpL<`�>�lV��uNcO*��
D�GN���-�yӏ/��}�M1�.��N���6[�~��p����a"@���o�:l��u���Z��z%K���Pw����s<�.��4`����S�ԣ4�Ǫ�'HF����/y��y�C���b����a8)�2nJ�Ш�	En�\ZU�6s9��贩"=�o3���8��Qoج�P�Ɩps��>���DO��Xi���j"�W�-� *�3�ϝ}Ɇ���@�*�:�"s&���۰�nfAU�g���#�L
�[������j	�G.�����l�d_MM���h�d���ypvz��:U���^BQ�7x�D5k�솬�w=��1�]}~���K.��@o9"��888���l8n�Q�z���Û��7lF��ۇN���1:�J�� �n�I V�Y�\~��s��+|QO���X��k덣H����.d�_QIߋ�jIPc����31�S��`�6�Q�[R�����Z�{����v�h�)��x��δڟ*����1g��ހ�{~�ß������P�s�a�&�Yh�o�>O�ᆪg���[{ú ��yW�ع����LZh���	�'P���M�%��Gk�OH����b8t��Q*�8VmK���40�)%�PB�F7nq���$Ѳ�=il����_��r����BK��FC��P�_�)��bEE��=y�B�^��%z���9�;÷�b�+�H��O3rQg�u�U��E��u>� Y��y�]W�}����>;R�uq u(�|�ķq��9�6j�뿄?P㵏���퉦������CA�*��%��d���[[խ���� �T�@��a����YmU�>��Rj�ª�8��#�@h��so�R�����c�0{dr��ĎnA=�:����K���)R	���w�GD�?�ۧ���.-�y[��o���#jz��6;m�Θ�nz���Y,rq�(;�o7��P{��uW�z���	�@:L-q�\��Y�ퟲ�r�2�(Ű���}^qə�♀O�\Ӂ� W�;zZg֕�m��"|1c�p5�(D��DÚ�Hҷ:<hekz��袋dN �I� �B�pU��B ����X	���.Uo��SۻX�R�'# ����8�d��1�����R�u��.f�GE��4^�!=�B��ɇ���PH�bD锡����Lv6���S��!!����-��.^��vjf�vgtܵ�w�b����D�[�N�l�g�����4O��c�P���#PT��4����y��v�1I��ϧ��+��P�Y/�1��nŷr�d�N������n+i٬$iuVx7#*W�b��҈c�l�h��E� #[ܥy{�:g�mR�8��p�g�b�T�hs�W���nx�8M���b5 ��%+�;�H�jE�$x��1��1�/@<�F?H�#�~�S�X$�N	���K�ِU5^�R���A��ĉr)�-��o�U���*����TA��"�?�X��(Œ�^'ό���<9�(��Cbӭx���XwE;�3��)���(�;#*3��p�k���"�4�� ��S��o�P��E��p˚�[M6k��v�<)
U�K�]�y��Zf�7܋�*B�H���ل�@;���Q^Yx����ȇ0ԝ�܎Y�&&�D�P6�_w�����*� �vU��^z�t�'],�Pdl,?e��
�tBܟ���͛T�����C��i��+r��M�ä#� ���R�K5��&O���]��wh�9p0"�t�Ԫ3���Qօ��g��V3�������1�fU!β����~���r��t��eEw	����Q+V{��?��Q�^�5@�cg"�����7\o��I?������	��Ra.�^2R3;z��7<.��kQ{=�6�͟= ���%�R���ۍ���7,�T	�蒟���~�C�@���c����w������^pV��E?���Wt��tIJ���8�"���q���͚�n'��D���������$RWG��<_@���*���>��}˲��P��;@��?s���讻��T#rx��( $���52G���y&@���3���o���xO������:�J�x8#�.�=�I���һ�6B�� �^��s�GaA���H�?x�u<�܅y#̾$�L�LV���<�7ş��Y,��#J�x+�EĦNZ&>Iw�7j!z���*OB�3������o"�&����n�`:���r��6�����a�h=��ԗ3�+|r�[�j�L����t�72�P��m�?]U�5`�&�����z&Qjʝ6���ia��wC?%�ݱgg��Ɲ����j��.?q���M7V݋P�g��y�A��(�iI+N��1M�?H�'	{�	k��F��N�$��\��k~C�����o�<��`�3;���q���^w�O
�h�
����ehҮ���qp7M���U?�xY�/��zyj���IR�U�ij˲ք�<c!Y�Ȑ!y��a@vEuc!�i7�d>��޸~'>D������C���[Ha}-;��	��b%1�a@j��Dp�R��; �/,@uMeA����Ar/��dt�ԏ��ڑ�����e8lkW�O���n��:����W�H���{�.9*��)�Oe����>�d�9t�r���NϦ�@�<��]��,Y�<��Ӽڪ�hlق�otHRJY��[��N�W�J*�ѐ�x��&$2\�	�ݖ�zI�D6�"=M]�w������P�~?1teאz�'O����r��mϻ1��ҋ��&�#0iZ�h�p!���z%�x�&���r���85�U�"s@�۵�+��;�;��v~��9{=�z0f�ͽ��Up�Ѕ�*s�I��o��><��,���0t� �8�\uS�x�
�F���+Q��P����<�E�IT)�y�.N��/��A�
���|���C�9�Ρ�_Y��ǁ�;�kMR-=���.���`��ڏ����F�=���	an\+�`NF�C�D>I���&�i�Y�㓊���'��� X/�?���l�e���s_��cL�@����MBoz�Ju�CٷU~ѷd5�"}\��CfG�P�m���0�x�o�ѯ�8d��A�ǽf��Au��w�\Wj�M��������;٬�C���S��E���I%��d��/��)mbP7=i��b&�rʍ��� ��=1͘�OxCR~�zC4��m�����'~�x��f�R:T�->�#�:8����Ԡƶ�%
�z�}��:��{4�����+��:�T�7�7�u��Q��L�y�*$(IwOMY�uIZ�i��E�T#���?�y{�r�<4r6���s�$�)��dvRֽ����p�U<f8(#�pN�!��D�hk�u;�ڷ�>ܰwe����&�q�� ����F�k���5	c�yMv�@�� k��vE��h˶��-?Cr��e�O��E1��5�S�M|���.	�v^s�6A�*$^�mD��}nl���+�$F=��-�bpk���i�$gd��Gn!�%�)�jR*�=�2���[�Yl��M�-�,} �$������6Xq�yB,U�AՊp��<]��|��P�	�P�9TB���C!jg����&��sH��@�48�C��g8��5m*�Lnk��td�_p5��Tӥ�� ��ٓ_2��]��y�$BI��']��sS@
����,��=9ص�%E6������k��+t�j*���Jk$E�J�ODx��f�@�\���**i�P<:~g�3�,�}@�f�Y�p:�F�J���h���Hva��2������p�T�����r��KM�,?ץ(���_khK�n��J�P1�>��B��N�3�u*�!Q8~��aM6I.�!w�Z�
�bD(Kp��8J��� Ѿm&Ip
8�����S��U
c�f�ҥ�a�c&�{��dVvd��]���d ��qy$۰��KA�2�����饜HH�H��$�Zn�t�=�iFy'\����"\���_7�54�l�TM;(}d�)�]~"[��!�����4f6�=|-��̢�C�Jo<��������I�e��h�C'���p2�ӯ��X�V���"���+R>�^aT��B�6�^�Е�:|B){�W�6�J$LM��N�o��C� ���$|9���5�W��_�f]���OO��N�F�f���	q#.�.#��74��fu�/ų��t�R�̇�=._�q�䃐*H��I��9������,Y���\e^�@��F����2*c��U��p��6�X͍�@�[T�q�1ppɋ���{&�4��D�X����k k1A>v_;H�6XTR�{�B��k?�t
��$�)5>�ME�r��!��kXp����@ѫ3tg�S[�� x����"��>���&��+�	p��6�XK��^��݃�/Q!iE��rV�_�c��;��t�z�{�T��V���c_��NV|���G��;o�2Y�kH�+
<CS����_�=�21{}i:������8�Ů�����u)������J[/��1kxt뿉�#Q�c#(�Y���n�	�{Glձ)	fݘ�2�]:�G��z��ʱ�R�e�?�8U����F��R�kљ�Zg��j'���7���9��F�6�aBjQM5ҍ�~J��%�I|3苑O6�E���1 g��߿}΁W�]ٗ�>��N\�����? �����y6��K%;����~*|˥����i�H���� ��L)}I�t�CE!m@1..�@��w$��S�+X,7����t=&DHB��P7�F�-�N7K��봼�N�AE9K1��W��T�O��UG����u�k>��b��<W~[R��Ɖ��V���<�g_
�d{!�|m;�6wf����T��êS�d?Q��j��^�s:׬q&���鿵�!��0ڧ�~J�
?�C^�.����("ך��4L>��],��9~.%�8Sh'T��������)uc�:��I��-�D1�+� ͋IS���}�1U�p�������1\�.�m!O������E$�"��bċ�cF�ٶc�]���{���dv�Oz��@�S?�[�-�7�'�d|�D��ɄN7�G9�0�Z��uA�S��-A��	xQ$�}�n֙5	�����ִ��.�YW�-�%�|vbx����R���#>v���;��	�M�n{�PͮƼ,�HL�?
������w�Em-Ndd�S���Aʗ����|�2, ����C9�PKؙ27~kr'AmGW��K��X�R�T�y9���83?
!9��4q�U�	��s�n�eaN��W��H�6��5q-�'xv�$M��L&��9��I��4&�O�p�Lm����X��������k���أ�yv�4���i�F�`L�P���
��qeXp����ù�?U��!Na��Ȳ��3t��[Xf;�fM�KE#]�X�,������Z�!4"y�oϛ�����i��Kqs�՛���8�6�nz�G�V��_��2��u�Nwd)^�?1KY}YT#$mG �j7�8j{ �f��%�Y��(�c3��� �b�ZG�D�Ɣ�r�
	2�У��=�p�)�"Rd<��`3��7L��?�x�C�GV����m��7�Pj���%�M�vǊ��7������)??�]� �i���7�c|+�ͼ�����r�5.�[z�����8lC�L��_�B�H�L�m(~�/Z��{�qbMbt�&hq�Ȃ@�4����Ys�{ă�o�_3^E^ �ZZ�>���O��ES����t/�����L���Y����W9TF��lP���J~j��� &�P�por1�M���]^����/O���D��4
ľpB�fP���f�U-"o|@�k�����L��C:���ʧ��ݧN[Ӫ�����c�ī{���H
�7�LL���1�~�}pv�Z�_�^0�rD	{����}w?sBN��fhA��5�.�>����1��Vl����E�7
����U�po!3E�w��6�r�	tf;3Nn�"��bA��uχC3�H�l�%Ec��oRD$�4��T��+ �h���j H�������z����b���ø��j<�=�t(�E6<6V�d����Z�G`��e�n�<�Pq9)l�&�LP�颅��O����̥���F�H��;����rP�Q�Aӭ��&+o��*���,�`;��'�8q��\CX�%D.�A\�|z�g�e��.\�w-����[��Ae��BjHhŢ��xv��#��ߏS���=��TzЋ��^A�;e�	���r����B}5F��i*tN���k5B0��*��c��5��kZ`󺷊 hgKO����"���W.q�����`�͈���X�V>_�BVK
�)�x��Y'�_)���{-8�MCI�����8x\XgGӍʓ�m�~x��+��n}0Fc/_����\c���ښ?MJ�� m%O��RD�ډ�h���+�Q}[K�[�Fs�d��y����K��c�"T�
�>Ȼ�����f�Ш���_#�w"�4"�ɾ�ߌ���go��h�b_~ڴ:�`�o	�h�Y��ǰ��z��ˤ?����je����h�ylY�˶ ��p��:�����b?
k�NX�N�!r9E�!��[��#q �V�h6(��e��������b��Ⱦ&�� �?�k����c*�q�8.[�������%�E��
�/�`�{)r��jS0�[ݍ����L�R-��#�/`x��;� ƴS�!i�Bl*R�Iî��O���rX��ؾiH�a;��B�z�܋b))Ӥ���0"����
�Gj�$=m��H*�u��B�'D*)B��CUV�S�#av7 j��oM�_\�Ӹ�CX���|z5�oe
��F�Y] sG;��xQ�.t8O�0���Ҙ]	L��
|���H�q7��Ҁ��܅V�z��V�lܡ��M��bx�H�I�6���P���*[��<��C�k�"L��3r��y��������ȎW�nQ*v<�t�5i�M���ل���a�h�.�y�-��g@T��+~��]�i�+�Ԭ+�x<���1�z̊�߷�gh�Dn�ܺ����K���bd펕�����ؾ�n�<C�,���e��>�������5�Qy�W���-P��l�¾￢�҉4BV����4��PJ״��f"vib�A1���c̺;�q����#'\`̀gE� �T��auc���5Aӥ���hW�zό�Q�����J'�{@r��7�qrg
7.��!|-����+V���jsp3����C}UK���Znbf��TD\y�*��Y�!oLW��HC�^7R�`	A�s����迠�.]��&���|w��?Lڞ|��� 2o�r�b����x���y��*k���9��R�6�z�EΨ�[���5��`	��N���=���[���I����OH=�(��{�%�1�g륿r=Kyr8s,D+'uy���;��}��G���8�0���=�v��nU.(���XiA��ɯ���ª�~{�.�TW�I.nfȋhA����))�p	B)o�Q����}�C/u�LyAn#H���[������g�����G��ʮs���|��C�S�M�x맨���p
����t�%������ҫ�!�/ '=�2�c��,�Q�����Ljd�s�W(�70���h�3*��z!��Ws++s��� ,Q����PJ��>�T�/���<�]�h&n��R{e�vc���:
�l�+�y	��"���6$����Z�4�����]�S���~����bn�2�;����b{�,0A���T��*��$�ŋn�8��pBB�8�����y�8�ӏgG.���,^VU8j��p�������A�J�0I���1o3�t���"|(�ޭQ%O�F�'�D`0``i�$2��0qY;~�W>�&�G���1j�?Dn�9ˣۃ9�$R�;��;�千�r�!9n�;~�!�],�!ڄS�-��GVW~����VdGZkHܛ:�z-@k{�!k��A�p��!e��Q{�;�}�媍#���9�Ň��(���}n����K���V�L����H��!ܬ΄��UЫ^���e�cd$�_�"��v�Z�j� �Epȡ��
���H;Vi�XHW"�Έ�] Iw�������z�\g�3�%L�;�]�ZSZlHN's��DV%=��<�"2\��<���>�^��/���A^�"f9�=��x+�1� ]v<�T;'�� Lk$9�g/���D�rX�c$��x���2��$��Z�#�����i�s@�?�I�w�m@E����\�<72������A�p�4���c�w-�&Ʉ/}p�9����
'8��5�Ӡ}�ş?T���S�_jYL~����@��t��Ԥ?	O���V5�� �r3�r$\������K�2&F���9�a�o�Q��i�E�x&E/�e�xe�l�M�^�ç��0���0�/"�8�O���trE� Z����<m)g�v�n�K�xq|H~�s�G��qo+��@��Sʃ�S뿖�⭦�){���&v�V�����B�e����	��s(*�g�S;\��T�����E�iIK�o��J�S��*^w�At��z��R`&�x?�
V㌷ɋ�IS�h��wQ��c��M�xE3~,e�y���C1:-��jH�Nr���5*C|�"���\����Ǭ"����K��^���Do'��-��\�n�����+lv���̤�[G��n+6��C'����]E���]�m(��~N�z���x��6��-���3~��+D�u�N���0�<�Fĵ*n�KYq 8���X�f����y�Im�'@O1�=�m�#S�"'1�s�;{�q��Q��iM�
9�BG4���B�N:/��L�'=*�ڏ�+�&������_5y�i\k��IQ�i�>��"C��5o7i��~��Y�}XbQ��kVb��7�.	5rTCCX�~F4��Қ��-%ɋH����P��n8s�=uBX�H��2������`גBPhh{U�L:��ȥ�A�"��bJm�,�P8�}�<����#S{a>���:��q�ĳ�l�[�oH�a�+����(l)�\�yP����)��-�Є�ַN�A�Ї^L�id����@�)��u��s�Z@���F�UD/�APjR4W*��沯��s�����<S�2Nq���Wf®M��Lv��o�Ð�Wvm�-5ZE�ҾU���L!�sqٵ�e�}X8�v��:H1�e)��d +gr���Ǣ0~{��̣��1\���:��=i-����M;w���L����}{ơ���f�{֖��W�#{��8lH4aE1�� ��k]E��M��yS�}����������N-;� �	�>q�R�I��0�G��`]>���bC'�r�1�3��&R�s��e��4�=*ȹ�-�����]x�/n؉�� XCqvP��Z�"LQؾ�/�k.*rs��FЍ�7�����P@�u{:����)�j�N�2���������pG� ��U�f��>�@��>I�eX�ӠI���:"�+�0�5�& ^�t��G꾿�{�*j&��@�+"�f�3����RT;�����8a�� ��n�/�J�����Ȗ�k���4ũ*q��X�X63�!������`sk��ġg)�e�C5���\-8"��V�*�3)q�c~�)���O�
��䤱�d�U�J�i���?�����qjkA�DLSN�A�q�E��8$�U?�9:�j� QgXA����':O�_=�Ep!��䍶��$��^�@�}ɉ,��2/�y��� ����~ܦ�% �`�+�������O���,�ƍ��R� ��`�JZ,e��ud*=o82�������)�^"ŴQQ2FA�h�N���2�8U�@�w���e�RT����Zp!��Yf:�3=�9������eye�'�T���/�y��!���#�|�IQ������J]ܓ��B���䮰C&�}D�kMl�	ײͷ�8��{r�\	��	��>��^���,�B���$��sB)���¿��{����a>�6"��w�m�P����t$�AQ�nj��f'���Ǻg�����t�`�Zꄀ3J=���Z'�i��F*�1�ssP�t����
��%�u�`�K�?x�lX��5o@ĩ����W��e��aZc���+	6�T�����F�L1���Hʔ�'�Vvs����
�A�!+g.�|��a��rg��H�'C���@�x��9vw�n�9(���]����l����h�ES��>��w	�CŅ��C�!4���?�я8Z(�WG��f�]��C�&�p�!5�~r�;I�*��o΂��2K�l%�*u�t�L�W����~��3��l����Š�.@g�S���A�y��*����@�ce-�&W��L9oJM;�z��I��s��X�D�����\d]v�rn���v(���ßB�d�a����+Q]I�D����C��Hn�g��8R� �� u�aK-aB�)��}*�E�5̠��E����nԉ���+:f&鉤X�a�Ї�]tdWa|���ƍ/4�]q�e����G8v�~���燖�һ$˺�19�m���f�d���� /�tPo�A�ɡz��Z�-/�dFQN�.������V$��UK4��׵]s��AvJ*۩�E��J4�_���5��)	Q"�w @������u�_� N��4+fǭ�ޮ�DO��*�
w�ҡ?��zB�'2p���*5���0���2�㫎�������K��x� ��yt���p�� =��P��D�I��nc�4�)w�(�zM:L��,ئmO�Zl���¦N�	�ݟI��g�Rx������u2=�a
��]�+X�#�5��S������J�O��Y
�
"�bg��AP��_k�́�U�8�oEj8��d�BCl���N�Kf�Tyԥ,i17@�ԼŦ�q��t�\�>V6�L����*:��Lx���?#����D�i�+l�h�\C��=����&�����+���!��胍/�_��a^�XH-ҁ�ܔ~�$��Q$o��,��,W�������v����wO�pb��`y]�E�Uݝ�8f
p�Oʍ�s4a��*�
�D��HI�u���rU^Q��k�.i�c��~1z�>@����J�z��r��d$b�\��� G��q�0�Ќ2�6��gt����\���L|�]v.�;����"�Y/�y����hY�s��{�6&�#�O�`KV\P�B���tT�tn�KW��3�z=!���M�/*����
*��QLk��.�ip&@�_��!ߤ=Ҝ2�,a��&I���V���85�e�:Ա��m%2�g�	?����ii��E@`%1Ib�����@�='�+*|'[�Z_I؛-a]��A�������K��T�,9����4�/�H�i"��/t�T٨��n$���v�-���W����o�U�I���y'W���;��i�
�8ƺ�1�l%���l\����0sf+)E�ڱ��'Z�J��D����(d+�Z z�\�2�
��� �P��E��ʏ���8��K�.��` arF7�Af:�����W� �s��'��_5{��I�0H�G��W�9y��,ݚ���U���m�]#cʃ[0��-����5��u�:3_�yR$��*=>gh��JOk����7���HN|s ��T͘{
�|���⬽[Ä5�p
/�!]��H�WOŢ�Sה���5s.��Qty����*E����;�Z�u�&����Q��1��S+���d��EB7���|�<օh.z0㵁� o��ׄ�ٷ� iQ6LΑl�_*ENuq.�d�t�y�˦z�D�0�IP�7��L����ކm؀1]�N#e��l��g�������U�Y |b��*]͚Ǌ�����i ��L�����3C�T����O���	t˹��\�מ?�;���Sҭ�N��a��&>�'�Ú�b�[O70A����7����Qߋ���(��s�{F�o%��E����N���Ek��w0�}�;gea�L��_t�D�4^��dT�V�����"4��~I@@W�r#�y7�M{p�8�����w��|���?���Z�J�*��m��1�U�@k��?F-l��	>��ˇ&�'��Ca�poE�D*|��)l��vDI�iIF���ͧ�茐;*���U����Dm��^z��4�d-��;O���	}��b��r� 	{�l��͎�:β��J�6�d�"hԨEE�Gt���Zv�ۄ��UiE�'~i�r,��r�D9�<���U�����̲)}tY8K�fn!˳v�}0�*����*|е�X?^Ѐ]r>ʷB�O�[���{�2ȑ��'y��*�23�BUv�/g^gBT�Q�Q�O�(*��,�/4IY���g��/��={0�c���>���ɽ���9]��bvt�%�Ƿ�j*�Oa��k�w*G&���s��v!���%�@�&��%�w�u��0������N�.�4/
Z� FҐ��"�G2�),[]|���ӋC��ԕ����r�C����)��%�YgN��7k�x�kE�<��i��a��ňE�K��s8�������2S���K!o�p�ȋ"����m:��n���kd�<7���K��֡���8PD��P
��K��:;�c�c�A�p��daZ�(���v�?����48a����y;Z�\�$�E��F:��)c��zX~��:���qu�n.'�1'J��}���ҋ~"�(��7�<�w�&x�Ss}9�b��}��l^�|a!t���<4CpA� G�����0�����q�z�&�(��(u2в���`ϑT/62��LtS���qEn�/n�I.���<LQ��p��˾�}�,NK��2��q�����ŻRB�{Q�.�F��pH��'�o {"��{ᱩ�FTɥ�q�*�#�Q>y����)���DY��8��ŝq�"B x��`��	kN�P�~ ��M�Ê㛶1ᨨ�M�'��˘�uV�'�6��q�({#jb}�,(�0��'ml8�����Y �\sߑe�%K1��n��tŭm���-�"&ִrQ�j}A �_9'L�P�H�7�f���G�xM�n�uh��������y�0���;Ӭ~��a˺gT���?K�7&zx����� �bЫ��{e�`�rD_���"��?=�|��d��I&Φ�J�v�o���_���.<��� mU,4�P�.!H�XJ�w����a�8�<�xoB*��T����cz}u�ɇ�e���U���v�U���i�48�@GV9���&Y�g�oӗ;�W�-�m:,�M���W�5H��1����x4R2A�-4�ܬ�;!s_�������fGw3���7�E��&��X4V�*Ow�/$�[�:����h@p�����x5�]l�~�g�S^����B�r��3���U*�y�8��
"�?�[�_L�����ł��������8�u��c�X�↞����7�S��2�1U�bvŦ[���K��$������A�E��v�3�,�k�Cu�]�t�i�T�{#�!��E�'���Tڳ�õ�.�:�r�~�:&:'`9E���wd|��2]��얠�9t��9�A嵪�+��������?Amv;�- �x)��O���
B��Z۫o����Z��E5s3��D�K;Q��p�^)1�cl+�\�r�^��'���j�/L��@UҲ�����觥��f�;HcQRz+�O%g�8Ľ'��.�,3��`�yԳA6b{�Ћs����9�]�	�y�s1���1�.���;R�����ɘ��$��<o�y'[<D�jĝhp�4woqpQ4)��ߚ[�%�`6k!om',v��\��>0����>E���	;�Z�P�iIlU�3f�Ltc^��o?jo`N��z_�j9���TC�v3�m�t��^���YG�kg%5�E�{4tK/������Y�g=P��릨.�M�4 M�o�X��89�Ti����+|�x�콄8ڋ�N�3D�J��}�B���K�Y�������k�L13��4��DW/�Mr�:��t�x���B��cA��k�xbm�QQ'	�\M�������zx��/1�qC�aIh3C3����;d'���٠G6���i2ܙ��K�z�É��D����v!j�``6�,VǺ$�5��5�I��$W�s�l]���E��Mk�����n\�!���&_��x�{h�<�`F'x���hw)�{9@v QKL<���dnЪ��]��l�����F}�}�9�H^��ʉ #��"�}M_��')q(bLX_�u������� �����}��^Q_�E#���Ko�bdL�!͘��:FzŜ�C[$��2��[
��YlU�->(j��5:y�2"'�O�oW�L���ڻ4r(���-��I���������v����43�Y�����n)z����1Q���~����k��޳9A)�㘲[�QoU��wd\�W���ʋ�?T�2�Ag�
���4�6-��e�b��F�TR��$kA����?��:̯�_(�eV?�4�Ǫ/�[�koy������8;�phF ��w�`���#D/U�F琽�A���jr�/�)+�Z��㎥N�|+о�U� ���,ͤ�����%:s7w���}l� )gcg`>2ҍ^1� ��}r\�c��� %�%��V�f��^+��K奬�!f�M�;�����*<��Af*yY���^ ��nk"�3q��.��r������ �u�x(�Y�_;�����K��"}/<|r�ݰ��Bϵ*�c�y��� ��a�Z y�b ��@]Jk���@ң�27U�j*6��̋��<A�=$�in�2�ta�-��#d�chTH��'�iX*`+xuq�q�z?����W�)�f ���0��1�`���'�'��P�KQ�=��M͐ۨ�b?�6��$���lhx�}*��<�󡦥y�+{T��;��ar�4�?�z�t�MȲd�J�p�-E
ªq�1m���|�s֞� 3�5_��U�?��4��h ��,����|RYh1�ό�ZAt
&�j,6l�إLr�X� ��<��&�������Ŏ�ɷv"��pCǏ$�v�)���Di�9N]̑R�>K�y��B���c�z�
�Q��!�g!�'VPz#ڬZ�w ��V^{_1xwt�+�\�h~�ʛ1!��9��# Z?L;���/�f�M�:���Vέ\zhPHDꁱt���.�p+��$��S{�Հ��~� ����:�@g������X
��BS ���w�:�0�F�LC�v�I�&FJ�瓤:�s�\i��8�:}��rs��(���C������!+!v�� �[��$�'�#����y�CA ��~�8/^n�n1I�1+w����*#/��}���hsOS���MO^�U1@��F��Q�/����t�y��Z�*1ms
�r "�MI�w�S��k�X3���Ո
|��D.,�I�{��$r��I���RBm�l-}��-�Psxa����9j��Ɉ��+J�t�������O0-7d�c�Wa�-7��so��>��4l���ھ��P����Z}������|�2��5���6�,���J"�a�?���ǜ��B0�c���k��� 
��pƴ���-�|(
&E�g�g:U� ��'��KK������/��g)���C�
���u/��?�\
GN���e��֮� [�Ի��hÞ F�F4�F� Xz�R�I/��"
I*6�_�[�����>�GIT֬���#�������L�]�of�R";q�_Ь��G*S���	�b�9�r[BJ���k����kw�4 O���h�Άg��s���dZ~F{��H�>>s�\��F�Sxv#����{� �е��;���y�a���7��I�7��D^��}�4K�lEo���+9�M����}5�o�J^��~g��=��`�WH�堷��=��e�H:�����'��B��j7���ۘ2�t�k_K�U[��O�w���@�{61�Ve���tǜ��s�%'�Bł�A+����"}�����Էt�omIT|�$��6� ��f;�ؔd
5w��nx�H��.���\��[b��]�������{�?	���ۆF4�n9�9�%`�U�v�J����nY@���S��AM+M����:�B�^�ʿ��,S:E绋���$�:e���$Q����>e���x���?
����[��W	���V�L�C�j�q�2<I&����^�W�̀��/���4�:ه\eU�H��!B�%�|��w�:T�U�#P �%i��^Oj_�d�*<�U�_1�C��0̩�2�x@+e%SN9�����Eu��tVt��Hrc�n�Ġ"h>t:�7 ���Ux>>�%��D�h�_I4�����]S�R��I��^ɹۭ��h2L��W����n�)W��ϥ-�zQ�R�{��*�r���y�����$^�Mo�P.��������VU��cZ�6<���d���*�1�<q=G�A��Z�p]@�4���x�=P��d=`�`�H'Ś��1g� ����[������r�Iҽ��3!H��0u.u���f��
���pX��>P&DG^�v$���(��2-��e�Px���B�Wy!��In<�i����¯EI���U�,�V���#�0���{��6�Ph�(>��巜�׍?ig���e�i��~���}V4����u"�ܥNʲZ���V��5�MܞR{����l�T����B�|�\�j�FpKJP}$y�F}8�.�M�mǴ}����� �+eU��kq]���Lfw�>�, �(i�&|%s�3tC��RЏ\��sO�F�4�;�'��1'�S�@���K��A����[�x�T�i�(�e�{#�5@dc@�]�)q����L�z�D���=����b�H�0K�i��4�/�~z��l���TIAZ��\����G�}�e��(B��RuM�v`d�#=�[��#�e��o�L	Sr�;[���ʽb%�w��t-��q힐�`�E�*R� �8Ҥ*���h���7y�΂����pJ�s�W?��|�Ј�\N�>������ �I��2!�4F���gi�A���,sEVD��MFabFW;�7�O��Ͱ�\��|0��a=Q���L�;C&�x�����[[+(�(�O�++�* ����{NtD?��Mg�����%w�s���>�bTݖS��(��[5����A���x�\��t8B���v=��C�f��Ђ�1<7���-ӊs������!~K��h�g5>#QO??U/���w�x76�OZ˩��E�U8/aF]�0���3��C��=�#��,��r�^@J�8M��-��8??�x`�LC�>+��.V��{���U6�t�-?�'���狟`ZÆ��E�wZP�K��^=���3+����H���k�����.u��ك	���c!H�h��t�Z��f
�,��HD�-|�-g6�d�Dl�yzDg���\	���cL��G���.0v"��V�a�tc�κzR`��N�*D3O'4���]�`W�{C@6�,�Ē0ϖ�30*���,?'	�@��e�������a{��~_$/������13Ye��q<����L�i?*��R����#�>#_
����G���fm��7u�A�Q2d7(��5����/g��b,��&��[_ޔq�C����8+'�F�D�Q1Ծ�R/�)͌�KiYkr��4��4���R�Nm���_�����?�h:�k��}���Cd��x�dd�6p����D�e�R5J�D�sw�Ic�Eɀ?�s-%�%cw,d�w�<I`MRr�\���4�~����W��:�G1�����낻f'%4��~	��Dkevǫ�I7źS呖�=�����|!�Ks?%�����^�q�cN�����
���p��ȿq���Y�L;�ŀs��k��eM�ڨ�R9.�	+h]�v�a�0��^gW?Ôz퐋9��2V�$(=��^Ҷ�y�L�,� �_c,�ؤn��D������Dkec��,^}v[[���9Q���-ľyv��1�?#�q�O��7���V��g�~|�����R��!J��Ra����j|1mL���Ċ
��a��ᗟ&�,P<�ǂ4���ʎ�Y��c$��8w^<�V������O����?n�8�u�B��Uw�-�r
_�y��3���L�%�	�1H�U�LZ�}~��f��=h��n1� M�`�z<����֝���/�ꑍ������~��;�-�}�Qq���Vѫ�Z�x�u���p��mh �Z��i�kK��<����O�"$'�n�*�BY�ֲ��*�'S>$�9�+jz��F��/ BL�CO����$������m�(���ͪ���Lfh���A��9��!�I$���SzǊ����H���{�Dn���T"y��U�9�"n�)��Sw|�\[��c����0ؕ}���Xd����!��woq�<)�:g��5�� Ʀ�ҡ>��2ߠ� ����$ ������|�i�����#<�}&}��xy���oj�����"�7��:6W�Ӎ{*��dJ,�������/���ӕ]QO����p��?��\GǛ���@�Y��yӠB,ʝǱ}�!�I56"Ԩ��_؜@K�*ƉQ�ࢋ�雅�
w�"�\�sVW"�~�_U��y�����56*�����t�vx:T7�ϼ�+*\G�@F�� ��Q��o�b��������wB?o�M��&P�+�M��p{�J�Պ���w���s��?�9��{K���gv��m���贼Q>�U��`5���I�Y������Y�����y��`)��=�C"%b����p�l%Ë�hؚ���ysR��A���8��~��S� -��y���	FCI{���J2�$Ák���C��yk����dz?��nk㧳Q;��,h�8{�ǻ��7v�����b岷*�1ب%��5{��7��Bv����/��=KA�!d�~R�(�썗4ς�Aݧ	�H����m�x!��u����Rٗ��}�2z�ĦU�
�<~��O�Qh�^TP�Oڧ�v�5���YҔ�3ڐJh}j�(����l��)���<K�0�1�+�3�g1>mٮl�ʜ�Yhl�'1����W�B�8�JЪ|����X�q�7�m�~-�;��.����>]�"��=�s��T��E8�;��у�"�1 �?0���
Y��}mC�"��ݹ3&aA�pO�� ����4n7�H_�W� ���{H%C��n��1(�K�x�T5.���kp����(:�޽�+6�ޖ1i�ќ
��K�m¼��i�5�W�RFXl�+�H�x�'�2]���ŗ@��h���k���*
����Z���]�U����Ly�k?K�V��9�`�n�]�x���n�#��;�q��VJ�4E����G��ݪ�`��鲛���t�����#��f����M��hq�� ����`X3��_�߱56��� �2�E^�ӊ�*_u�OY���K�U��J. e���_n��d���9c���xs�+�y�y�c�����8X�:>��B*�@�}W)��?o�n�� %��KiIu1u��0��D�G���f��9��mN��BP�����uS�a=���\gA>Z�CZ����a��ַv*.oz�2C�oMޟ3���ƪK!�%��s_nh]ki���e/*�4�q��]b;e�*W2E�-��gy�I@sc��v�bTB�#/5"=�5��~��꽙ac�rS�����W�e�����S:��U�V��;�4���#/�/-E��kg�V�t˔����2���u���R��4�=f?aUȬE\>� =��<Lַ=->�o5&��UP��Q��Bwy��XO��A?O�hِ�?����O���d���ܺ]��{�U�M��s^D�J����� �F��*���b�~|�'�9�܈=P�v ����OV�0�&���G]�Y�<}i����{�㾢≮m?T�s9�l��b���=|�'�>�� �5���C.8�a��@�?�����v��	�y�
MFt
6���;��8m[%��&6�N���/d��r�W=��p�
�ys�=���b�,7�^���e��z�2���2%2n��� C��x��vBN0$��-X�i	d��^}:ʶ�����OI�դظ��(�uI�Zw�G�9��+!<F���Y�����%����ѝ}���i�ދ쎖���0���s�e"�Y��A�|E��,.�S�0�%�q���~�_�`��jl�@+. U�^̵S͟6�g�(��y�dΛ*�K�
]�u���%��%�}O�����܂���X_�X�`��x_����|�KG$��~󐺐1��=�%�U�����}��;v�=�StD�꓿��cd	:�xKx��z�C(�����&l��9�$ͺ�]	/4n����VjPx�d��ɠy���iAL+���R)� �X6��>�|�\���P2@\Nu~H/�$���ϧn!^(���� �L�W��Hb�jr�זq9�!?W�2�6Q�o�k8��� ��)�xj��F���P>�n����I�I�X�ߑ-{r���7�A��b�5y3_��r�%DߘOR鑃��j	� �;1�e�-��jz��]u�V��H��s;�oG�
��+| �Ҁ���M�}��3,��1_��wSjh��t��V� <����W��e}�u�Zȟ �������0��ԘkR����`�~��ф}D���Lk2­�O���� Tz-)3�۷��v���b���>��U�Y���{�8�9/���������G��
�*^��喸g4� AU-�Z���揚�G(\���z��E}�(M�T숞��H6��!� m��5���\B?�/V��>;ԯ�4]��M�u$8�%�f�J�~ kR��gB!�MwP�N����g�۩�v��p�;#8�UH�TA1`���N�q���S���kN�E ��%N8����_��.l��<M��p�tV��D'{��M�=�*]sr�ȵ����k&�  h�5	�-]c�T'�o�*qJI�]c��6$�C�J�7�r^y�c$��pl���u��{�y�����O����6s��=��1%��xy�~|���(^�l��lLј(�ߤw9c�Y�b�IQ��qǺ��<C��AE�
(A�1A+��@QrX�W��eG������0��2x�W���f��~E]�C�5Tؘ�;z*,�mn�I#~�q�nP�|�ź�q����ET�E��Q��u�e\��#Q��6�\��^B����۹�8<4�w�Y@;L=
�	�d.Drc���S��Y�G�\n%��1�w�kY?���墇Ւ��5D6��҇��J@[��8&]���(Y-\R�z�����u؎��p%�D*����d�i;E�MCU5+%��"��j��-�-9a�p�����{�?K5u�,\�����P�q����p�#��C���w���tp�
��1�Yzd���i>��c�cK	��v�ff��b���0��=�w����9�̌M��N����mP\�D�����"�{��rdvh�Њ\�iӂ���,� }��/��ij8�@����_��ϓ���^��=K;�LYK��lv���kpʹb��t�ۙ���rO&�/S����j�� 4��ĪA�4��z��j����:3J�:�V�yb�K��h��]�����O��ɒ��.;�^48�f5tSm��Vva��A�Z����=p����\Ϲ�>�_&ʅ��d��K&�O0��>��iK���V{Z���E:�L�<Y�@�7a�r��&�!M�ita`���#��eD����C?��a�ދJ����3pW�zt���2���O�w%�� zw��$�E��@l�bM������1�T+R��\b��ЕC
c�#6�L�$� 1�9��αd�~>��9�����p�a;/���S��v��9���Euq���_�k���Ip7g'�S����5a$�t��'�uQ��VV�pȎ�	4D0�W3d��e�>�W�p߆@(C�k���6Z�~��\�UW�n����aO׿h������1�z\B	�DW�q��w'�a@���-E~��b��.O���*��UMEIs�Kro����s��=�Q�*vSH����M+�a�Jd����T$�/G�p�h\Bv,!u+';evu ��)�s>�?E��_<gy1���5�3�5ҟE0<!����\�h�>R�c�E�/Xd���Yj�>:�L���26�0�6�p�C��3�Y�#S"\6��#(<Eo�r}��z�l֟��׽gp��)q^eð���e�Mp�w���U�������K��)�T���2����nښ��k��L!g���	Y�4[��p�b��U�<Rda9Kl���@7���\��VEa�l�ib�������+1`h��­6/I�.(�~z6���K�n�*�j}�Jy�B}z�\^c�O�z�6.�y��$m��me��B�K����H�e�2��ek@%~� ܊Q�(�@yCj{�1���M���1�$�����}��`xP�c@Ԥ�i��H��~��%�H���P����=O�)�ƕ-��9�	Ȇ�򚹵�����Gu7�>% ��	B�&��z��%��c1���y�aMhu���cJ���)��.$J��e�0s��jK����i�#�8�r]"�9�����#�l`�-���жo1��O����w�Q�s4 ���#�x�f�r�I�1�A<ᅄ�<9�W�~�ͫ�7]�W	�p��3c_���G\F\p>�?}G(!!���{�F�L�Y�ͻ�w�����A�s���`"�F�-b�x���jC���W����&�f�m^E�{+��/H&�3%�D\��P����M4�u��0α���uw)��:��{�!��bt�˽���l�"���*�����~�v��x\��k4�_,Md�M��Bf;EqkF����jc2(���S�����bd�y|"Փ�:����ܧMT7S����#/8<	9\��������$E��iÒvo�G!���.s�T[��rCaT��:�S�W��%x��^V������f��j�b�o3��&��'��c[}�J[��ܱ���I��˷��':<���T�s\�ƌ�.�nT�'��uۯ�Eh���$B?9�}0(q��a����c�@h���?Lo�jxV��Dz�$�[q��.�
�N�yD`�}sU��T�	���a�^ug�6d2t��.CQ�)܌q�pt�B�%W�$�o��S�U�s���|��3�Iyr$0�ǄG��_�=*+�V�V����6�c���D����Np�_%&�FELw��7��$�����9�{*�@�_�ר��*�s����^X{��7�DzP�&����No�~��9����^�Ut�J+� 缓�8�ŞA�!F/�	�Q�@�0*`���"����RA��J�;��{u�A���A�����O%��D�G��ٶ2��x>����o��L�e�2f{D��h�cPK(3��<�H��S�a{�P��b�򌡳���A�Y=Q_���dW�<nm*\�F�q�M�"/�&׉s)��%ײ�~�o��0
���@%�Q�ӌ5�趜�!"�܅�2R`��,�	P,��Ěo���1�ǅh0>l}��'�z������^�յ�,x�.��l���ѫ�X��%�'��ه���_Yl��7�M@ԽE&�EF���hQ<�t����ɬ5�w&�T���ws|��������W;��x=Նѯӭ�V1��2,�I�l-�$^��NG�9|:��Sϔ�[�Q����C+����z+��Ѯ$���`V�Uoh�"�Mf��J��aKH�qM���s �:��J��Yۡ�&��\�D��^�[[�Ez��{����QLK�h��̅z{��P<��d�)%�#���z��8��a�/�1�l� ߱��������t��[�f��3���֏�J���E��U�5�&�LJm�<����[,#���BY���X~�c�g������gb�'a� �������;H�C�E�bc�j�\qq��=��d�#�7~��}��wg����w��n4.٫�����\�6�J�t�F>�F�X$_P�	3�a�|���M-�p�N�hz���-E_�L����B�i���㟀�	.��nZ
B��|֏���eQ��t�������);�#-5]ߺ淬˦qr
V��jT6ؕ�bv���ɳ�P�<�Y�e�ި����H�CRoJ}L���8��z����H������48���m0����$��͚���D��&6j<��~,;������-+#gEj4�
������0k0�m�%ص���x�E'U����֨t��)U�K�:�r�
`�7_9��CR�i
��iR�H �]�22<��g�]z0l���#a�q����vB
��T�6�+��46X���\���'f���d7�2�l��㤣����s$m�]gun�?McIsX}�[���:��pUc���� �H�Oέ���$=!��/<�r��A��D��\_���A�MW8�_%���F �:�^�pH� �@c����j�+Y�T�e�H��f#���x�t�+P%d��\���x����X%�:8r2����=Ρ��"��x�k���&�)e.ғ�}�pN�kV�{>���~��k�U����>i�d�������RH��1<g7`����π�ݜ���!�j���mU8#i`hە�bI��q�nK`�����0Е��Г�x�t�/^��{���|.��}�ã�5]�wt���ΰ���9Ц�a����B�;g��q�杕\�斫9��+EN)K�Sߔ��X�r@������=�I���r=�����R**��~��Y�����J�xn��7u�.��W�6����φz�ㆬ�� Zb;�����ҋ��ws��+_Y�k��dۮ��4D���V03�`��D˂�6٧�����Xc	�%�Se9�o�a�o\��T�zFf����@:B�̜�b��'��0irq]��8�R� ��Vê�Pee�j�ɳٓ��m?����<�VDa�+
��5S�-w��:����c~�-o���-������:lk�$&�V�g��5�'G�i�v~e��FV1�4��@���V �ԼYS�$�>�Vx�Ns���}|������o�AZ��f�+l�Uu������V�r�c������B<[�x����㌃$���J&�#��ZN��t�x�ܥqZ�d?��s���*��Mh�Ui7a�W��&\�>t�D<�E��P�R����
e/��|�1�r�\Y�������"�Ӝ'�0oU�?��OQ�*\,�U�>+��z��	�M�A���{�/�78BZ��Wj;��E��M�4�f��>`*R����2��yPg�I6��U���<�A�_�Pد�ѓ��h�U���H����кӶk��5��R,d��&yd� ���E�_[�A�9R��y���h��O�Pj��]]����Q��FJ.\�?f�����a|�<��'I/�^�y��	�: _����~(V;ݘ���uc?����*���WgjݠA���c�-]u�
l�����Î�ΈtF� ,�n�-�����ب����{��A��|��3�]u�����b�
�� �۱�S�$������3�W���#f=��5=��/R��z��n����{_@�yw�ZPыpץZlb� �R�`��Og�浅}{�HЫ|��6(ۓ�3�0\O~���k�Hu�����_2�x�j����,����dyw����i\k�Y�BKD;[6E�����:Z�ח����Y?��8#`hQ�;���i}�����ªKj�7	�-�6ũ����aZ��R���UH�o'�ǉ�Y^^����n2@����@Og�x��BHeF~�7�b��o�}gx"�j��}ܻ�ll<zUA��Ql[���f^m�]�aa�OJt�S�mqߠX#A�r�ܹ�� ����w]�u���^�-��E�׋���Zm&���\�Ll3�½�{�^�}����6���ʯj��"r
"���l����j�M<����h�������ڱ�Kتr7�m�Q��I���B��g_{����KuO#�ɄB�\�΢�%8���S?�-�V=����=y�Ƕ���7�$R�48��w�����hpMO���"�$!�r��u]�Q�C�T�m~�Y\�A�g���z2T��B���R3���E3�|�M�v�I���(J�E��qld=�I/�Zd�?��,�/}�Zˇ�8\�.���n�ONau�י$fm�|���^�[�4��/��> Ot��"��W�EK�NO;�������Hbg�$E�Վ� �4��b�=_�*���8�V���:&���*�i�؎=�Fȡ�I���0�(2�B�h��,_�H���e<�e�����q�u�����E�$C���`�j[ߩ*�;	E��)	t��Y^T>ш�|���$�2+��7dX�%�u���vu�vCu�z5��3O�a��|��.�����c�7 Q�=�a�7�9�T�;����Q���ͯu )\!�������bdE�K�X�v#�L�^ef���p��{��L-a�5,�J���}'Y޽��l��K�
��a��l�M�X�d����J♧��"���p®k�*D�-�����!�������GQ2�L�cG�P�<b��'�\zY��CwVXE.b��z-���n��Z���l&~_�'D���(��c���}u���{F
�'���SПt`�c u���j�&  �A�_�e8-��B��%˼��7�i����f�HXx��"��$�X;K�7��Q�萟�/���L���D2�kئK]0T4�B zr2�!�� ;��� ��u�0�%xZӉ��^�i7F��d����'B��A��i�P��uO��P�7'	P>,��AU묎��ô/��Ѻq)�5:Kuy�~e�z͔R�r���U�����`Hw��3��N��k��@@��(��u/Yi�K�o�d�F��4|��w:YA��)�\�Q���6�)���2�r�&2�/�S#� �s4�h�"���[�aR��dHԆJN>�0��)4��o^�G 5Yb�����0`���â�}�-���g���c�q-��JV���[�B�J��I��Lm����a%���y~�~����E� ظ�щ�D1��=�(��x��~7�<(^���%�7odP$n���zW�����$]uA�p�|p��@R�B�KM�BƎI84]qw��5W�/���_҆��Э�����{�=R̚DJ|V�D�Q�b�L#� ��k�B�F�6F�����=�
)x�䀎Ů�m.`p"b��_��5CU����bx������+h���E��TP���94�D-�1�4|�'��t֋@W�x��z�R��ׇ���Q��[�R�M���ynD�p��`��U��I�Uri��'�|J�s�L��)�"���kJ
�1�{�ǊI�L@�5��x"D����J��kѕ��(���bhP����w�9�������� Չ$�x��l��s>�	���~f�7�*����H���՛��<Ω#nuN�g���.�:�7
^��gR�&Ԇ@J2�K���jR�8��� ���v��g�SG+!z���T])\x���'�ڡ����T�rh�����`T�	A!<W;��@0{3�>0�O�KsE����2���{��o�vo=M*M��2��z2@�j�=[W.�ɉ�O�"��&ȗ!H9��MT0"����x8�D:sꦺ����f~J���DR_F����r��5��*_"��2����������$?�l��'[x+��"v�m�#�'��kH��JQ�*Qn�
���"RC�s�
1=E�'棭��Ś�E�	5XOOk��me(� ��OT� ��[�m�1b~M^�'��p����!=w��R�=�+'yhad�A%�~MR�+�2�&cɩ��5�
]a��K����$6+�N!�j, ��af<���k�S���l���K~��e�x�+��"`!A��V����t�WJ�.�h�;�U����Mh��Iv���+"���k��
��wr5�C�[�
9|�2�?7Z�-��V�'˳��[o2���Bb�vy�D��ͮ_��ǒh�^}<�(�d\��4H���!��abϊ�C��L8ӄn.:��^/��1�`�C~�0?d�Lk��Z����H5X�ĽTgg��0�;�VO�O\�1'	�� ⨈ς��G3Fݵ9����ų�;���0��ٝ��4��&�.�Z�\ !� 5��9�wW�:�j;�?���PPB�;~�mj��t�&��S6E✉</h���l41�)�+�)q�XylH}�U.+�g�c)���s-�߇c��5rG���M<Cƻ����CO��� Y�уDɆ�buڅ�3*�b���� �r���`�hc���4�_��n)>������^H�Le(3Y�F�ߧ����Wԡ��kZU �w�@vui��R��FI�t���ܯny:�G���Z��;p�]�,ݸ��lTyu4�q�+v�����v�5�"�s��K��a��`��x^83W?kaI��c��=q�?�_Ǵ�uܛ� ��۹��
W��NH�N[E��S�K�
1��&��ۇ|GЮPf�xP���
���Bi|
2���7V)65,��8AUԗ��A��[�$*�9�n���������G�d޹H �_�-Ka�VU���D��m��Xd?*�y�voȟ3:�{�"��;�[���gxV��v�C7��Q]�4O�k�V$i΍��@i�Y�?�ǅ̰hwq׎7���B��}'�cD�3�PW&��>�7>��δ�kE~c�0�B�tPļ�>#��B�Go�j��.	�A##'A��E�ѱ�EU�x% bqF��8x���G�� �ӊi�n�'8��K��$�������x�3�i���֕����Gl⮚�w�`�z�w�����c�p�G��iK�y�aQ�,q0�Z��Ę��߹GGŸ���u�Ak�ߪ.�Ұ��)LS0��7C�̕8YoP����~L:/��"y���k�_K�����иO��#}i6!���V���5U�j�r�t-&�h�tf�TQ_����!vs�f�?�[��Kqf-C�Y�,X�dk��E�� �>dk�}ʈ������E$!�I���eht��q,uJC�W�����1h��qy!�u�q	)�L�x y�����_��<KUM�<^=�+T����S�2�	E��Ղ{�i��5�`��Y���n�y	;�]H����C	�L-8�4B�.R������i:�g�"I�C��1���(�O�!&�����<A���L�!��5�$X*���UP�&PP٬)�O���p�
���q�Z��#�����s�����7@�kxD��AI�ph2��8BR�۲��t�Bv�a���R�p!�M��O�<v�-Q��oh��2����Y%��=��a�=���n���ی�@<���W�:%�ط������+�ی��$�0J�O����8�p�4X'L��]Y�Y��;Na�P&{e@m���Ӻ�P�7[��݀��袴'��K:��b��'�b���i�,�>c��@Q���>�Re�A�SD�����M@\�ХdT��p(<'y�9�E�)��I�}F���g���||.% 0"}zs�#Em�Y���R��h83��:A��0]�a�������7ei 0z8�OW�t�`w�Hߴ��d|d��N�ь�t^i���=�-�1��9
��&U��̱�g/��:��t�?p#��b>�L��X)��E�ھ:*�y�nvY�F'#_J�z�4��Q����0׼֖�`��T�Z����F.�Ds�i�T�$�T�1AB[ D��xr�u�?KL+��z{J��qx�Ԓ�Ij��0a*�DB9uُ�nO�
Czj~�!�u���\��W� �i��V�["���ŁYA����e<��B���t�O��$]/�U��ҁ�v���"�TǢՀ��>�U0�����*�v��1w�A��4%�Oޣ]d�d>km��i�K�Y;1�����G��8�w�����w9=��`�8�<�X@Жru�`jfOS�����6���g�C� ҋ�7�C\J?Y���E��FBI��#h�3�|�D�$��oWsk�n9�3j����pI4�½��o欙�)'E��1D���A�y��>��]�@�r�Ѓ��B%�gC��I.���"윏o��zT�Bg�i��l�a�Y
]�PS��*m܅TYɡ�UC9Tk5����P��8�G�SF[0�4K�c���{e�蟅�1`�/B��X;C�/�l:�ٲ,o/�5cw[BY�Lv�4܂J��e�Ce��jb����3 ��P���N��J��������H�?up�7bL5"<��Ȝ�m��Csh�*R��q�#*�&��}Z��GwP��R��sl+�ǚ=f�@�Y�Pq�4Z_i�Sv��5ǂ�Np�ʖ�a��ƾ)��)�K[�� X���	����T�A��>�],<N!��j�ӷ����b���7����g��l�u�LьB=�B���X�s�f�ds~�o�>��J�����}���˳��'�<�2��}�0�*8H����^%nٴ�m��f�m�\�"#��j���4�o��J��x����-I4$�4_?��.�އ�Mc��S�i�D�N��6��"C�w*�4�)�%���D����'������F
RX��YD��4�V#��AA|���<~�����DgV)%�g��b��ĩ�M���0���r�HFYC����S/`�G�[����pDā�\���AQ`���������5�Xp3��X�)1K�M� ��5ߜ��w<�B�|Q��C9f�R�oN�5rJ�	m&��#���K=��xWj�i���z�8B�/�u�,�!��hQ�L�B��R=��QLA�s?����WQ�$�RR��������A�m��f#PXe/âX�;#���MԲ �-�T�U+���v�b^
2	1�N��z���0"@4j*��sh�IsU���H�V�L$ӿaܰ��f���V�[$�@(/��R��\���SZ"(%��ޫ��5�P��|/�� �e����4��f�nH�]����E�q"�l�O�l��>�m�E�=؟cXC]�)LI��%�NE���Ҟi�]���D��QY�G��Ә�_�Ⲻ�������%�!�����l$Iz0��:rH�"ztjS����]�$�q���M O���g�k�/�ђ	��X�$�s}���e v��?^šx�����	+8�Q��a4B����������h�Y<�,��@'/��dha[�><�÷�m�>I	n�3�m1�y���CP���Ϫkp���u��R��OVk��e�Mˠ'7'��{9�~����=���'WtaZ^q�Wj�3yC�����WGQ������5���#Ͽ��S*?3I2;⑿U~���x��I���m��e�Δ�BA�X��I�*������N��(�4�2v����&Dqs)�UW��gf�<����B��{��ƺ�s�
)�ۼ%u��()RF����҆�
d�&w�$�S��+4��T�Ev�pp��3��8�Q��NGfಁ}mB;]V'+����ȸ��xQ�7�1`J��P�=���S��2/�Jی�j�]��ё�Y#��h�z׼�!E����LW��Eht�G%P�9���u��� ������2[�K���8�W捩ڋ��+K|���iT5�cWA'GKK7�i�}6���ِ��:�Ή��x80Qg�߻��E������E��k�r�蹀�O6I��O0%#���ʷ��1n��}��s���ͽ& "t*0�%D?�׉�P}�o�;�|^�B�q�ʤ��Q�ed�46l������D��	����?�Vd���
������߯��r���Z�Rs�?'�e��W���_12�'�+m:��p���cIm�� ����l��{�EO&�a������m	%��f��@����^�YL��&jZ���o�xϓ�87x�'�u�>�{�I���L�9�7�ԗ��0n��H^�m�-U���yn{��cS f�v*�Z�D��hմfz~/�#���>����®)�g��=[�
My0$?�Ř���*�����%@:�#���4P�(�>��Z$<�;�s��S������c�{��Ď��7�B�ߠ���:D���s����a�����W{^W�&j�8�>orf·\R���W����FO.�T�OݬQ�%a3����iа#������R�ɹ�r��ev�Kn���vC�{�L�Q���� �9&~j�u炣�6�����^4#��ɨl�;��Jz����qJ����UL!���[���{=�G��E�]�@���^�����u���`a�i�8"�/!m��W*��U�N�c��j��I�:mH�CC��^��Ӣ���.� r�'���8�޾�a)a2z+���[���H����baw�c��W)/L����p�>�ד �����w����c����Zq��x]pep>�	x�
���QP=%pa��_�J��_�����o���e�b���X�e�f�AfK��{L�����S�,� ��|d�K�gM%�%FSg�m��S?0 �/]�H�iظ�FR��)�3��  ���s��;֘������yMHț*�VQ��,d���&L�L.�ү̷YfE�o�S�U�����F;X&PSӉ��NJ��j�75j.�hd�X/�+ōavs�ę��O ;M�-�B�7 C�E��\��B�$+�j�:���iȗ*��q �%z�`�nh�9j�l�8	�5<O����W���7	��/y��.�q|�J�5��o��
��<���漐`��bM��&�����]�r����˽��%���lK=�0���/������qp�+��u��S��T���Vl��qۏp�B��)�?��`���ќFRG�r�p*	R�U`���)���Y�ύ�!*��!v��A�0;k�y� �b��'��p�k3�����ۥ�8m[�6�G��g�� �2��g��˵8ܜx	�}�~�+�O�`ʋ�b.z��1�M_�i���ջ���kj0�I��0������˭o��k^w�f��q��ȟ�ʝ0��"%�/iY���� �&b(����<�>��b՗�iF�)�?L��A���K�����bc��W������VX�p@6 d>�����{��x쓃���w�!�ou�s �_Lk��d�@��+�ÈUY���EG� Ǥ�齼�䅄�Zx������V.�� �B�j�~��>}��w$�]��ʳLtWo���� hk��JW���cՐ�i������.���c�zMBAc�Y4B��/�#�=�̻,H)�V#y�m�/�6�YY��.��`�bi��Ӎ-BI��
�8^RO�X�7��J�)9[��~��Y�M�Y)���v�Q����:��4���ؾ���ɏ�WI��Xm��b����o��mƅ��ڂ�s�`S��3�S�=q��t�/�����Q�5�i��Bw�0���C	]����!!&��M�*֦�j �K��B��Jx��6[}�o[�u���g0� n7���\�@A�7o�!V1�4f�A��|-b�j����i�
���<·�2?��r���D�YЃ\��K�-���(�x:��X�3:G}t�q4��,�/u[�(�j��i���?_�h�\�׆LCQ����%�x%��Yb�/j3��0���=<;���v<�7T|u��E�d�=+���vŋ�PGC�����b�@�A���g������ğ�B��{�׈�NS��Z����ꂿT���fJ�D��_�\j�c*���L�����J*��n�v�AO���k�qB�������Oa�ۄ�Ma9Y4q77e�x7^:ٝ�uk�4�_r�"eD�Y6��՗�%�j��j(j3�EǊ���^krq,=����~`��Z��Q�eyx�U֧M����2L��	�S��X�[���%D[(��=4���a��H�#=6	4�Mї��C��C��O2�B�Fc(%K%��)�c�vA{J�]���<>����<��i,E���B��4"`B�P�sVXED�@9/*���-���{Nږ���|��_mߢ���+����W�<�?gPʠl��,
_¬��m�<|o������Ke�3:w����o�Ć!��*7_ޱ��aa�p;���|���kĦSe5n�q�)�5�hO*&#�琸�kU�I"Ki�M?0yn�%�ɡ��>�_�p�����5�(�:�_����Hr�7v�'r ��Xo�Җ��σ�ԉqI���p�A�sT�����@_�D&HQ�V:>HM+ئQ��������Ű7h��*�P�U@qrp�����p�����8]�r߻���Do�B��,�xM���X���=��g�L�;�;�[t��;��e�r�=4`��#K(���W��X��5q90��˧B��·S��_[UW�Ib �ΐ�/2�}Ih�՚��W��&w�P���c�ޒ�9Mh�XD5/SUg��8*�0!�� ���nM�௾��f0Ulk�j����8���"�o��9�G7������M��Z�>l���۔}dw�a,�^�i�e��B)�f-�K-��'Ǻ�〚^b��Q�`�`�h��&H�^��B�Sغ!n�8��{(�&fp�
*ƾMgT��+���.��]X�`"�Uا2�v�@\i�@Ӓ%/�b�D��Ev����u�Q� Z��'�p�D�){�H#n�̲<��[ό��n�6�7&{�؝�dTA�d���ӡF�&�lz���!���b�1ѯ7�zY`p.��X��8�ߪV!>Fcl�)]%Y���)@W��8Ss`��qB\��QH:�N;6B��IJ�-MZIw�9�!�q2E�1p��׍���!�=����ќy�#���%�������7�R]�W�\B�_�=���I�|�E�iIX�x�n����wg�y�D��Mt�  ��fZ~��b�'��J�Z�Z��Y�w�m��e�����&]@q������Y;1�5�9�H�N��d=yɡ�������)���9DB�͟+�C�>�N\շ��D�u��`�%A�ALTN"ʉ"�!ݺ���1Z���R�qS���Z-F�j��7�7g�F���R�k�%������9��s����g�q�5{1(KQN�e�q���Z4�7i��e`����*�/�#���C���TV-�Z-O�����-"�ܘ��c2�5�81qL�`��m����ֺ��-5]񈅃��޳B�@���F�	eؠ�]
�G[�����=8� xM͹,��\d���lS�=ɉO���0� /�;|��z]�D�{AJtP����Q�+��x�KU�"��BӐ`�v*��k>0Շt�5�����F���yU1�X��6�X�t�A���C��!�ZP^.TͬJ+['83�´�������H�:��.HO�*Ŧ~^I9�4lr9��� >�ƭ�f�ЫᑎUf���&Q���شp�)=_�o�����B�̣b�U��2�YQG�_�4���;mf@�wh������:���F��%/����<�s8�%��F�3�_�}�������;����x]�; 7V:�UA�(����G#�}'8��Uչc�$�V8�w�� N�Q��va�#��a��Q{��W�� �l�69E\ʺ�r��:��f�R��:rK�P�[Jx�J��
A��b�����I������|��k�?C�^����Ѧ����ٔt6�R>6�J�E���7C,(�������^�uk1��Ev�tx�}��B�~oW��vR��dsB.w�C
����7�<���ꉖX���nF�Ƿ{S���M��n���F�
.b�2l�I�A����xD+��!�@�.��%F�����8��h l�l�wz�wl��Z�d���I��FI�z��;|d/\<�,�9u�it��/�P�dTm��?xI��4a����y*�-~�Y��ɛkS��>�G�;���|)��r�cb]���%_�f?)H	㩐K@(���)Vz�6m��W.@v�@3<�WlS�KDGq?��7l3jJ:�G�,���3V�fr����	��E���O��F�3\�?(��#"#&Aa��u`~D�����c���ty���F$R]�FP'���@Jyj��zt9�)�*���2��-�({-�k��_��2;�5��dHÎQ�H�3���=�V�ǽ�M�U������(�f�g~j��)H��}�d���6Oe%��VK��� R�:�	�^������e=���7� �"?��tT�"?��l�~�a�kŭ��'d�p�J5*	k7�p�� �ސ�e�Fo��`��*��F�ٔN2���($��e_<��@��p��tO��CÑ|\���ehDR��3�{9zJFdp��P,�%C���
t�XE�g(^�X����N2�(�"us�6^�.$IzL{
�^ɹ7}�l1N*+��g0b�����"���D_$0��Zi��ܞ�i�v �#5���pl$��q���tJ1ãe_��<�����3G�c��mM=RGl�r���� �6g���y����)��l��vol� &mc
M�˖єNy��d�-2�Ax_���^�m��&x���Mw�ҧXC�>dq����CM�u��N�)�0��|�H� ߭�} �N��5���!H'A��rE�0�;'�l2��X�M��>p�;��_�y;wGƞ�}���Igs�"��k������Nu�qC�˂_Ċ�y p��H�RS��ɡ�6��(�3`i�Z!��O��2.I��m�e��7Y�Fw��J:c9>97��~�hk�m�6��_6�/ �j��ҝ�1+]�Yh(���cc�E�[�h+|C�e�|����cg ���y	ʒ����[G��
><�3�=#�T�'�x��r�$�.ݔ4����FB>��)ٔ�����]�ʛ���^'���o:����j��9tZR����V� ܈Ca{�`���4w֒����LǥE^����������j������^���x�1�r� ����ٹ+�oY���{��M� ���X5�u��& �]LOq�ݗ��MlE'-�@��r�n���$"��g�i�� �8<3���T!B ��	��@^�Xd�S8 �gd�wl�i�I`^�I�`<%՝�tTY�����3������༹����z�Q���so�˶�d�d6�A���`�c�;��hצ[.S2��>%B�X*l!�N3j��rf��U��b#�-@y%{cAe�?��� ��V7ܴ��pO{����F����Z��ڨ��Aht^I�=GJ�Hq��;?����׷�S���#�	�������c�*�<�ْ�Li��zWc�s���`�w�LC��u�A�r䀲����r�\�4.-��$���2�lP����7�U>�I�ˎ<�@�8c����#o]�/ڝ�&�S��c��H?)0�0J*��4��O
N)sz�5�2,GϤN��R!_׺f�PFu����]����x�t)b�No��9D�8_��8��o�����Sw��S�
Y}���qܸ���ꌛr�bR�����<�G��D������U�#?����u��şE�����2x���Za��Ⱦ��h.HvR���1��(S���N[�\b�����gB�vVSa�4�<��j�i����nSgt�"HP�ʊo�zw��� ������h��K�c�4ƺ1^
�&��'F33�'
�� .ȧ��Z�ٮ�I��:�T���*�0~fկl��;m7���7�VA������Lv��Xc۸�~=��DA�^̏G��=N�ʴ�ԯP(�'����0GI����ȸ�Y�7����A��L�{%��җ��l#����j����|��0a�!�X*�_c�$�M�3��m��|�W�۰$�[W��
�n�k+Th��Bq����P{�6�0]>������L�x#��| �O6���)����E���aH�A�����*E�MOX����78��إ�җ�u�-�:�VQ�5֪��7����*/�SHPid�;+���=:��P��6�˛����mn�E�ulv�v�g�ub$��4�i'љU�	Q�g��u+�͘�m�n�z�+	��&��T��e�b9}�`en0i�P�u�G ���	�8�g�HǼ��>��\��D�I�9�E��ɳà`��]���w�LYJ�*KG޺��UA/�Y�� aq:��A�`�U�o��B:٘DRXC�Ɇ�*����-������L��^,�}w3}�ŔQ��Ϭ\��f�ll?�Z�Yy�h��4�eOn�h��}�l]KLĥ�"P�ʗ�����1J^R����
�45E�PlOA��� �<4{��5��F`�N�_��º��Zz<��ָ၈�(�6�;��D0PU\mv����{w�v������4�i�ϳg���)ru[��>f��f�7�RRW���tqg�x��<'ӓ��d����W��x�OZ*O��(� ��BE��Yi$]}���cꬦ#G��S�4�gC�`�F����͢غ��`���>�*�K��	F�I^J��q�'�M\�����x���D�M��^���q@���a����>T���|��	�����m�_�W%��6t+������At��!Z�F!�DiF��e4�(�T�?�s"<;�yqg�a�^��E6-�$}�*mޯ�⬁��]Խ���T,��EĠ�eEƯ�R+�(m�8C��O�+'JQ��{Fc!ͫ^2O�*�����e��m�7�]T4��sU6DQѾ����i���E[�l �, ��3x3O�QJ�$wX/|�3g��c,�/(5U���R��D�?��n
���;�X��,�����Ĺ$-qgN�߰�*��J�ɂ�{W��g�@_}� �~'Ȳ�P��q��Sp���=��7�UIk�7=i#�������=+�Z��͸*��C�n��{��|������Ҏ̄����e��G��J�V���Jc�p9���?R[]�!���R��.Y��FWE���fґz�ðK^���ui�_�b��+Up��.�)=x�WY�R �Y��/;`Ss�����n�:9t��/�c�/�I��2�e�WYD��'��I[p{ђ��2��%(3Y�/#2�ުt��ʡ�zpA֘���g�xx�
��L�,���I��R.)'�aj�w,m�9"S-&�+�r�Fb�`��]0�|jZ6�łk��`{w�99��%SC�d�9�/�D�]�#�I[D[��=`�=Pb���U�M\0|�n�W�|*�kPx�BD�R�6�C��٣Z�[`���w&0�%�<]uD��2���'�eQ��LW'_D?X�`�*�C�#	w�3�A#FB�'dc]�e�B��.������?`mJ���k�sf�=MD�`t����vA��
�HA�殫����Ih͂Y#���w�Qǜ��|�١ZG'�"@0�=70�9x<��[,Q��@Dٿa��N�[c���S���{��5��{b~�,0�f�[��ω���U_Č��[�
Y��}�,c�ô Si)k�[%��hù���`/^^R�kw��׊t����&�u���	CD@�t�گ��@W�X�_.9N�,�7�3O��FG�9~�amP�0~��Ͱ�E������I���ٻ���x|�O-��,�d�*\K��v�us�������tߣ�?���6��/2<T��� xj�'�M3B˭0�����dM�R^OP�* �?8i��!66���^�����5���}Pm�	n;��w�p�}�r�Q�;M�Jn�M+����AGuӀLE��Y��i��PdH�s������qB��lҤi���2IQ;�%�N�x�[br�M���-�}_�t*�R��9�dL8
?k]d�imq*ݸ�\F�ݽ��ʲT>�ܖ��8E�	>��EYN<w�Sܱ��w��\�7�Ѱ3L��Ws:�#s(������n��{���0�C㸥۠���S�y
��zyyoO߇�=�D���x�����U���ҍ8:�� S��������mX�ko	@2�q�^@'���J�S�h+�Q7*j z\N
�9K@>ܛ�_W�0�A��$#a�xq���Y@�X�Kt��9��w]ݾ2W��F��P<jP[;@���l)ͺ�U�rlI3#'1��ib��O�Z�� ��9l�����)� �"��}�QCj��_�˨���{��0�1SA0��C&Ԩr3&
��N}�خ��UR�t�d�PdH���{��G��hR��2/-ìa�Ɇ��(E��7�J���!��u�I�~����������&�Υ�t��Q��OmXw�g	� �d�o�s߉`Ť��J;��p1;�
z R��W<e�J.����Rk|6��02�:�:������\3�S�ל�yUs䬝�b) �ъ�����n�Z���
�	�?���?��m��=E��*%]��(�}��:�t�a�}�~��F��_\[�^W�6|�,�&}��-�,��3��>O�����q���+��'��F�u���2f;�s���i�4�O�;�:�9œ҈r!��Z��wL���{=9����jq$!{��ߣ��~C�4
T 4V���p�u��2C��8Ozw|���ڳ�s�+h�4a	����3�2b	��F�8(��+ٖ�'��n�;����H�H ��\��R8����C�9U�G�Vy����!����<�(��K@�מU*��'������*U����/����3���ޭ ��G�#y[C�o��f����(ɰZ4���#���F�4�]|M�&e�!���Tv	)���c5C���ǋ�U���`�K�E5׼p��)�A��v
(�d4I"n�Tk�j��[�-i�)l��Q��2�O��O/tc�.(u�`�N2�qɆ`�����w4$��X��y�#��,�!F�ms��pD1���mr_�A���G?Eh��h�L�߻�˭L�)YfI�;�Rm{��j����M��xBj҈C2B_i�*d�� ���c�g
yC���p�C��i���5r���l�k�`���b��T���	�De��δ�'IW���⶷u��m�]D�z?ϛ�iEേ�1�:�W�E��:��GS�ĩ&�"ñ8�`�U�&�W`�*ji�(�=5]pN$�ux�LU]���J~&�*GxEC�M|��9S���k7�|�l�ܥ�b}*�g��_L]�3���
���AC�c¯�Y�>F�tȃۄN=����Fx\�=��˦�7���m�..E��gyj�`�x) �v�O$+�L�@�R�x]�����;k1G���FB������Ŋ�M`|0��S]��e#��V���/����/�TLQ5�r�ˉ+2y�z���@a;�Ygձ����j�?���J$�������z���&tB�~X�u�U$	ؿ��5x�� ~W�M� ���>�~���a��(�p��R2���ǤuF[�z�nZ������X��O��ڑO��tS�^�[y������ȑ:iD���G�#*+�Q���r��Ҽ�γ����ڰcz)n�ui�c�Hi�P�Jy�=��e�v�ٿh��B~Wc�^�ֈ�������Ԟ��a��+������#��D�:�n�*{����Ky�>������Qx:�)�^��k��c��wC��������,ö���3��4���-q����O��x�#i3l����C��=g �.C��̤�!liJ�/y]1�JW�t���׆�a��np����*���i��8Dp4��D2�?%��z2��@��'��JU����������Nj% �!X:�Ml��~����<�\O��	k:���֭D�:R!�>Ѐ�'0��Ӷ���w����`W��t��B��;�^{R��J��G��^��,��O�[�6��wT꽝�w"��=B��"\��n+L�QV���U�6j�YJ�"u�_�������T�@H$k�I��Cfv�bLAf���g�6	�r>���w��g��UC.d�G��J"9�7}5�,w���}���N��{ߦ@��m�����$*}/O�.0�̘	Y�f'A�Z�M#,�τ����8%[�P��� �8t$���Ӗ+1��'*}L����Kw�r���
C�hf�|}\�x��cƋ���=v��vE���W��7��!TN�@f_M��؇��?�0�F���B0��޾�]���L׷E]A�UD�k������ɯxK_��5�j���'6�0�F��jܲ�H����	9O�@�Ek���y�[9^%_�a�DH������u��/��*u{�s�{p��1Ɲo�w��g��� �f�����qo<|�Q�-���A�G�;��X�'��!������z��=g����Q6�/���@Ţ�΀U^^u코ܖLM��d��X���&r=�����tby�\?��?^g���X>J�,�Y���q?Uy�����[b��)O�O!��zs��+T0T�8�W)3�$N�6����@04�C���i<8���8�/ع-�D�3��]���<��;^�\q��(��d{˔�L�q�o�}^��6Þed��RX�M9q7Wy�����!g��`yƊ�z5x[��`#�����3y�:J������q� ��vx��da-RC?�����RתZl��4@�*���ơ��}���G"��
��\�̴qR�6�̱�q��4U#��u-���C�RN��:����W��F�|�]�I ��J���揎�Z��Â��2v�	U׆��a��h�d�f�r�9�����K��]1��'�1�_���p��	�3<�k74�h���#�u�X4^Ֆ
���a	�.\H|/�l�̲S�d� a�i~���b���.Ό�#i�IC��U�'��Q�q5+�	�f#i�%�o=W�@�A�I��$H͉����u���5�2�΢�^��GTa\� ���A��̭��
�k��֐�v�f�=��&Y�QVw��� �-H�]�����6H�D�wW�[��I_���R���>[��-Wʫ��w�^g�OnG�V:V�}�u���*ey��ak���*�e�'���VwL);jh�M� ��c�&=�Wj�j����������.��DV�a��)D��l 8�|��u�n�Xh�!��R��D�����f��;�\�t���2+'���	ô?n'hNF���P�׼de�
��\Z��
?,I�i�@]�߆$n�"���:���O#L��Z�(�� Za�dQ�Iʘw`Dg"�������9������KD�~�P�����[��J+:�6������R����	�'en-�Y�����4am������AD[���y��7���rB�z����?H$�뺀'��L�5!|��J�-}�6jƟ���
8eQ��#�A��ә�?��&�����aX���"���k(������@�-#`H���)$�AM=�2�ȿO��ңȣ�^vP���74DX��D|��tZwT�>d���a�@����)����K|�-�h�����n3��Gy,ew�+e��}��2^҅������m�չ3�8]���#�W6����p��S����XH�5���w)A';;F֢���T8&�{D�<�z�N�$����D��}���L��/�Y5*��Nm7փt*��mQļ�JrAPT\iV��:(Zn|�{�_�c�&�8�	�Ht4d5Ǖ�^��OfA$7|�Ȁ��
v9���g<���H҈��������!`��x~X�Ȃ}����[�T��<��|_�]�.�9��ش��7h���ꍆ���(��%8��f�ޯ���������?:���9�̥�,�c*�����x�Ua@����pB�"�͈�F��x�\>�����}����^=�O	�`{������ԡ�<T�Po1�Z��P#f�ζ��^��xG� ����>k���V�m����ì/��T��"v��6���'ҝq;&�)����Ӓ�c��[���>r�@�v��pPW�.H�܎�|�[k���U�S��;YYw�؉M��Q��m%��V
�s��0m3��eJ�-�&�v4z����[h��jx	�U��Ƕ��!���Sr	�+7���;���k���o��܏�F��Q��]F0�G�[������m1AkI[ :l�n@3����7=%d�O��I�ʮf�}4
��l��w:M�|��[�E��%��0�}GQ��V��@oI���yCZ�����e[N�Js�v: � ���ac/���~iP��D3�����%o�6�"�h8h��H�t,V��^~�̷^�kY����ɸ���ɩt�Z�T�
V��(q�o0|CH�(�v�����N�j)%E�|��;7���܉�����;ݾ���9�c��m��z�^ �|F{�=n+��L�o/��;4����%�I���#B�:0襖H��#)����x����F��r�������R����?�s
��b�<�>Ã�<�:�>�J�X7��?	���~��"���Z� � ��N��~D�X[�5�W`�uy�ƕ�	�Q)�&��Ep�{ ebLr�_�܄��}'�>�!��Z�É���B\�K���H���=���Q�˘���."r<�5hNc�w�c��L�U����Kf�I`M�hYHˌ�N7@9Rr�h�Ŏ��K�͗u�/ĕ�ʠ�6�U	ZU�KP�h�U�y`�c�69�d���/s�c�K��<<~d"M<ً��Ӵ���]?��p#�^�'^h�O��}��K��zE�$��N�`���O��uM4/ɚ��_'��V���2�M���#�Ƨ�W� ��q��Қ�n%su�t�O�Q �����I����q�M�,��[�1�VkU�A3I�I�����Ƞ�@8�g���!$�[	:�ЧA�y��98��Ol��,�Ը�U���9Vcա����{����X��*��A���M�H�I��K؜�7�� T�<�,vR�x�M_X�����U�w�{3�'V��Mӣ�v�ݳ�t���H�J���e5���w�j��%?&��:{�i���Lx�3��aw�ub��sX$��jCd{ܺ� :��PP��o�����@D}�=!L�Z�$$��/K2N�W�� ���9�U���7*��m��͸�l���ƅ ޔWQai�M��M½�Ϣ�R��1HǪ4�����ENǥ	Z�G|a��](�|s9 Ҡˊ�ܖ<�bx��W�̯LU��6Z���)��K'O@��]��0�_��5���G:'ȇd|�2̈́2"||�Ez��Ο���H%���z���)�<{+��)\���J��'�)�d�9�� I�8��f���&���Ys�w(",V����gh��䉕��yeIn����
����:q-(�!;���o�Vc�1��6\H�b�<y�U4X��r�V��W��	�,�6�I�_Խ֌�&)V.s��@zw|W��$8�)���;�5)5� ���_��S�;LrdlW�z����M�{6�%եPO'�V�RzY�pJ��yor���cb2�x`��Uz��:�s��E���R�GŦLф^8 ����ʌ+Q����ŭ>�{)f�m��0PG �^��k��V/WFpu�샓?y�4M..v ���k�]�$��D����|f��U��������b'�����m�,�GE�4u$.���_�x�<�v�_HդT�q��XYDI�@��)�U�L̓)�Ӏ��$�/�n\H�Ɵ�Y�{sc+�#�g�
=w�����H�u��3�u�����)R�Sp�{F�$^2zB���э:� �KWM�<�L�� Q���G�'/.LYF����3�E 8ۖ��2��E�6[v�y�1���Z�">l�[��wCU(�%2i9��o��r�F��JL�Rf��jҐÿ�a�j��Ξ!ے3g���o�_w�k�Ҍ~�~H�S[O���S���r/a�#1&��5lX�[/���~��� N�&S*v���f�=�W��C��(�OF��-1�w�8`Zi*�O��*���Q^��hRZ���[�zC"�}�^Sp��ݟ����A����KC�cS��5?��A*�n�5��jc7Lu�:"����Hhi��Q
V�s��/��B�L���;�T�`������^�G4���F2Z7��>O�6,����g8,\���@g�&,���]�BA�j�J,��$��{��乘!���#���R���IU[^��f���g��4������ҭe�i�vp��er�)�}6J�p�*���Fn��ʓg|�9X-^���yY�����DM��3�ko}ψ�:�bwYY���C�)e (v��M˹���g���؛�D;�Ʒ$�� �*�w�>6?�?����0���e�;�sAT�X����[���c���^8��Pէ��y�V�*������ا*S�t�ό�q����yg�G���������
�X!������f����Ƿ�B>1姗�{aL�y��`8M��9�]X��˴��w�˯�>3E+^���4U�vm���V��55��ӧ�"L!���J���O�?�;��NT�u��ǅ�=�9_�/��&ϖ�z��o!ɽ����O��w�%�?R���3|����%6	��u��aw\Q{l ���Q}rs/����1G]	w�y�V�~�$\�ߓ-�Q�4R�t��RP�m3Q8(�|�Wm��H���˳*�xY����B	굽�Dh��C��[�f##�"�)�ge��A@ci�%.f�RZ	�(mR릊�(�eu�~���tXLM��x%�
�.(�u�ed�g���|rx�@p�!\DAl��B���ȳ��9Q�ʑ�$��稼z
�h �&����0*��ĨĹ�� �u?��O�������������E���pb����	T9'�GL���%���*@���fU�B���s�T�d2���Gb�.��r'@0<��h�`T�JX:��ٽ�Vʹ{������'���*����1A�u_I��L��e��Q��0�)�ٸ��v�Hm
9,��_'��^HF��R���3/�sW�uq"�lϲ6D��Sk�Qm%�_�90ȕ��UL4���t�����rD��;Y���a;�ஹ=q�����2� {dՋ��2q^T��Y��>иvQ!`��P�AÒ��C��G���n� ��4#r���dp]x�� �rU��_ ���y���K��#n[�&C���O����ɫH�"LC��9l����,������(�RR����.Z;7h��E�Fc*1(F#�g	NR�Csof:��W
)
�|Ui�u��Qz�,+��ٟ'r�J6����Ȣ�Lۡ�%�h��8`/��&p��_��24Y�-�aX����Z��3!`��4�{d��Ʋ�,�7���^�w�)�9^��}�Q�r,����B�����%G����0˶�L�ø	�抱�|�YD��?��ff?u#��O��1��n��m'(K.�"���T����(�=ɇ�]��!�H�wFfB�/j\�c��޴Ϭ΃b��("I�,��'"�=ݗ�>[�R�]��K��X6�)	��v:Y��;�w�짔9���f4=cT�(����g8[bY�=�\F���P����������a��@�C�M��M��<��"b��>v�]@(��(|�ۉ,�6�%|��;ǵC����zߏ�x�a��ԜM=�{B��������R����߰��m��Q����!�yd����'q���0_��5)&�#ި�N�*�����
�����d�X$��v�I4��p�a��z��I~p��T�*o�ʶ0.b���v9��^���^�t�'��B2�
y�V��
2���3ܨ�jx~=�A�G�'bm����y�*k�j:��Ct[��H�ȔX��B���}��	�O�����XC�"U�-�[�b˞�=���0�4H%�N���%H�m�E]���q$���<L��0��5N�@Ҝ�
�9&-�[�+���;s��)��P�
� �Wc�v��LJ��ٔ鋨a�9?[y��9/��4��\	oƻ�$�㭞���}ع�'�M�oQ��u�R�z�D��j׈��+pG�+I.�s��G����u�nm�@�L)�{����m�
0���lE��J����Q>7��^�"w�j� ��f�|d��e��~��=�S�sD�s�pc���V���-y#�ڥ�b�ԮD�Qqϻx�.PkSs���a/;"%N�{�V!f�2�LyiI�iVn����Vp��xS�3�tMC]l�_+�u(U�&v@2��I�׽��5�ʒHx�mO�=?j�O��	�ei��Z�"zhDDu'{��_-}K%�f�˞*x:sg�!K2F��n�� Adn���m-ٯ����<�y���{w"�\p.@�x�v_~=_���Na�[ Hs�r���\4���l���-mf^����:�j\�^��E	��!�EQ��!�cLKI�Q��,�;Ɂ�q`���.���ZX�{�7�޼�ܒ���?�&�h4���&x�B!�<�v��-�n#�D�����gG�Ӈ�}\�G}K���̚�6K�:_���>�����������=%�!>;,񭻿��t�)�O�kD����{�����
H;E�\�]��p ��߈�EL��ȷNF}�l����U4����rC�C:���O(�Q3%���$s鼵����kʵO�u�"!��Wa}yNp ���\7�ᴆ ���W�oNH�5OO:Ϳ�Ʌ����~��c�Z�o��~ H������c`IK�� �K�N��-v�X��A�ڧ�c����g�W�2p��kI{���~�z��҄̂3��"�"�������AZ�lх�������*H�&��QC�"�Ag��K�f�*�E6&�⟚#C��<��x�k���W�_uӿX�����j��Y��6����WV%�SH��r�J�+a��Az4fs�m6Ҿ�w�ڥZ�L�*Vn�ii�d}ǂ����B�%,^'S��j�1 #�0���g�?�*��V�V�M��p╟�6T��|ԋ����^��i����	���A���{P�yn[�iupj�\��
WФ�\�k�i2�ʉ��i�Y2s��.N7i`�ў�nC	6(�H�/N50(��i�r��_�%mJF����Wc>�z'.�0��e�&�H���(�a*թ<O��+1p�$�u���� ���w���8�����$�;j´��=#+B0�lZ:Y�^��S��1�.�dU��+��H��v|�5��Z�'�P��c���C�t��D��+��0}���7eu���%%]�̰&@H���=bf�iz9V��#.�D/��&�ϴg��r��)���%%�t���;��ρ~��?��b�b��£אG�v`㍪���
�a��+:9�<���rߘ�(kϮs(�5���V;X�|4���S���m!����;&#�B�$����ug��#�2S�t��Ӗ��|Z,�M��(��;���G���X>צ�lMw����� �Q��
`��f��� `k�z�}z8>T����IR��D�C�`}����8,2�4S�4���[��{>L�=�Wq��k��n6�ᯂ͝�ey�,�ND�$����(��YM0H4��N����C��ɭ�%���F�=
�,1ށЯ`ú� �\�#�;�oz�������~~���? ���[z�M5,O����<Ď<�C�X�bGc�_�;�K�t���b����aۏ�E]��39{J+�� Ѝ��d���ㄝ��x֚�J� ^T�p|h{�t���7R�,��D*�V6��ut �(�0M���{w�/&��<y�UT���x��}�������R�S,8y�9�na��{��H["��<Q���iPY�\��Yv;Qoh]����}2�X����o����ݥ�j���Y]���ZX�?�N�Ձ��<�%������Jv���	͘ӆ����Ɍҩ�H�V�::�d@��q��	~�(��1�L���Ypj��R!��������w�˅�y�􊉳��Y��)}�e>g��ʸ^�4���S���/b�Ҙ�D��hB���D�P2/�Z�U��֙� 0�+�?����؜�^�ޯްu*F�O�.����g3㵞e�/��������z0n�_-$Ok]���]�B{b?���]�7����Q1��!EjZ]�#���>(�U�+�s)�E�aS�s��+�W�	�hϤ6��Q�K	_���Mt�,���Q-۳����n��!O�~�s�h4�V���h �!�!v�l�/
�;�>��M2��n��E�ǲ���xNb_!l��JS�x���n2Hzd��x��,�ޓ���ܴ�(c�fY�Kt~ R�-����I Yc��	�`�ײ�Հ��d���I�GZJ��cW�>d,���%D�΢@�es��5�L$�c�	n��z������Ώi3��*��V{�_�O�K��T��U��A�	v��c�r�b����*KC��'��)�w�����;�>X]��yl�DT����]��$����6���[(Z4����N�Z��Y���?��\��2���W����d��M ����&�	<�1��j!�����j����&�5�d�el��Y�� !�T~4�>��&�F��Ɯ�G�! B����c��m5�=G���
}��RU�������u�m|_Yr���qE�X��}煮4�����Fe��6M���a��4Q� ��}"�,��A�NqL�'�iMB'�Dxxrф��γ�Nj��Qʇg��>�a/���1��v�*;�q�d�6��S���MO��-�ZGil�=���]g��_+[`����s�},��%pMu�8�6G2Q	�18�Q��9)ӎ	`$�72!pxS�v�����oB.qǪ�X*C��-Ɂ�J�^a�Xh�w�ޛ���[��i��+,�k���q���.S���qP٠eF��V&�����2��J��+ٳ��\0Ω��+�1Kw�.f eY�� �@ ����-/�Z�οF;p�>��I�jO��*��o�2\G��uqA��z��7�B�f���/�I�ߞ�/N	
Mu9�~�;�V��z��7��1��c��$�Z���˚' ꐚ�7��V�0��DH�K�H)ty���Vq�:G�i>o��3ya�<��<����|�3���J�BP��Ö�km�ҡ�!*���n_��3F�����m���V���A᜷#�,��^��o�R�	<m0%;�5$�J)񸺧zZ��shْ��w��J�w��)'�ک��;R(�(�#n�]#�蛤^�M�ǡ�c]�ax�}j���׉t��I�F#�V��=g�TB��ݐG=.�F	0�
�w�ic#�Rg�8�jc�v��NP��qМ(�X�AZ��-�Z>sD9�ǃ�>�v1�̾U-�R�Ln< ���e��Lg���H��\	H��抠�8 p�;��Y�X3ƾM��=�� x�㾏��Ӛ&7J{�Z�#���d�P�w��>\�=M��9s�j6v��[cސ҅X��Ͼ@��dq����<�X�Y�G��,����Ɇ:ma̞��X��V��H�q��� �h}��B<�.a�J��M���(Ё�mmQ ]���c�_5�+���Hju��%Z��Y�k�|-x�m�O�:4�+RE��q�g����{��vc��\!�`>g�"�a��k	)n�Iq��"����%���S)��J���?-x4hȘ����?����s�VH�F57$����؎�͊�و�l������E`���^�3Yf.X�c���}#���`�%�H��E�·���E@�������:Vt���^V�1����!���~��b�)��1=r��H�:�c	u��ګ�N`�8���Z�ŕ ȗ��r�*FvȘ?��U�닳��mE�GvO�q���I��I�x\u�3�+��!�
00���TL�f�v��Rl���\&�О���+V���}�� 	��PH��e�O��C�eY7-�=x��:�눂	e�ћ��d�g�h�<��\��ى�}��c�f�iCqz��JxD���3'�R�Y������C��̆�/�����->a3�n�H�p���1&�ƎL:�.�e�ķ��x���i2n�O(�y��\�R��j*���	��n���*
��F�8�G���9�*e�$G̷`Amj�hG�����T2��2K
�I�_8�����Pv��FD�s L ���=�9'٪e`�B�V�oy#��*��"�0����.��ݫü�Z6�!y�ƮKs��=e�E�|�u�M:%�W:mض��7�I��'3� �Hc�1�ω�8�W�N	"�#|�ߔ1n����&�ø�z�{�(�1�	��ag���·3Z�pr���̼鉇�8�y��έ�>�����ٱN'̘��`��(ʊZ�Է�Z�f~:��u�C5�f&<���\MU򺬢�t�(�1F��6�bEݮPKm 
���)�r#�c�_���;�Љb�,���i���8�1$p3,|1\$��z%����q5J�㤻�3���bv�����I0��"���6(��wT]O,?uY��$����S�?AV�Uŗ�i�@�7иv@y��/���!���!]��~�J#M\=�*tm���w"��z��)��kudp������+���v_?K�$c�6˜S�x^���E:�F�RC}u��G�\n��պ_�p�f#>tl�J����ѐ;�6sт�MvdG�u�ҹ-a�Ud@���[|枙p�]n�c?��/��k�p�Ҷ�y.���!��	^�[�]��ߨ�'�_�V���Y�Ў=���1%/�hWǙ�5u@��g���������qL�"�$�{b���P�^�p+ʥ��^)c_� ���eZ t#�a�0�ʳx$�~P��ϔA����+�Й�~mƝT�nYP^X�����j2f�7���)���@ ��P�2�hi��\�P���?��4�������N�aq����P�8��A�Lf��.�¢��V�ڸG����P�lץ1�X�J�q�r�~a������.Ap,@{���Ѥ4���9������Q�ΑR6f��Z�[E�C�`F��̏Q�C��%'�35��$lD�d1�U�`N��"�Zfk[_���<���YN,ƾ`� 
��(����f�/��2�W��J�F+ۊ��d�(�޲4p�G;�U/�_m0�\���7�Z(D������ǁ9S���!s:�#S_��d�F�]�T����Z$�\���n��8N�,A����Є�1�u�!�LY#�8\�gjb��a�����2��߼�f�׶�"��h�������u=\|��o�3���$�(�bѥ��ר�	s�[�@c�b��Gb���c��ش+n@��}�p!�q*�����o��Y�[y��B��k��&���5ր����p>s�I)G׋ ��C��=�̇2+TpL�<1�ɧ�?�[��\�"�����3N`t�^Q���S@
�[��7U�L�"�C
I�喙H��?���Y�ʜ����Z`�a����9m�S�c&��g�#1@a�ȑP��9^b�?�TVt{�?7:�e/���X�������½@�k^1W^�ѝ0=]��R'K�;ҕ���8X����(��[	���H���O��Y�J�\bI���x�|���:ֵ�:�"�ǻHOxg9��j\��u�R�C'����^l��c<�	&>�9o�@������`̂&O�Zm-B��m*G�BI��$y��f�c(�B���`\�JT���2���Q����މ	c4��W.U=�Y��D��8���i)�\&�z�3����O-�����&?Q�L�<�jzg��eF(�,^b�-㋫�3���5���� u��<w$g��~(����F�{��@ڞ�	LE$�#�J<.1����_h��^��1�9[�GQuJ�h���}��-����5?��+d=��a2WSBc�v�b��R��M��YB�}�ϖ��u�9�Z�N�/ޘ/�T�"�*Gv����3��<�$uo�
;
��ť�@�4L�E��"���:_��t�t|ʵ�A]����Z�
Bu���X�����DFD�֍5����s?|4�<a|겣t��}^�b~^[P�s�=�,+� 
4u �ԠVN'{m�XP<pԏ�}�=|�_�l ��C���>;EA�O2u��qi:�Ks��T���R��%��W��;�V�1�u�A3�N9�wֻZ.��!����|�R��S_D���Z���MOJ�F���}.�����_oqc�%����ɞ���MU#�5:�,��0x���+�o�q+V�{�t��}m��tv��|�"�b/��,�9��jO�'�oY�@�^\xq`5w��8@6"�k��P8�%X��r���p9��8sk�^a��>�Ks�S�yF�E��d�0,�c˅|��k��!f���~w��z��[ ��ܟ���*���[����#�#x1�^5�lYY��5����#�Wni��#�|��l?���P$2w)3�u�����0/�� MN(�m��� � �i���џ�ڷo*�p���	3N=?�3�R��y���{-[v�)Q��F\���m0��f�qX�ՠ�ѭ���/0��񥖄��ß��>�}�8d�8���K�)C�v�w��Vd�ۙy]i����F�~�O���.Z?9���$p�a>����B�S.Z�
#涼s~����b�x��i|pU9�����Y5��ﮯ�y,y�%M*���P`���&�p���a�0��\��s�(��D�A����>��U�E���� h2�
��^��!��a���ۻ�..?ݴ3�w����:׀��Lg�Q���_�@��qU�gr�+?�	8��XS�h�� �8T;�7�{{f_�4��s��౮��Ʋ�+C:���(#��^g96pF���9��l��Ko|�:��ϥ������3~�B�����Yy��%>�Ou��|�AT�kp˭'�e����E���06�����0��iKX[Gb�}p�D!b��҅F�/�e^CW$}gq̲Tg������V�f#�F�
d==�%�HF'�v�9����liO5�4A@�������W�9����[�F��hl��m9M"������xOocnQ���,a���2��/͑��̶#l'!��0�[1�~j[9��;FLU�ך��I������0ݜ	:�o����9�qGx������D*5XI�=$��4/~�z�7�R%5���_�\)����]�4s<�ܮ� >�k�$TR�?25�T�$o$q�v�9��&��йj�o��7�i�������6��*.=[.a��1�d�3!K�ءة�b���<�:�I'���=��Dʹ%���G,̸���lV�if����f��|5��[pa��	Ou�t/<@�^�Vvʵv��5�r ǵ�����;��[�w��*Ue�+9����;��=�O>o�C�_�u�G>�&E��'��V��7,��
�%��u�,mr��t�V��1�v������p09N���|>a�Y.V�&?�^i$�-
�������\����~�=�e��ӂL��n�������cI��1UK7�4r��y�EM74��cb�X^�"�q�lI'B��KY#�� �+_��@ DV�Z�zɱFX��[��?��HAJ���^ڡ�G�z���O�"ň���}�����U�(��c�R�~�(�˵噏Ö�.���
�Q�g!�O\�6�ي���%�+�(�їNz����Ϣ,~��y�P�����3�
��.q��QO,�_��&W�;������Xⅻ|R��Su�1����M!$��ϏW�X8y�P���<�� ����K�>ywT/�~������zc��[�+v�����ѱS�N�O�M ?R�$�N[���ȇ��������cb�����US�������Q/�Z?,�ǫ\=��ї��(~� l;،M��D�X���q����X�[j�,�����$A1U+L��O��D��i�,R=i	������Ii
Dc����ȑ_'�)��+�]�����w��z���^��
�e�Z�w����-G	�	��)Ō�q�f*i��y�Qi!���1�ˤ��03�`)la�#B�s]�[P��f�d�aClj2���%NGrEĹ~�7� j�7ʩ�u�n��JeR��v�'���=<6<�X?�y��!�D����շ(cK�j�b:�eRV_G�^�^����v׬P�q��O�C�a=4�� ��fFЮ��,J�ω���wL�h\m�m���,���f���k��78=���D�w���KQ_ 3��	C��8��VAa:0�QuE_�\��%�~�P1n=��yC��-⪊��9V��0+fh/C9�qV)6��""�WX�R�}�Щ��v3�z�儫X �>��hSW�]� ���>D0],��.�b�ޓ���m���ǣ߉���/୮7m�.��ԏN����n)aQ�e��w�V��B�iʨ��)j����}b�Ȼ���Q0
^��	x�,�h�WQ+�!
�9o
�~��vS�yY�vx-����a8����1�V�/��M�D7��Y��Rb�(W�h)m�:�d=���g��D�gQ��\<�h,���
Ǐ��i���2j����1�ײB�T��+L�����9x�T ~a��G�
�}����f��ǂ����1ƹ�����0?��u�����*�xc�Ez����fkq,����Ծ	�̠���v���-�]��
L�L�9����~�Ϋ�)�Zp�՞(8��s���9���MYT0o�r�$[�A����^{��B5������S��EC�!㛹٘��z� 2�v��@9صʳ�٧ߡb��1Sf)�8e���X�O�}��r����O���`vS)n��ojm�]u6�@̺��ێO`c��Y����A%�O5�ܤ�X�HKP3�vQ�s�gWutuh�ࢪ�
[2ls��x��Ğۉ�!^f�48'�&����/)T11|�
�^��[����@���=��h��3��H/c��?�	�x(�\���6҂�1���4T�w�nY�j[9ed�|��֌>�6�/=��ް?K(��)�%�b��۝LM�@ᰍ��X�����94w��bp�v�	�������A����Һ�j�o�f)9��Cz����ćL�Mb��P�%A�Q�����gU����{&m�0�e]I�K������l�w��RI���c���Z��t�ߔ�o�M��F%�P���Ԝ1�j�qP�Ϳ�[0"�C ���h�헒��X|�-���8��70$�aj��,aƌr��s���Ajσ���j�0��LT6��	�
LP`":��C��4��Wġ,"������:�9#���0�/��S�	�#�|����7��#3#�����!�UJ-���h��M>4�q���h���"�UK�T��z�	�!���?�eH�Y�]`�%��k�Y8/���g��>Em��x�� ܟ@�"Գ;������G��快Hh/��&�ֺ`s/��6 *������nRt�J���Sdݿo�פ�^$	O���.1��CG�|�>�O4C�|�|�2T��&��b��tXЅ�m,4�����px�wK��	ұO�W`ű��u�+Q�z����&KQx�B���i �Bb���#}VϥN� f�:~�맲���R�?X��V�:��1�w2&MO�bt��LG�n78���̾��5��N'w���{o�s�3lk�����t�I{?e/g���ЪDp�%�D�}ȉ����-j m}:�|=��i��UJ�?ѿX.gRm����|Q����䣐��Yԗm������V�J-ߥ34xP������jA�H�_�`l�}�����Ը���۸�͍0j�������E�n�c��f��W\ف���A�6h�í��]��0t`%H�ؤ��s�˷'=*C�/�۸%i�t{W��z�*O�n�&&��@d�C��S���0�Y\�rV�3҇=z�5T	$���R�_ܜk�H:�O�?���PF�_�	<UqM�e����)��(O�籙���f��y-���z���"vEL�k? .P��w��ь���n^�7�x�G���n~w���X��vx%o����=6l������m����T�0,C�1;��T#E� �����(��A�x$uIH����R.�hSGJ��B(e�ulrU�%ρ�m�N��i����b�yŘ�$���"܉�W8?����>�=G�x�y��5{P����Gr���86���fL��T&_"���o����<V��Ii7�� $�v��L��<mK�[�#��Nbłd\Rv�U9&��p^s�Q�lX�G�W�R���D����G�D��t������������6e	�4IL�+(�:~1+��9�T4X�IƄ��q��Y�}�ȿ,��sr#���Ȁ3}j-
����(��)l���:\�(E�����5,�Z��B�j5�Jm"�
�	'�B2(����v�a!��=��9����(܍>gfܴ�Ξ�X^Q��_ǹ��ޙP
�؏�;4�|��U�w��D����(��b�AI�c�0�t�_鴠��YI�*	Tm�#+���Zȣ��5d��J�Dң7�H�;���`(Ƒ�%-���!f�ga��|�u�.�����a� �Z��k�z,��[�E�����dB�oژh<8�\T	��l=Wm���2�*�9}v�u�DOD����	/N#iD�JPc]�P����
-iL%E� �~6��&=R>1�����/��Sjn�bS2u��@�T2ͩ��d� d��ob�Di��+w�E�̺T���������ʩðϾ?5F���H�{?�ă"?����]�v�e
~��4o?N�VTq����l� �}D6��z�����%_�@uL�t~�m�5�}�����ӵ������-ͻ3�DH���tg�4�d��ntJ/j�,�@����of@�����I8���rz�H���#P>]z�R�PYSTG����rs!�&�vY�d��р�o%�Wy�G��.}�	�ϫ�˦n�N/��IoY�{�1Va念��w�(�cC�)�)ፆȹ���g���0|A�s��^_�z�iyŐ�� ���[c�=�y������6)�^��n�n�:%�g�ZB�M�h*���M��ƨ�@X��~�*�W^k{�R�P��;&��*�*��]ӹ����G���cS�=�|=I�g�9s�y��m���r�]��ג����8�~baEjA7� �l
��!b����3����RMi���N?�`�5�,���i�m��e�s�w��{*��~;]kQ�+��0�e����1Q"�
�5��"�^�+����VD��R�KP�'���쬪e�r^C|�h�D�Ac�B��3ٿ˫�t���5|Su�Hē(�[$SH������#5�r���Ɣ�6�/��I,�%�#Y����>8}I�"׳.�y~��%� �����r�����CuU\����^�KZ݌��Q�X�d�Փ����|�_�$_OF��X�V�埕�a|���f�L��Y���}� �Y?��U�&g��O�n�Z�w��{jԗ^��5�ܝ�'�����c�����J�pi����+�ޢM1�����2���K��r")U#�ߝ�����o����"h���0��:}�%�e��ł�Iu�Y��['�]a�ʨ6p�,O� ��5U�	?��Í;��p��t9�!�7iٜPF�S��P:�_Js6� s};.����,�b�����U�^�=1~�m��8�QV�
��uk�%�v�9�K�Q*-�)kXr�*;ER��W(�x�*���o���aY����^V�h=��jϋǣ��*��݆[5�\���*H1����%�	z����n9Y�1׎����
�<���22KĠkOl�`����C����d8�d�&�t0�&W1��-U+T:'v����F���#LS"�Ե+��8<e'��y����6,h��7�����{�_gߚ}��j?R/���Wr��,d%��Vsi�m�x�#U���sq�>���N	��2�%�-�w=����k���u��zFy��#���&R���B�JfGu*�����p�a�B�{h�ZRC�t��X	`��&���:�(;%��������^S��z1�DZ�!�(3W6,�5Ғ��gf/����񽒿�xjr:��"��!}2ȿ̂�f"�r�����(�c���LH�Wʂ�j�t�#\�LlY�c�!�����;@���yE?�.k����ͷ�K�F�!��tY����$�վBΞ�/��l0���te`?����s���Q�}b��}��uo�rŜv��5D�2Aԧ�N���OB9V��C����f�U�{0�ip ��a+L=��H2r��N#d��I��-,X�LAV
���*0<�[�w0��"���y;8Y�5�T�����������*#�"-�󂑓�WQ#(��^<��a G���)y7�Tk���������v�2m�,�@ɚ�kI`X�4֧q�Yښ�[�©WB('?�/z%�*������ ��t��kL��3��{;��x�kO�}R%��I"�S���`�Glޥ�^f�(�<V�5�	��Zî�C��mbG��|���ʔ��T�@Q�xxH��x@�f�x��fw������n�?�Ʒ`u���nm�s����p����f��ELx+%��t���E��dN�lT{P�P��a�D�k��J�QR��?p��uH�<5X~�~�u6��K����ݯt�y��z��K�
s�F ���Ͷ�^����,9�|��dz�����k�;y�o���x܇�e3��%!E�`�I���h����m3$���Cmrk�0h*B�Fu<H���'�`���[�F?�����@F.Y��46��dk^h�|�Vw��+��Y�H�Uw0��[�o�E��(CpG�,��C�7�c�*�h�Y�'��	2�%�*�G�b�tS��Ӌ3�=3J���O�f�w}�.��)��.����7��!�.���a���W{^��n�p�� ɖX��ǻ�b#iA��c|:*�W�fR�����Ch���zFV�~L���T�F�*gZ�n�p	�)�7w�P4�������X5+�OQ���PrxK\Cht��j��p��v�A�7���c�t1H�RL��Ԣ�ɗ�JZ�2�O	�S���D��o{�cȢlē�ܷyq|!� ��"��Z?=�#������^{�i.ü���u��0�]X�(i6ap7ˡ�$��"'1���IT�&�R�>��U,a`�O(D����i�D��P���i.5��&�iŭ��z��AArr���˵�4��L+�y��yꉦ�+4���
�.f�1&�l �ʳ��_��il�<��ћ��A&�{�99Z� ��nI#6��{���F�c��X\z��a��bj�����5萂pC7�Ϭ�\&\\}�����+)��.���<��}��v�a��}��@�âtj�H]�ဠ�Ŋ���cм�Ӕ����w�.9#7��Y�i�O~N��n?/a�����b�١�%��Hl�<����B !"�.���ͣ-�~0۵%�r�@���UV)_�*�/yZ1�c5�1J�aI�"$;�	|����NQ���I=�=p�񴅒i&ːQ��
�t�e���ĩ�B�5?�l'Eȹ�.*͘@�#��q�������FP�g�C=G@J�?�D�Ǻ�QN�`��L+^g�鳀���w��.�gS����$H-�H�\��U�1�B��z���ps� Egm�g�/ck����%����z҅�Z|�M �{�{����!ۛP�O�H��^Eg`J�#!�iȀ[�6~�z�	�]�ږS�q�[��*\w�i�mU
�T�!@<��r8����,�h��u�<|�&4��x�ElH�դ��!~J���>U(Mj�^Y�>uB���Y	%^v*,˾J���ơ�ElC�r��X�F9z��O+7�H)������&��L����������L��׊���� ��pOi9��7�)j$&&&$5��vY��D��a��j¨�*T�}F�Q�@ul��I��P��RJ$��T��ӏ������mC#K�~��sN���r�e�c�j^������[�C�׶�t#�N_�J��z�%�l=ٰ4��e��#Ͽp�ʓ������8��` ��컛��@|R=߈C2q��P�/f-�w�6^�p����\C�N���H!X7ܧ���c�� �Z�e�JD<��L�D�{2z��Uo����c����#�6JWM�$��<<�Vu�c�5��O?} �6{_��MO��(v���Y�k��~ά�cA��2�c}�K�%�N�J\xB�F)k.���u-����+d.���Ō�Vb:~G 7��U�x/�x�Fc�a����o������k�Vo�".��dR�z��d"�$y���;�<�C:�yQ���}���Y�~��_,���bL��c�	�ͅg��6�{w�W��J��~s���'Ǥ)�o��*�����]��W?e��3pģ~)��*~�qRyBzB\>.��$�J�K��GR�k蕧@�8_+%�P�����-�ïF]�u�D d�v
}��5�	K p��c�o��J���VM9H�	|i����w2e��̿
K�j��:j��F̋X����FK+�'�:zI� �E��Ź��2|D�#[��h��W�z h��l��Ϗ�W\�9!�V�D�j/�AJ�̠�L�����X{��VE�� s)�+3��V'�>�����4(�P��RUz�$ඪF�]0ci�U�YÖ:�K�km.{�q��`"lï��������øp�*���#|b1���q�[6���6Z*�#�#�e}���1���pV��j�젠O!zR���9C:�	�Mя/�p��{�ܔI��L �K�OB��hs���\�L'k�˃��lŻWo������ �D*�/��T�Y��)�]�z�A|b��\^x q.a�ͧ����~pK���3Z�֟��ݤ�g��$U@���"54OXc��!��f�M躆��w<�!rv�B;���bCݟ�����ڹ�8�l����Bgװ˴x2�n�O�W~�	��E�s�,.iL�i-4 7�SiQ��]I�9�����3.��E�=����� �`j�R)��L*pg�S�Wئm,����-U�0���hKh��4'���A��;�N�FD�(���)^�e�� Y�j���z���Iс�q���a�R�в�:dM��V��i���UTt�nh�+s���G�r�����Y�ْ�ݒޅj�IUƬD�Bk��0JQ*Glo�b��\|Zʪ���� ��C�YӷK�s� tБ��#(+~���>Ы��c��؝�7�iF���;ڇ�L��z�&�E����zD&i*˲u,U�@�!3�kh��H0���h�e[����0��!,}��U�����"�/3�]��2���iQ�'��B�]W�L�oƿV\ad�����3�������ٿ��ձ_�2�������Dɬ�.��>3zA��F�t��o�QdL����C�2�Nc�"�=�6��Ik�$�*r��o���#����!�����m�[��p���υ�L�8�zyKd7���_��,f��E�@�vG��U�Jr��������?�*�G�GL�	�q�D}���[��UM�@4܍�ʶM[�]����|V�2;�ǧ[�t[��ٗ��W�),��:�,��,%V���F���UE�E���`J+��9��B�Sv�X\z��L����A�LL�	����� ��,&��w�팦+�����#����;�,t�u��T�pp�ƹ�4��_�CԢа�1�ˆEV#��HMz@����RbT��k*bf%F��[�k���7h��4ΟY��Y)&���Q��ZF ��8H�o�y 6��w���Qr�A!��?�i�T�/�x=��P�X	Ю9"��5tJT���ZP������/{�/I�mLЏ�����#L�]Xk�[��^���Y�˭�-����������?���[�Do�/���(�rh|E��X湈�\���Z� �w|�@#gɣ�� _�Lb��}ۜ��MشV+�zQ[|��Qba�8(�~,8[Cjd ��wf�c�
��d�)�&d�?<�|������,0���h�C�q9�;zr2D�_o������7��A��j�C���KLa�����ڃ���u�!�b����C�������ӇdT?~��&�"8��'b�7�Cʝ���"eBQ�xYyȎ��3��8QHdr�R!���L�6clm��_s�Z	,�cXJ�l�D�pv)��z�mcH%�|e4�%P�`.-J!�s露mg�n�F�X��SL�\2py$�G���	�z������V$Y���s^��?E��M��gA�����D�c�T*�
�h���`����5��ѽ���v�,uQ�k�ʒ����u�(A{��֏�MD�"j��.D�N<i�2�Y-?���QW�ۇ��Wd�a_���1�F0KJ���:�������;!~\"ݻ�3�5���D�0̈�-��"�(@D�$.D2���k����C׸ՄD��	!�i����Y���)<���,�Qk�l�W���ŧ��8cYN�F-�X�ܵݗH�Q�xq(MA9n�ѥK�>Mì]嚈ػl~ҎEY�O� ��;6��j{4�֪��D+)�~�ȍw����5�xc-G=c��L�&�����@��ߓ2Qv`�e	�T��m�uHM��#�,�A��q`��']ݿՖ4ʞ}�o�$� ȿ����B�6�?Ex�����B��jU�jh:��	w5��)�y��l^��}�*Tz��kH��m���!e� �_������HU�"<�ىZ����~��~;d@��j��L�YĆ�b1��vt4)�oa/8hZ��ʤ8w��+Цh���+�M�|��L�7�)�V���R|��y�쁣t�Ci!٢U�]��h%���'�#�Y�D��Q��3g��w)��
��d�����[	�Q!qȈ+ �.H4p���/&aá�������
���e	��0�1�W�	_�g� 6��ܬ�iݾ]8v��L�U��ɄZ��vS�+�u��<	������R�Ka�l�;2��T���*���7�Yde�~O�j�nӷ�@�}��F�=�Tc��l��<��y`�x��[?bg�>Ϗ��L�w���n��5���������-'��)#�E>Γ��aF�-:c�G���`�4:�X�������]=�~�΃���~�RJx��K@#Qn��B8n����k���O�����)�&�N�P� �a������0ج��0��H-daǻW3ov�\Lm�����'sn�{�:�\cY�i}�B����Q��T�Y?3+��4�/������[�X�A��BV�pJS�"��Ke�����Gd�wۍ-cT����Sv�$<{�bs?2M��8�1��^VGSv���;���r���G��a$�_�#���U�N巜�}��E�rdci���8�>5��ZtAt�r*{M�52|Y���AVF3T�j{���~�LC8���7?\�X97��Ɣ��^n�#�p*`hJr\�W?�h4�,��S. ct�w�cs$�)��~H-i��Y�xH�gy.4�v�6��~�}@�Ӡ?`�!{���fWƼ�t�������z��Vw�L+$$���O��3�H3�a�e����{"��O>)�k��{�|�J�a�4���9ϛ��=w�H�d�:���$����It!�a*��=���
������U���.�{W��x������W\��-����ͦtSǕ�C��4�O�T�H^��ZY�״{}��Q$Q!�S^�t6�����ŀ���l-dc�7��s"�zf_L �2h[���-�I� �Sq�-^�E>e0�C�4�����UMx���9�v3��FAs��T���%�� �ѩ���G�Ů���{ �O
GwT�h?�X�ǘ}�`�8d�q-УF�^�����:��J�o�����*���p1�	P¶[�wh1ע+�^�c/)�W�Z���Y��k���
��"�'����� AkfD��|�ws)���=�������sr�=z�u��&���6us�C/W�bb�O9����u�&#.]`c}&�h�?�sd�F�l��2΀�jx
�_(�h��x��7r]����q��4B'����\Gk+^�Ď��X�n�ٯ�?'�%t�,�/㣁Yl)�>)s%����(�+�G�B��L%0/v���� <�N��s��ej�կ��*y۫�B�`���R5ĕ��׆>9&�P:,k�2�}�ߨ��=\��H�]��� �bQ�c�����5q�
{Q���t���2����Ee&�3�P���5�%�2����Mfk<��6m+os3�0���s;]o�'�@�V��/~���J�0�c�R\