// LDPCencode.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module LDPCencode (
		input  wire       clk_clk,           //   clk.clk
		input  wire       in_startofpacket,  //    in.startofpacket
		input  wire       in_endofpacket,    //      .endofpacket
		input  wire       in_valid,          //      .valid
		output wire       in_ready,          //      .ready
		input  wire [0:0] in_in_data,        //      .in_data
		output wire       out_startofpacket, //   out.startofpacket
		output wire       out_endofpacket,   //      .endofpacket
		output wire       out_valid,         //      .valid
		input  wire       out_ready,         //      .ready
		output wire [0:0] out_out_data,      //      .out_data
		input  wire       reset_reset_n      // reset.reset_n
	);

	LDPCencode_ldpc_0 #(
		.CHANNEL         (1),
		.N               ("1"),
		.RATE            (0),
		.NBCHECKGROUP    (90),
		.NBVARGROUP      (90),
		.BITSPERSYMBOL   (1),
		.LLRPERSYMBOL    (2),
		.SOFTBITS        (3),
		.NB_ITE          (10),
		.PAR             (2),
		.S               (4),
		.ATTENUATION     (1),
		.TRANSMIT_PARITY (0),
		.EXTRALATENCY    (0)
	) ldpc_0 (
		.clk_clk           (clk_clk),           //   clk.clk
		.reset_reset_n     (reset_reset_n),     // reset.reset_n
		.in_startofpacket  (in_startofpacket),  //    in.startofpacket
		.in_endofpacket    (in_endofpacket),    //      .endofpacket
		.in_valid          (in_valid),          //      .valid
		.in_ready          (in_ready),          //      .ready
		.in_in_data        (in_in_data),        //      .in_data
		.out_startofpacket (out_startofpacket), //   out.startofpacket
		.out_endofpacket   (out_endofpacket),   //      .endofpacket
		.out_valid         (out_valid),         //      .valid
		.out_ready         (out_ready),         //      .ready
		.out_out_data      (out_out_data)       //      .out_data
	);

endmodule
