// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:37:12 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nXfP3F5QztkBKOIfGhxT7gZANdiKQJQv5QcLhUOyrE8OF1OqRulpRP9f6jA2SY5U
TVdi4ByNXD/aAC19LosLJkPLhCsQoCwW5lqDVphZMTi7LPG0ua0Ge9QfMTTg+B/W
7+eEJ1NqxDx0qS7zwkXlYRQIB7/+YH7hvBr1lIlY5Mc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 90672)
80yJzN3/5dp3+DwnmtA0GD82pNqgyO9vnRl0zOlfvLe7lr4XrlBSM36Hgx6fUHjc
bqF7f0J8Pnp1YAK8Y7mBLxiGT2ohyrEo4GHPGPXO9PwjYaB0Jury6V1v57s0fG96
bi7lbHrj6r/SAfI1b0nhRjf8lMvcSd0neLTKcEgV9q6/C8itiJY2PTY16VPNnn2u
PeU2ahcHPvIqnjBjUcWdlD6fdbJMDdfFerzW3eTI9lgQKaSbroMRj6gkPyCTVgI3
P6v2CmShnSlB6UdS+Av0psUF2YgYVAdEs/pzH08MgjaQHzyWNKZ/ImfNOlWaoWo/
TgbirS5wvg3X21mKJg1CEq0igEYjsAvPWz4+98m3UdMf/6mfTeKvA4QOmGpIv94V
g+f7MNTcbWuB5GCsOogKLktPomyVI8njj+gRN2NVt1aeQmMOO3UM69Jhw4naESQ7
Iw9UURY1WwVIPqhmKlOi1IQfXdtf4YUjAeKd04DEfvsigRJGRWjzOZt3Qjez6eKG
MTskl0QjlY3Krz2w6vBJPzGGh8rUNwNhq9G1ejKv5K00ZA4mBIC30B2w+7W1Blj8
XIVJ9zGXpkboj0jzXLA0SAiBGigzJCNwH9JpHnxR/ZDRWs01P0HcyIAQvvbgf9jo
gHsqNF4IClPXihh6MOorH2n3VUW3tvyZsHjiN+Y/wzv7cFHoRTop69cMj6Gy08LR
5XEAd2f+UdiE9YP5F31IHXt+wCqT8/cAjZAn5JIcPqhJMRCLUO7lKyLuv1UlDf10
6lZt2UOZL+iA+DhtETn2Crqq1iduIUWi4WMj+/AwXB9+rog3GtWQLY6B96x/cHXV
HX3ENHB9ayd2gIzrmRkRQ9XW6jibqdanb4XnlionvPAfRvQFtV992VY9PumtDl3W
WmCteQjqmhGN3GGdrMYHyl8Kr3eiWL6U2dOeaIflfxDJC0tfSiYx2vy+CIG2S2rc
1RF63cv+kGvgFQ5Dxe/ijuKPPuRcLYGxrCDuu9ba80Tqt8dVLE1KZ5pag8H9qN7W
qye/n9ZefhFHFRb53zQw3B2r/eCv7g+2ylS/U9KmjOEj93JXaHwCgK8oSu7ow5rj
IJDYkiHqDlCaN1fidirlhyc6PeIhwOAjdv5p5kX7A2hK2bAOjWj6tTM3DFQlTLYu
Q3RhQSW9eqAn6sbVGjsLi2Ait1Qscf5VzS9ZTi9RrvfBlkE7GPfvov4zrHZzg/6l
bQM9aUmFmdHhFJ5b0kchX3KGZuwNBYkM11lg4ZapB2COLKpOIzDSdrie9dXu8PHF
MbAI4osiMeW+DOya2v6DE0gX156gep+3nE7Pzz4AjVzn4dZQ7NfKUQFlvpDhA92N
GXkufTuM/SwczwbYigDpZmNdKpZaNQlobwbyikHPtq4PCPGktzI2G29S0PH4KMkb
G14Hglwfs07p/tB3zglvz92ANd5Uciiq0wfkkHu9chAmxXE32leMUysP8R9HWKU/
fSR8dqZ2hswnzgPzGyZZjvVT2rbqRY6wKKApK2iHtGzPRN7VvlYdaKPdXo0UplKU
9roZjPJ+ZgfKgnzucxEcJ0mcSel+KHTUdiF0t7BPRzAqYg28fKnHujXppEitx7Bx
OCdreK25VavDAdOubKUpHZ7nQJ4A0e/LIxa6G/jEoqmhxhpsEjwwtcs/Mkprkv4o
fkzbH1UJtAKIHWu6lLgZj55TPHdlopn4ZAVSQi/ujDsZMiFxA8DRKn/TTTOz/kQ3
U6sasDgOtXBooQxY8/7qZE04037HYdKi9+rU8JyoBGt2uqJ/3YyeCJFFllfYQ/bI
hzEhGP69y/pu8g6r92aZTvbyUV37urcnngYxe9DOZRRwvgdDUOPtn0g15zchK11q
MjwrpA7KROxIlOMwI1aUf0nlNvL2rExrFLrTmBA5sRRd+QrJhXQubMDidRffNbNG
cIiW1O22Zslsn1VXjkGKw4dgj450BTfWu/udvUyFL4gA2Mi+0tGi7es86ZvZqJUJ
ZNvwQO+zGBN8KrD6Bq5RB9y/E2SJpdtjvUgnbMoCJU+kdXJsoSn/Te+EoQHZpVSX
F50P++aANZfJJ3VNglACQVJQGJrWatu/TuZHqyHdGPc7rA6JYK2pgX/QmMA65yF4
SuKeB4ui3LSxGMpyS9b2cu6AK2O895wyzuyzv2bKT8J850aKAGwWKF8M1Lmym+ra
zrH/7r5Xkz5tCFAu9hIDkP9wlnJV85kxu6M/B8RXvbldE80aWwj9vuRfLn3ttHbv
v3bNDMIlLrf7221H/qRQ+ZmsDGJK8cX1qjLPuRIjPB3vo4ue/ErybDPTig+r5WR+
HMZ/3xL/yhO1QrAegerxW+3dwyIRppJ3YgiLbqmrjM9fPVlbAGsjhvu+nrZ4F7cf
cfUxw0glznKf/uXSwvaSJ/cVh7yfyw67++pNiknP3p7FVOGOGitYiETUD9YoOX+s
w4/TDYQYRVTOuxQUTNAdC9ONjdAILz8YYpZ7KnP3L4uD0Ep/iFubaNXGfLywUgRN
jYsY5EPluLXuTjGZyjVmBJwVTmdOBccKcAxX/OuQTLhAmxlUVOE2+hFBomzeUnGy
pfK7LNdWkzi9a0BJEcBkGKxgoVZeSEfo2uN0cBI2PzXpR8zGDomi92ifKYcpVH9e
S0vNa8xWOBWfjTtPOFut6eq599+8EhoMZjuJ5YlSgdPLMBTjKlJRpwL82If3Idk5
P0iDwX6YjG+IlGd+vKsphh5quCIXfJcZM5HvvNUEcevC3/+D6BEKf+H2vOkvjZ6e
tnG9HJp69uVZMe1LvjpHne9Xo6hokfBQIBPCcJjh4K5GcXhFbTbkZ/U6kzDmVTR9
QxgVvnaHtISBENLo8IgmRou1AC1Y+PszhhkYfznbuEi7VNZ91lnWNvc/2KF5Dr+M
uvxeqBYdeTFHNXEpgkzd0FXb+hSKqqL6tmE98yXB7vJjMoKD83YYybfDCloCccv8
ovW1Eju1JTr2h//aZUEx0bWyGxjKm2ANrFCKZ60HpB0FMCU2J0d4tkPEz5ft6sZ1
oKUy29j/hDtQjMqk0PCKmEL834sX1uhYHPk4i3l13rPfxA3brSHPLhJS1XTxbUkf
Fso9uA/ZtgrYR8NXYECQIuti5BlP6g1zxyRpSMB+84i4VwOB674HBaM4R0o9nDAs
bI2lNOHwy/poxa784tkVDAzfowm2gT9kHrRr+I9rw2UjCwMgxuXE/XBEna1goeMv
E3+ayvjQaECwZsAtofgL4wQ8Bdqxm7HOsCrsBRa4oRGDNb2gLoL47piaoRIlrucK
khqS64qwjy4L+fqQGPbtVpaX8UHil903SHTpgMgzJssaIZoSVJVYy1sxhD1qX0Pr
tkNh9GAIWEqWrl8mP14MHynMrlw0KyWJwR+wYUU/9Moj0cRiLyyH9C7VnPl9HBSw
4YEQFe0Au7h8t8ZAO+3SO95KxQHbslKDdfXlyK/tCL8YJKwX4clpftO/wxPp6NVy
4ZXYp5QspCUl3MzSjldT2+SQiNO/Bavotui6RQXXWE7Sy01hKdzTc33X1op8XOWT
YEFkNxvbWP0U+LXj7mX531V70u/gEOH7c/EQjzfN7DINf0bK1bR4lH/Le7VCtbo+
q95RAHvY8x23ZgUjPlcHK44ooXLLIMMxug18GUJs3UW25hmHDP4vIRmfQ5xdGXCt
OB8HOo4JQy0G+VPb6V2aishbyVYRP3f+l5IoSMWH7qokgwIAfjNSmmWuhIPIdu2v
Yx8RNZkFWdIX5zhKSjVUdvJB5MTyS2EyJ589Q9IaXkTvl6sgCsSRVchH5AplI1HC
zC2hUVOc3J5UEyf/I8HRw8Hqq2IushW4EYV9PNX+Vae4OKGAs3f28lNYz2Stav0L
ztdQ+5WavCpwDEH8KZnxXqGPwLLiiTszrs46z/ooJu3FK/fUH7O0qJ+nzXVgbXIP
Uv8zuaDSQsWSgRm+H76o0yExqp8q7QOSbrS+zxdaDHOPVIY8XTojKw2Mo+/DOxLu
u1tVpYPQMAcDlo4HHY9CawKGeV/Lge9MrfbtXDSU9dPZFyDaAe5h7R4jTj6Gf44E
UAgMXL/KY4vjlnYof0x4O2EvF72UB/UjYCKFxOSPKdwRCg82i6Pz6TWI8nXzXFhQ
v4SVzDh/TNDCEpaDRtx9FsLQHoaGkw85L8iX9c/blMPD8fzWskT2Z9zOUfDhVujB
bOxqc/REFiZgdPiFNKMYuiRdObCL3YzPpTOo7Dg7D/7zutftMHFi1VeNjQecQJ9k
P2X96sUbI2/AQZ7LRstMDPkG4eoU2JL+vr1XJ6DKvE2xtXMbSRKnQ70xk6wjirWz
7666vBh1dhW7Oie4W36cVp3mElvl5yfcXlpzbDIUaCglwENsemL07fMQ7NkBUCQ7
2+xN7CoyHCYuNl4Xk6GgAEWgIBwkwyQQRb8pFbCsUx+ntyTci0V/BGrvgHn3zh8l
/O3D/tHGT61WBPdcIrDkFDpQeB/HeYaGLRmSgVOSfIdnnITAYJXSC1F/65OlzFaD
y+A5NwXwyQet9O4D7AINo5aLFdinqwTKyKddBWD6h+IxQzArtE6nmumkCqHXqlkR
/wbWowwy+MQANhcrBIDCgGdauSlURK6t59tzJT197Bnu7WHEwDiIlmO0QMbIN8ND
olJ6ZEvvIrYb+OEEhxek4JMDQMCu9W7KhU6UOwGP4MdfxSUfFtgmYAz9kGzfPceg
c9ttCybAi1aNMB49/t9AtFpaNYyU+D14urmI1h4hyEGeWltFm5liyn6YSJBcSqQb
lWDKC4xHDISZcEqaOy7+b8miixoGuCXN/dcegpHLSQZbz/2yixCtfuSXkLPiQtGf
/9T4dh7LRWzBec6qPftsI1zBKr0XiuPxLbJ//h35ZNg7rpEWJJqKasE/BysmmGfI
4jDwyLk7j3H1pjXOQEMj2q90Swc1DU7mGSEUswKSsf9C5uWAXg3nx+tnmgi3WY2R
Rb0kDVXK2TbEvBrAte/5FEtjBtrqbbBFpu0a8qjihwZ+PpG1ezoo+ddZCScVI9g3
ubgRmS2EVaUmai3AZZa0QvgO77MeY7Sm07zazd7HBcO1LXQCMtbee1JQynBQLvJV
YnkENWS+h8ZeWuEnNXWVukW8QmzSZhZU9hT4GQfLtQ0sPhrT1qboBiosqbGTBnlS
t/ss7UQyoyYBnI3VNuYgQwFsMQyjXjRQjIeQEA5hOZt65UaRIKQFYNEglJIb4h0f
z/ZZBJ1x6QRFkDzmBXvthAdYkNywjQVKGmAJCUonE47/wYx9r7FE62wKF1N3QBUL
7njx9JiQ5xmMGwslxNC9Yk34LVEVGUDbJDtQ7uSaQHHgRORzwRPBqHxBuoZ46OV7
bxnWNrJROXlGxwSAsa2OoEtlPsHgqW+LQsegkHoEacLJrMzPC/0YvxbW7qJH9Xz2
ZrPsTlE4sOyT/1MtrVT6H8t7pPz4KTgxG7cDN98eR2XjB24fyf2jCPVo8fkpd4Ot
eFMWQ56kkTYp0KsnfPW+lM6wmo8MsEUFob+MBGp1tR81L0qMU5Zh/rZ5eK38CI7b
itFmmM/Skr3cDRL49YXrgBz39UpQCjC9hkOKjv9IhqkQlwtU4CNfwOJWHIwK3glT
5+xcdbrd3KxjUFRP06EzVld7X+GLLXn262VVddc/G+88UO/p9ECBdHAUqhJlDJpv
KGxRgmWaGvLxVl0jC+tnlDuHp6VpDdIMxVzMbGmqAkP+oBsU1lkLDXHZuCDc7VAu
ye7MzVSn/LMbiqLnkeXH2KXL7VNcnJwIVCQkxzGx9WYvoeW/cWPkQOanr+NuRG8h
Y2wyrKQe+a/t7d9ba2nFpukI1Miz25sKM2eMjewghKAkK/qoo03Y1E/jS/NQXIFL
JynLW3TtFkEOsKJMArEYFqRGLEHV83UHAmeSvkwxD1t2iteMj7hAZnNXYIRn7ILn
bNySBkNFincMNdr+oaCbVwxotg1s+KWG4UoQgAl9xv+8xJ/c2qmh69MMU6yR7mUA
0LM/fBfysa6qyf5boh6uiuL+HyswSVb4pDJdZ1GawtSax1XhTrI2bpV176NEk+y8
Vf6H18BQO2/vcoVR5may6V22eGtW6ihgIRr5yjYAaqzZwTmoS69ah24Q3pDaJACX
VTwf4mhJX1PhowWB1ceIU4FEEaWwpuM/TCLLiSaB5ZintGU+whe3US3M6Qc9cf7b
6fazOvREh+fZW2XKfj6VaghF8JJVDkwtfFp7T248OhX0tZ82yNjH/ExAdndbt6Mv
m1Mhc3eyjPQH6rbH+gbKfqIF1vnoVOPzGFLTZWPxuiEO+7d+4O8kbGGnF/Wjyazo
pQTaxbUzPWSNNA/YmDxYf3AcOxRzO7mfNlZpGeUb/l3YIzTCCNaKAC1pTBFBLHyO
0zlpy8JYAMFJnoP4NopDTT0M3sQgWfJd7TeX2U+gZRAiyHbS9tCsQVh33w6Vpfvv
nIgduujvawoR4jJH6K1qs9K/aHWm35z2Pi+SHEjNrnOaqgHxy/shjtzmJ1h+MKCQ
wGM1UZd8jNDVP+P3n71xjDZMTagIf1gxGpvIQT0wl/yX2WHI6hy7EM14mNIc3hBJ
f/vu3PLRU4iL92EapmZlvuXx0/saRIw9bNqUfVkQH5szZIlG1YZGytVeo5DskgZY
ti3PfB+dyOQWMJvy9h6sA8aVSvFc7amlnBC7vH0c1r+bLpyH75Chlq3IbId/2zxn
ms+qj667oyBle5DRH1Zb7nt5OCGFDC5ov0UxYR8C3n7M8PTiiXhYtZD5v2Z6NWhz
Vag9gQsltBNIBqELIdkbXu33DST7xPGVETvPV4YYgxq13qzgt/HZnPSPPO0YyfKv
ajUDgNnzqM25EgEk9j+fNKbWGcUJiGSzyG15TN9Fag2IqiD0+eWwDNBSsGZ/foND
grZKYoHNMY2xKONdeOp++x8+0OBr/94wd18md067np2LVWaZmHUIQ5oZ0qSbPxAt
hL19m7+tp+3mNOAHHnUak351fIZaO8IUSHiI6mDj/FDRCvi1uMw9+aBRS9SX8keR
gY7u2Tl2geytTqjsIhWCgqt+OGzffbfCpz+dTtFIi4Yl7lTySdk56WoMpCVf2jTK
13lIF/UpLf/C/x1lkxWWfr13neKL3+H+yzJuaEn5wIQjoxdLPbuRGTBilYfArpr4
bzrujB6ZxgJMcEon3YLT4R1C+v05rryAVlkSEg5QOmRx+A4QeOxaqFyCFkpcQMT+
7+O67iMx7HGfGK1Z95hA/eC0JLBNAVoMK2+66kKvQdbukrjHAKkGk4GHdmllCrOi
jt1HxGLHvPdwUk1fkmDxtjsN7VRKQaZYlvIrckVAUFXZMvN6UK0cWgNjTCksLMbc
xPjiXhCxtECUF7elQOhOAEwTYq5SJ9JO/V1pNtWmqNMTXmbqjvaJdQgL0Dbii4iQ
DqulRqpXUg5DMwb+sLiLNh5fEpYdMQegTVVRIwVu05Cfvbb1u4jU/gtdVXUbHcp2
2RLr8qvcs4+AZuou0E/oOfismIoFy4RwLc9kcfVO2pJth8vmq7PvReIfjv6rX7KG
sdw6JEbG+M0SJWvJzbvuq2Bsi4KdVXCGEcYxePBsi1INmEXmAGihPLuPETCC1ume
dIh0PIR3oUBFHEN99Q91n6En6AUnVd7cDkEGMGLHIiYepQMjNVk/9PU4ZlE57Cjd
bJpm19ZCgWXe/+OM/CY2Kcwk9iaQJPYsyX83V5fQ+ibDSRPpVvPdtdtut+B6f1Rd
ijBXkIH8C4mgUw8TMIlZBXqaCcYFxRqFKmy2fZ5BR7bAwVAQbhuAyC9Nazxzh6g8
7d9KFpoXzwNKObWGYa6DTmVz3/mYF2idoBGKxKkvr61EgNOxIbt7P7z8YqothEL3
WKiRo7+vSV25Wt1XQiaUYKTLABXDU7GK9gGT9eNEtDvjYcx58GLgIbb5ATiZgQVQ
lTjw5B3BooU7q0ffJvyV+XdjSpxT6Y1rMk9j5cF4m6Th9C5k1KZeocIsi7uMvj1m
MOf3OGlMHjyZQ5q5kap2HLB9lcO5fgR7LCcxqluLVq0Ad6lFOw3lsW3Wduxjfg4y
/4/lruzUXL7/lSwT4HduWRIDfL0ESH6aBHyotqkTIFlALDT7buXpdIxLw4wmAE+3
970l5Nz1cYzqP2tn4ZcRc0e68vUawbyKMozUWDUtIQ849m7zQM1F/FFKoXvp1lB5
uYhV4+RJv9sHeKeYjpOW3jajdwON3/eFy/Kf0mTPInR/Ky+nVGR9EqmXVIZdqhzB
4cAC2DhJzMxoVzxwpIArGtMey74XnBiGdaAWMHNzQjIIfn1al0CCcxHgxaRoZIOp
U0YSHFkahbqr3ht6VHY2vtOmkkXqEOoFrgoz/aj8pU1Pn7YjO7ZkVHw6QYdwWh9f
ihRloZqTwOYjZ1h2gfEr2AoBCsMf2l/hOtFE4DMiFbvU+J1iH1RACNwNdaDEjDYj
5ckBXhdfYBJ1joioN9uZJzmYZqU/YR7JpgJxynMIa+Z8v00NrM+snl9VzsvpdMk8
1AJ6mlB7BIHpR9tVnvooqUagkxrd0jM8grA9hoV6k5I351Tg5JVmTHqxVXDtv8nf
OaG9G1Xn36ADCsWKn0O263cE7VurBnfB/LUdnrCyPJqyKlrnq2CIaKXgiwWHALP8
3u45anVJ16u/FLSLDgtow4da2BdB6E+M6Il/M6p57gntQukFTSrpvoAIODBe2E7N
7JDb1chyR2AQqbGAEuXnbB/7YxI9S46vT8DbewP0OjNqbWHywjReIDr6T5n9N6jx
AO+b3Zkzsq1qIef2GQZcO40ZuCsOEhzXn4eQ2vq9B+xTuvWRN68VDUpFu2NEvZ/u
CI2weI139fRyghc6K2F3yLdz+iS8Yr8cjVBCFcs/H67s2ZlbsJuEwm3x4mdXfNVM
A2jTV2htKeuGt0CparWda0RghMzQfrbHyV25hp2/AGYHkeWyLFyTXmS6hUYPeIdc
h4jLKlhr+/rO5mtSrPNM+a13Q+6ZlbrWdZ+ElLtuoHwZ6CVqfuV8Ibp6KXFSeIM5
YY5x+OBk6KqyKVWSd6GRQqdQ7dlnX45y8Qagwn4P0fYY1OifiODjbkzM0oXfpPN7
1hPVEKyu3ZxrpCwmdabINvz+bqKoj8FIXa1RMej5LOCi5zu5+fLOuVMymi2GSq2k
Jhb+QB7afir4+U+lvBMntHeK4N81GGCNGu96crHkxsua1dO8oLHJsA+AwKe0V9Oo
7kuM5aquzJxuoWrcanIqMsr2tAm/n/m3EuqjR9okcGDUuk2P90o8r7Q1N1/71PtT
7vQXQrVToJpLPu9l+dNKWirMCB1Shzy56KJ88S62jyeCA4D2soy006d/+ZNeGEgS
7QH4UswepJWySpffN1eQcPnwHRDtx9N3dBZ5Oz0tmyupTEcAcZ83yEyXPU7mb08+
F4RtQOOzwbuhisuOgX8NbsBbOTi8yPgmG/vZ6TU4mCe4tQ3hns8xqMl3SQwa5zCM
5kISX6pH/HUpOLc6Npqp66+v64FdIi7w+PnqufDXUKXbLhEb+8+tMvkK4/gPzC7n
c73ny4+Z+/c/tgltvge1LzJ+alo/XX01u8znz06P6JVr+OuNlJbzfzH2fIHgZtGk
vmrp6un2ds0mAtp7PrVazEV8mFh3BxdlOyevWfM31y6DzZAi5imYsyt7ajohXYI8
wo4ajFfEVJjtpLeLuoPfUYijWXsNqVtNBwiDiltYMIledfC2nasYgQeto6XioVia
t1ESvk4bMvDOnjfZyiq3UOx96mNGnUhk8YjuldfcdfBxBRvS4f7ZPkLNTebb/ETM
fQNH4qRwLirmwfDSYNjl5qvmF6fj00sikhXCADrldZmBTUypGQjz/0KcDYzZ4tNh
99dxNwcDfbuMC2jfv8YdApWXLkwkoBX8ykaGFgNTd+AstNcwhFUF32WjiiikZH2D
NpUX4f+3KerpU9caPmP+0hSDgmm6bIYTxMERgnEyBxhubq3bVfn3RIaWXOI461Sm
ysDi8WJKs7LAn7Rrh2lImdxD1VFAjbaoudGYmogPOipChPL94pNz3nXLsTpJ7RXq
QSfcTDnsXXNQR7hdjMg80NvOoJaTWDD0OXRAISgq/LRV4ueiLTCtlOWWhxdww9QK
FOsuRdyGBPna497MYEoHNKsSEb7J6FAm8KxGx9MfaSbF45Pp4v1SiWXjsDYJN3rg
IzQg+zp5K3SMp8tL3Yb2vF2ez4G9IfIDaOvV7oaMy2LcXSYGAkud4MQqK4CmB/hy
NLUulmgiyyY56NppKKcWfwnZjmhWXfh5VZcwlIWxLMZMIxzFu7oIEOYp9Iq2CWVC
SajW9mhtD2RoyFDfQiuHcEulWf44VVIkJo54mC+ZBU++35LNXTvdCDUeCMFmTlFU
pTB5ZuSJJf9Ptbwzd4oTsefkV0T6lYgkZdKAVhbUypNuw2m/vfojuWrKD6v7ugr7
/y8xXcJzohg8XBCtzYXClh4kNxtdGdgrM/5KVP9bFmSG8zP+vatLWjozKr4aSjpn
pVuJaJZ+rcSmhGnYfNrPKLFJa55jCwYDZciTrgcKgbXMRO/XqIzQjLvvYj5P/lIo
Wr5amW/eCrLqgdQLtqeT+LRA4SnDXjwjBx3VJ8x0AP4XMY4M5zzQaDym2/mPq8Lk
08HsCET0ae0u1K8Rd4VGO3yAV4LHaSNJPqj2cgzZ9HkZk5tOKvb/cLKpW7cyf03V
bJbqnSyBkStMVESYe8WBKW5Vkr3x7I+ux4epq8KRxoggRREVoNfokK5LdGOW9USt
HDlsXf8r+lY299wZW1KhoPr9LFiUIcRFecvc2oZVWcM3TChU0ae327XVhFSJ9SGu
x8VDW6/8d+FGGYEk6r3EExi7VKAi3zrW4UJ+UDN1O8zidqavRcPVsAE88tyBvSG6
vTFT2q0xm3VzVhgw/F4IeJBA45BfWO0YMi2Eeqw+/bgpKert0R+f4+E6VSGp5ck0
iP8kjbPSYzfeKwcvBneF7IMammdvbfQczmjU2ulZ8xTM7S4RP3GtKhrqwahtUKhj
gdfmRkLGpsYMekD6OPOpoGjI7y+agMGeK6PmQ0Aj41sWgzTz4i30jBaeUqkGrEoN
PN/gCCxVe/pIg647yIRPxlKfZVySx60gBL8lAb0uaKUD9EO/3vr+9sAC5I6E1wo7
Utys74yLlj5peBnxxicgIunZKVDiK4c1MvZx7l/qX309aBSBCJki27XsZbKSkXjX
x309SiAjMOoSYJJ+vIDPx90c5AgSuq9bQMVF90vFba0PPO35G7TeCGeYwfwrm8+W
oboXKa5z2mdlWInz4U3mCPe3E6LAhOUQ6SAdPUVXcrnWeikLl7Z6mB6Zzb8XNooD
t4OnRDNquJfOXiAlMcpK59ufvSAD8YH63walm4PQT579MX/9Lx+z/2rNOVQwp+L8
f35NEhqEU+4BrxAP8uqgg5/tXE5Mlc6f4T3W4rbjYr7V1TASIq0yvmJ8B9YfpyxG
7ghitK1B/QX9KP0v62R8KHUA9JcJtwjMakUSvdQgtTB/JuTwKLu1oo15D0DHGezV
t6ggeZ1DtLIEXe8v/7XbpntVp2QM1IqLVPVHnzehjyA1j4MjBnXCGw6WhPoJFEDL
zOvLl678Y1mnaBqxSdFI145SHXHFoJclDmLvmQpxW2tbyPgPWRtcd+mqePIqSK9v
j02OalvGAqkQqfUI1FCNTQHToo/gqyjVwHkfIEzC4qPHSKnp5nwBU3ZqigPu9Yrl
Grxn3ukNBAYIOmOrIF0I6F/kFzAyXxPglwW7FAGvoK2EqqgnD/VV66uxmTY/0JA8
p3ZDpJBzIRCBvirjsYWTGHeK9i1g5efcPIXNSedojnDumii6P6pn7w7cZ8bzdPhX
H3eiG0KS94ACZ0oZosEnR62BJ10zLrokz1v5PL90qG38V6LPVhnf9jaqtqqKn2Mv
Avrn0jYAzHTwcEtWdmYyfRHk0CWcPdK0M4M6VebH0i1/kyApdDoPFKy4chrM06x8
QlId+eZwUylcxp95SbBKuqDMac4pVGt0X4bLWRoxQhImzaiwtLZ9wtvaxFxGpB0F
lFAPvKCG7OGNxJw+hN8eLiN48Fp3LlitdlLzdwt6M+J0Yct2DBSj8V1VMsbR/Ry1
Z6ESJ8IJ+IOG7YKGpoPY0Pji7gL0i/9hoi91wpD/nYjqYviaCTJPsAJe2s6Xhh6F
SLIafloMOcbmidGlzwPv81aPq5BJwtIWMg3po7aj7DHWBK3HDj30sV8aPF3yXTXi
pIELN+VBkE2tRSw7P4thQmzJinpVeI9kws8sjhObLnuRVaCz+P7PclODTHTHwSzp
Vz5o6Kbu8v7FoCj1E7AsUH1vQVijuQ7F6Jw3Gd637E4f0lUhWYDCtCmYBO1IJI1C
bIoneyhhyvZktmklGsZPAAy4CVv1V0ZrfqNgf9KHU6CMoW5eRPxLm+74wSed8v95
xysUqRDUflEZRGddxAIpWGVj5rpbRaSZtCxmySPobQZFbWs4bFrAg0IvL7MX6abK
jhIMHG5Qi3C9FjPPgLyXrhqV0bdlBvpB59SFfDX3DFpv9Sq9QOVvYSv/8lv3U3/v
4gUg3deE4gDXYflLnm57mSg84fGNtt/1f2+FuKKZ1s4PA2O8/0yR1j0lMLJylg+a
YLWJBv7JGOi2EI/e9lo/F+SD/JTZnHTbtJzqT+GZFc5+71a9RDutDNML6DVRqKrJ
rdZCLmqXG3f1EhY7OSXfNKjBnh1QmWah/o6sKDiqW6hwKW1bnky8qwJkgSLdb/9g
B8w7dKTdXZw4tqqRRNMmEe3SfKofmlAD4JQCmRgaWAErUG34be8ebWNHT5wvDwvo
PT0w5H4xYFXdA+PupPO+rOKIDiEETt0KSP935H/JurJAsMIX4lEyIBfiKvW4oUtr
lECeQaLFf3UReEzv/VUriXywAM/HLA6c9Tnf4F1m0ttsAcBt2x39bjLccYe99ea5
IkxscW5vShP62KURnk9MxdUX25dvVeb9Y0Pbit29nlHBLIkZbxLfeQWUSj7+vgV5
lcDzPbrPO7rFNR8TRF8tA61rcvKdoVChD3RgyXxd3ug42V1QKryOYF6zrilR4uCI
8xl+qI7eQWeYx5QWDOr1MheR29k0eiwtDNbBxH4HO/r93GAi5K1tXvEBsB4VFXHj
h1MdtRmKPKFuXFH3EP9N2yexoV+rfeRuJLp90QujbfXAVGUfsDQ/KGCjV9tXK0zr
I0oqHI/Lju98bxT5qY22R2buOyPC+PpIDaG4I1LNKr4ix1c49kLdEd0hj3v8fQv1
GCmsCiZER1XHV3LEzV55LoR9kZ5EmMRXZLeqnYMK/UexE9Ef0SvagJVqh+5LRU9T
nYbEYzJEADoVtSlkBWlW+y03ZEYSZWdCmXBCMwavHx62WZhl1xFBn7LmSZO+Tues
hiYZCQtucn82UMgnj0ezxvHOD7FMew969AzIFQpgUqhL97rY3Vg8NbdraZ/zdS83
2737qT/jCSDX68JbJLPSI2kU5LI5cHycFho4UDmV5O5QMVHqhDLpUr/+/WWYneUx
s7rubTQX9PUgGjQaUyhJC3PK8y4e6v8m2xIgYQP0MHCZTYsdC6b9t0+m8UYwClh2
cije4OLem7MrraY7WZgeNQHmHsnIy/HRn0aNa+vadtEjo4o81f3D7gqUWE17BjHY
bR0uizlPxz+kE2+q7G2QSR+crcVxehnk/umuGaYgPeM2rBYyjJ2To6HexJeNtJLO
dmA/tG0P2NQhVFL3qfhophocWx6/48GNnGVvQp9GmLyYi+c70bdFUbzDcLGvroTY
UAiYT9+HDnTyf+cKzE8ThfM+kiX5cpaS6Tc25haSghGZSIZnQz4uLboe80q793h1
45U9IqgjIx3OrJJy9383jVJ5xCSWr1P6rwPOUFX4E04LeYwo2LQaZNhDHm1Rlndx
E8hjQpYtA5r1AVySEe+Zhrek6x5zrGen1gSYbUpOeTQrvVfXTwANO9Thrkh9k9Fv
x0xsh6gbzqJqiqliRurtVWA3ftUEWRuKgC4ddMBqwNoP4F9DGtgRSJG+q7Q03Qks
8zVfrF/cNvCqqP08wFjRjfZRfuWv1VwvzouO+LA+zf/mvjQD8aHfKYlXlzcu8vhU
Z5vNuTnnDggGV2E1XAtcAHN2OSu/Mcs6brbzGuG341p1ObWYmakp551nb501k2xQ
Iph6NteEKsR5oGBAsPvIVIOMrJ1QfGEYt03IW7JJ/lq1eQxbcRFdNb5UOVqFfxjl
KjGx+4OVLhgETRVvo8qK+EQ9E0ocwyu0beGVZi4bbiEdXpxJtJLeJIsfi3ferRGL
MbfauKkZmIjwqYOargnfZwYAne1Sd5vVn7+pHQsgvDUAwUMglzXqg2jiTAAQRGwp
Xom3Flf2KRAtgeN3BQdXTdmZCg7DVle6bbJCdR+Uf5dOZ3SfVekwr82JUfRBeGdT
8npHSKdig5tjUPbRyzQa9Vj2VOQc1By/mH7AS056nFHxDc13euX/D0eO1/eBaf6G
zdKjkjivSVvwUPFcgeoA2bxX9PmZIcKbigYYFy/ZtFSt1Xez8aWjYvjQLS011dCt
QuhOX5HGDaTJIMkyBJhwXVnfz8/ERE+tw5aE5D5rBKRV3OsSHi0fURIO1HuzS54z
IQinwVRfncDNqqnadpHpBHFkJDFWMdDYUUVH1W41dR0UHN4GZr3mwyIA2JQAXVxo
EGzslytQqUzUJxvkkIPXlVjSXAF5L5cPouKgIZTAD3dD/4uhIQYZnXs2mhXB2Vl8
/J/FJ9K7iVYMjEY4qQoFVSmHOYwveYuFRrTAkvKILDnebNxwdCEX+T3N6r6H+FnT
LHoSu+Qmfb2FMhz0WRgR3LXt1woQhxdT9H2bTvTLCdsiTvyLQxuzOpAujEuj2QjV
dl6nPKIeTkVJ9sRZuCOGbaC8dYf8jULKRMHBGBjTRgl75SHl5ZNRn0Hm1GEuQGR+
T0aBWRol4pKm8SmgK3Yuw7U5UTlko45zLpbPeYUKvPOSLhufzwMoS7vYZP/mM5Vy
r5GZPvE9tLq2Q+Vb5vQsEhRRRHb+qZKIOGezb3frYdOtuDdXHTF96G+KQdeXCU3K
pR9Y3pU/V98VuiMwkcir9LIwc8GIyH18ylbovJr+GTMqQNcE8gF77DdyOMpCYBeZ
XMktCCoHA7CqQBB6uQwZ2fWGijwxoM1322paw2KJq2lz33vKYFUE/Hvz9Iy+tilB
iQQ7w0A36UDaKshqBADH7p31MKw5Z5RYUccPvuwB5IBQtaUnwoo92X5/PJldF8el
R01BlTtXS79vtP1h/1x0xjOiPd+cfApBgeccEbkXOg9C0/zFDNjwzP9vQFust4Jq
Ugn1ESxQZQxho5heb3CkUl8oYSQsi9Coh+ajiqUiTxhltfkxpoMBAbt5bQc9897L
XSxXeGHOEQ1KsAfjU9HGShFWlW9duvi9M/8NhZjPjnxIcsIB1a15ecFhxY0nN4x8
vX/zCO4BkzdTG+j05pJy+2p1APOihsr3MA8+/iuyKIsjyWAbtVo5lX1FolxXpJdD
mkM9Siyf9YYbxyCzTa1s720UaVtNS7n8a5sSi+OuX80+js/UosABnBJs94TqBDNg
x5Oiu5XhRugs3xPhQDetnc87P6iBco4Brf8fuFSf/Ac/MAG+DiscZ8ZYO0+hi/NC
9vJN9G4S2XS025O6nqm3hjF1aMH8Efi6ZgzUkbYkSYJgeER83A1GzqCuzLThE/y/
q6g9yQWDqEQnuYFVuBa9Je8V+0iPb4GSvZYeSQrfuU5JVrsFUtgZ7c3d7BgXpqZu
cVo5BKB0SNlYo7+iI9R5pPih9pMy6NfdFFKycfage9FLsFPGU1vcxbh9gH+1Gpos
ikgMTGkBjBSe71vzvE/eKw/tDWd9EuEkrweZZYI5swrfnYMOb7Bh0WIdVazVXtMW
GYFZZoYU79mLpYGBZQGNQTUhaazTUtSCwuMdXpczAtdLVLdJCX/Dagr+Gbts1wRN
gRtsqWUpUh4nImk9GDTwGEDzhpFdL+ZqSD0yaDdCmK844i5+fGgmmc1hdO9gEJje
Oau7AHJPG1+p66vSkugq9vS09SOAb9Aw2aGoHeK+Fre88BzlKojniAGlQu3Y8D+9
wvUjd3NdlK0BTvehsjeYgVawooR7BwzuWruarrpTL2yBFrkpLraSx0hxYdbwm6L+
Akd7SgQmhMVF/n+oFbFamJjs6mbpjumZ01wSbSjIJKz3vm1IOlzWZhNOGl9Dvev/
KIzY4SQTb8cfkKTyb5iWVyGPCcE26DkHwBIQE6u6Vd7nbKyzF/DAS1TAlsTkpG6d
IkAb+7s1FSjFVqGQ/AWYRqm3llDfDuqFjeRsuGZkbvJ1LKV5FPr0iRGe2ZhjA3/c
pay/aDEBpED6NCD6avDy6fL3hoysilyFcmsQxhfKs63LSWOb7K5iLnraBLOEdT55
d5+iYJnjUseFHGFX1GazriecG03EmvVnvsAmPT6lpsJcqUUNY3ebriTBDbLkdpMh
iMMIklOjQg35nN1nD+ZEdbaRnSQo6qc/VHDU3YExCOi+BehMQ53yfdLkXvPzRi6S
oQix5QJA7Eiwx9hEyNsemrpkcpPWXJcDjtqWrGnuWgy3QFku5qKSa9ZovXZPt3Ut
E4cc5gcP86rc55D6DXsfHHmzUCm23ccqVgahgQ0Zk2c6UzmLU1DsAtKjC0sMC/ti
0hMtjikVGZOOfvwmfTo3AngiNNBKaiprCLl42Z0w3S3x5jEFAG4AvvktjRI+Q0oh
e79NWhJL7M4J6Ib6sXxOSxS3RW7ZEN2VI+ZQumnhaXhuLlcAuY0BDxWcMAYwbAui
Gx5eYIdk8E5vFznaIPozOJJAYumTZcS/kvutJ1wn5JqyiA4H/2mxN/wXeOBHNbK5
aQQ8/vZEAejyeK/Ic9hLkQOPTUvW1BWXVdvxhyFntRMo8GlPkfMkR7UVh8ReAuQz
XflKzQROUao7SHL/dPMVudATJMHHib2h7g4CmqnjqmTlyyT1rBmomI5cxpaA19J9
i3yO42Qmcw6o8U2irTLe5KyB4UnnrI5N/flLATxZjqNCnuhXwQ2/TSykpKWdK1xP
HBY8czmelT2rgK3mZtTz5Z8Y8a1ZODUkBTCp4RxN05RQyWZBnbrt1IKbY7AGHo3v
Iq13prSPcQVZleSiqEnsQ8dkmshA6UAvtQ4ljVgpxFJhHcgLd8k3X+rOVa/pS2fj
ruAuXB16uj9b91Z8MwEjJmPJCw8JEKxxyWNizhYO8R6FRViCRcksmeyVFixO3Nkr
ferab2VaC4fcHYCCykiJ3Tkw5DzHLTtMwpRzVumFXKgJcrQYcgY6LzltkKlyMUh1
0q8O70H0QSRgFAEH4uLv7BFyfkfQEAjKtMXrKhhjY/Sj3fY5E0rAtt1ebUVH7u0Q
I40KPkLGXyBRVguTe+vmBJfRHYhXH9ZyAs5Y8vCkb213xwzx3z5OG1zy36HBjg87
mi8lg1H2yjlMwZqNppWW4K7+vdiXyBH5oFmL1FIEIRwg2f+pQMieC0D1OIIO4IRv
v1k7/aSAygKfEH6SLtX+PXB7bt2bHt2EVWk9UWfyLeA3dWbrggWi1O3oG6qXfi4x
Lu1TdQNPZSQtA8M629kxYp9AKvGJTuchUwM3QfRaQUEOH074vs6SZVENFPEaLZpN
/28ee6JqLkKePLzbVO6dh99FIPDr+wl/ZuKvB1FuevnX/P5K1T4uEIsmFfCTiAUB
rlH8G6sjsC+3kWSfjwle6qcrMaqJObLR/zNXyD7MIFnb5i+4F89bRbzEtxQLHDiC
Lh8X/abm38vn5Fjyw7fQGB/0Ysql2ox8dkwO/lE5relyJFxN8eegNTCbpbth/naH
nlzm0xWhVSeB2xkWQQUShUdR0LBRSpMNuNKGRB5ENunOU7+5BsRGpMilT18vq2YI
8vHsjnlsqIOp5JhWnUeeQ0ZEjxcNtp9KQk5gmFuZnC5y+srEjLtcBSUEv9L8Xrs/
AE3SwDedFjg1eEw8TJ3gYxvmE8sgzW1sV529ZyeBnVUcfNpYUd7rDzqeBOUd8Nqt
VWRlwQBA0qrnsFepAnqfm/naXsce3YanyWvK0VV560CtcB2snqsqsg71sW+VJ9DW
b4ni+xnwqRWl+uVbzAS/XcPtVDpGFzT4TABG4N5gxRzWqvS9wbROAnvOWs/yfb0/
ht8XiKjeFQ3dBuWI5B1vXJg9qY1ICI5yl/jeuLKSK1B18F37aaCaI24PmVsBD8f8
qMqW68L0kkweMqZ2eGjGaHf/tKKtodubMsyWQBCm+t3KGTWpp66ohiaiYOkG/7S7
d1DAcDeGA3EG3ZQ+cG9bIrXIGVT5NdBJOzGF4OaNFYxxc5FEV9aTZpg5Od6BBci6
8W+GyitBNArMNYFQEDqjKo1TMBtS7Y+WSCexYDhxC47SamJblfvgpPO6iemYrIAd
wcy4bEONpHYJdyIFmb3IVwy79Jj1qjvkbJ5bRoRTBrEC6Pf7t7TMULhUBxITOgU4
ge0JE/CaE9GZJl6HutDJN+MOMAEK+rRMOzNyYdpcSAwxgAqnkPFrDhrhFXNqDc8i
k7t5lafAO6GA/NzqOQq/AgP1FushfZ7JrKUbLFWT/RYDXJApVlParVdwi7dAtToM
oJiesEIdRclmP1zzAxPcNRVgFDA+KBFwnora26lQYd4H00QD6kZLEjmlZHW1LIhK
9S5uX9os9BWQ4kjfvKrivfq8VsO48tbjgrNpiW4jB1kdE/D51+aeBRDCrC2bbBhZ
YJSH2NPly6kRufaBiZFKqSH31I2DQTRSc2CSadsW47S1vSFUOvsnu58yEscQAByT
cViQGNep9TFl5jFMVy9Sl6IaCrDHxFFl8l+gujEQXM9D6nQz9X4uB229+t2wNPWz
2o7+mnGDkQCjTk2VJRkrycjuos+miSR4iKSZX3+FRxXL0A4vDWF8Xs7ZqIBTjrCR
wxfzFjH/ndaIzDHJ7AoHvMqRwzD2kjib7QUUEQmeOV1wBW7fiZxwyqU3BN9UvKTs
NMDLbEUqzrWJcVPWQdT4lM092U/y3E2mkqhjVpf3OKL3/Zt9gEt0D1ekiFFyRpIZ
kk2JHVjGg7BcGE1oUmr034lIqmPD6iui8Jctn/0gO7ADsBLC5nqX2mjyIHmJnaeU
YVOPex249J1OT4lAlzUW6SzkOmi8JS6iA+r2xq1g5Q55JRVYNzPJ2ODu9B+b+C/S
Ja+uiS/7NtA8mKA8T/RsqO9yAtPW7AZgL2sepYFXFPi4/iHMgoLDfy9XRuL/9jnR
f0A7kGoYoY3q0Wx49N9w0rk/iHozsUit2TatGJmJ1+pE7gEx80hnRcA4tt0wnY1n
tpRI/4//LwEXpQR0awtDoy6/AbaWDkxjyF1kp54fHo9A0BqYP54z4/HAS6oxUftl
r0wAQvwCf6a2XM3sLXO0XMySteJbgz1Sa7A7LBiwIc606p32TVvot1BQV7s+Ry7s
AYj0MXV+BxO4V2Gk5YW2zX85LnBfY5v/yZsTEIKVPbSy+6nGsHQ/Nae2tWrFTaap
i7ROTW7N9qBxukDjVarUpaAi9eySisKt+1Tb7H4gNGgFb4y9opP2LgENhDmbBs76
63G2V4riiAtVQVlGXLmEE1SRDbKRP/TIZmdT6DbhgXol6MDYNfQIMGIyjEbQ5JHt
e0BjAchZyEE/IuX0GywRPltsFL1b+dImhqzq7o8YqLn5zeTdjzSNUfdq+apVL00h
+AnKqMIgJTFq6bbScaXaSg4X68p1BMli8a4CogYXGZnvanZfCugDdv3SthCPEF62
aBEYXLuXi656hIhx7PoxOB27P6PixcyLwP/o6nGpk9zzH94jDXEBMWKiJpmg+8dD
h9z7jhCdoF2V6pzjLqghtnL1xiyuW/qLTLnXwE7XNz1VIyOYI/vEJr9MXWOvlIOr
WxZota+43xuMrI0mctCgpg1A+pDCiMdsIoHITJPmM5qsl1wxB8bnitjPWDjWmouW
Gysmk/jx4XK0S9/7MwHrMSPH3+iMkTHWksZiPEu0UFvxKtLSj+nsgNbbpjlogL9U
dg57t7uQN6x0ctaKs43EP/wvxOdY2XE0lfEiS3MkA51F1Yn+esrpV9ru+Ate6HMb
xQ2I0r0Oc7IYOAQAdpFr5uzvsyWs4J21f0BFHwYUs+IokfdR7FSOCthgvCiCCWLM
S36urDFNUkD3v8S89ueXzLEmB6gI4rWEIQtHgdqYVKdQvJPi0jB4RhL9cnrlPOhM
0sbFyMJQVyY/wiCOjL33oq15FxkELc6aFGlYhn/FlePmo+HgmmCtw05Fh1vuF1gt
u+6Vgwm8R1cwPf9nYCCS9BEZbE60PrFczPRDLJ6ImiUa7tUqE5Ek8mMT2kKDSOsD
49xLg6kZMH0z2CoAkDxYT9dobMksRVvH2TLntYsCsmbgNeU6To4KyfLnutZS/2BG
SjtmUi8zhL32haL3w1iTRv5WIqglLl/dMco5A4h5YZw/IBCyEH7/ofpuZHdTgrWa
ZEPX2ff9Ek6bxSma0HQ3/bvjfSRNS4QwupZHUjhMB59waJrjLcplb43iEebneHfD
8uLp7r7Yf9+4gP1IC8bjRvTcyrCHOnnHJkn5m+BidKH5btaLF0pVNi6XSYwoQ8+z
oxVgUCtzvQHx+RlsJ3rhtxVkaouRsxLM2AZA6O90YjQZd+0zCSa50NlqLoIWcpT/
2kNqP+NjLyUEY3FdmEz3hdsxWILXTXLJV2QC2C+CMl8pZBkKyxD2kWHqPHtn86pj
TA0sJgSeu0+doWeyZi1hII0gyds2MkE94OhZjH5gFv1O7ZeNTf4lMHdzLGwKhLJd
whctkZTGSkwlv4Qbknnq9HJ3/b0HONMQYPBfgUFbRYW98MiiM14a8sEjHnWW2vlD
egZ+yBfihUnIeFMf4B/gy0pguig6iR7JYzrwsoAXK4FM6aCeVJGqRqldpppmQABO
JeWwdjlFtj2F/09dQsJmulccT1oEAIFrs9Jhg5P+DRIW3PmYIu6ow8pSV8Kdkewe
TmOH2CS2sEEe0vPL2uCyzSjDYNR297tRR4o+tZ9Yx2Aibww3hJpgBAwUhAB/qtlP
05HnPe1ifh3SwsohBKhNZMAZkLr8YvWAR65OxXgh7SicyMN3i6makMLX6CynV0w1
VB7WrPrTQ55ady6AJvlGEcrTeGfQKxUIHfEALGbpxKsCllDRaHouC5Ypirnuh6Zo
+cbdi90jiCLM7xg4UDsbUS8Ct/hTLAv5zLYYQNJyU/9S5uzCHaXQMvha9UKdo1mW
33ry6vikDreOFk52VYL6cbjRk86e3q+J1aTzAvj2FNirV6mFVVpDXhFez2pHZGvG
IEHkZ2qRv3rhGSTTOMEElpkN8SBtqJTbS2aUCTbdHmviVop7Ao3eLeXaiYFV2IXu
DVxkc9sH9r2/eZycZz8Gqu/gubBnAyLNeqdjodoCcpL7T+X3oRWR4ePHTLZrFavo
oNLGN30QEUZ2dMU4uedf1oreJhtEUXa5vSYsZvTK2OKdEATFU8jd4tUdACXU3L/1
/8jk3PhjseCNp8+G1CCKke/Z/OwpmiYfFiFB2QdmjC3KhYVyjGyX+Jnjd7oOGCVY
pGLw9gZoj50IRwfC6DD/motQFz/u/e/gJi1bYF2AnjmptkLytFz8PtRxlfmTHCqH
s16igUoe3ib2CX07yVWyvtKDeA2wqi5MDvazX7BD3nXVKs9FXDyKYvIj3uFB0R8G
aeBw1Gh/fNV8V1NgHbhmWbMqJy5VLB3C91yfUDux3Di8WOssJ3F+8p/VPBYwRN7Q
2b2ioP4upsXtiUkDYk+2N/w4ezDfT8rGajZzarybzH8kqAQnTySvpjcGu3h/4zG5
HldtpdsAPaTBG01RI6OGT9UeAawli+s0Y6jZVeof6DjJkEZK18hPqiZjzs5ctpr3
eaExMF4JLE+H/lHHO6q2LcZ/bWBXZroYdsbMxf9wKJrCJn0RrLc+GTBTowO2eSP4
+mVD2mzlMDcpAENITpnjhkrHfqGlQ/y1O+9gbBdkGR2YuyFzww3iD7Vyw8FiTGf9
gIu8Of5BIyDusO+8ctugRmO5CaOBYeyVfUb3L5P7iCSrFHa7EInPouxyApZ7gWnS
fEFYguol+jUmqD5Sp8IXmq7O9/iJqEaZc4ErJUVx3dOEWVSHjj0X4LpIiiVZtqb1
nEr4syQBj+uB/wLxn557jBT+/KoKybZLt4IUlmcZRqt9zx1ccmx0RNV736gpnin9
nMj5bVoidZO3fe8MbXZfOd/PRLzuu2uGqLTtraAWsmFgKncfDyFOlEZ6nnqLzS/e
BagwFrtjz2K/eM75HUzjZH2EuJzF8nGJtEUFnCLE+v1XlQDiN/NumiFKulq8ppz9
oFrV9fzyz46LHwKw2ZdrNotBsJhBCKdm+8vaaKTUas7aPRR3cC2ST6+uyKN87veS
Hrt1XmVxgeiTu49J83w+Uy1WDPqwnMOrDPiLGtorONoq8oBaDNhakOu81M6kGs6A
LVdtbQZiikXINyEX/Z7y/OXH/ya3sbdQiep2+kh6Zh5qveg2GtHMb8v4y2Vyzb6c
LbhGe4YFOpXPVIea2nG2mP8mKKxyb90NUVNzPwKkfwCKc0AOkYcWSrL+MuH9dwyp
1biRzTT8TnqeQK/0GBxJAzifrBTuCAp78dp+VHAuxHC/P1PJVWWieC1kGl7BJbMg
2Hnc6f9eGHyUoVwv5EgysxqvglIW+tX2i3ueXVRu7SfP+M7yCaoawFWlapdZchK5
WURa3ccSCv/3ozOskfXkMx8Xy3k30TH3pxAke7ZQR2A/Z/g79w/2qHK7gkiKu7D9
Q/uYwB8JiU0MNENvton23IUegu1KJQLA4b8/jPdXNuBqrbXZ9YlMkxBgDWL3vsZP
RKKP2mF/rgEMvvkiz3zz6KoqnoBoqT8Qow+R2pVOYRhZ3Xasa7FRNZYcDdhuEYQ2
Re8mvY4Kne9lsD88n+SkxjNX6oM9oCIgVFTDMk8wRsGigD2diF+w8jIKypvuGfnQ
F7n8P5T7gOwTl5Q69gNUrx/PBmaey+nZuPrDLBB9W5XgJUsljh67Kkj+9YbDfT61
vOt9aOpJlQFNtj1WGWzZnOV5/rG+kw+ADoe3sPaMR9r2LjF0LS7uhuQF9kyWje8N
jl+XoaTI5TCklo6sM9EsaLnefLTJohvvYvNXMaNS0MRBhzhGmZq6K+V06OeF3IZx
ViVi/pPRgS+rlV7VAbwXF/evhWAQAQZ5NuSCsUVM8seJt6354Xk+ib+PemwNxKV/
vF+lCmdMYmD6NOGG8RX4DKSSu+0ZBnkV4H7rIFL0nesF/cOqcj9bm4qEl2hJw7Mv
PplkwyxydfuFc/MMpfYqP/YquuQb3E2VLFxumBxuAlg0yg57iFoWY7DfBhBLut5W
ertql3yG0IV/ylFfa/s4G//vQA6RJAaf8mdzpMXltHhZzYFcBmWByh+uZC0oiXFC
+aGP3LQyEjE9xAeutyXt1ovyLaNYwqYjEJTwebjHgvm70Kiplwx+9bYVk29j8lvU
U9fpaoYMOc0lAmQxnUp8gpxxw9MfrolTk+hId/HaddH60waO2HXkfNlgB3azGmuU
8XxtNqmmWP8BbphCz5XITAG9ujtOu+eMYtn6IWYEUOnTX2z9s6z8vI0c3taAdlYK
6gglfhoHoWtJSyAeYIIHhP27GhGLd9NmkTOKm4n2UksCxHHVHNhr+Iy29q4hoHqO
D5CfSSVHkCsAh3EjWMZn/gVjBVKP9v8FBX+KLN8EFN374ikJf0qd50VyqKjcXlAX
5SOc6JMWaZ3QfWrL4e1mc1geR9JL4I4+fnyfBVwPNbR2Nw3CvW7z7NctZZU3lmg/
tLwUEbBLo7r/iCZrrjiQeSBoSt51RM9z3LG4xKBQ7pw+Qsa1DRoV6Zod6BbWjfsF
RNJHiFYerS2DbVQqnDZCG9t+jzzsLC5mI3UHfGNuLgcxnLpepK7MzEZmrE18bI4w
/iZq3ZuNtO6OwERCr5uRVAvg5lDrQLlFRhiZnqyp9nnNeFJxX5OK075SJDaXEtFt
Pz5NNNimL6tZP/MuvLePaHMQdK8zqIZPpsFnNTXEENXF8m7ogCq4gr9Df3ZsotOi
fB1yQ9uF4GQIlHBcHJ88lLTs9zYopQjsPf0wivdmvzai+T71z9n+ggQCALtb60tV
zhksfM4+5aEYBeucGwAWeJ8DvHL5KBss9jjmpTgecO+9BFO7dOFbKKL4vlbQ/snA
Dyrr9b7ph9ht6vt4oiDSdT1r0YcauRKo0xa7cfZYvUceArr4GklTHWWfjgvXSPFI
N/bUEkYyahnmpW/IELk7CtvN6jUXqcaf2sC2Quvzt9kTQMTJKJFjrwWCGXMjARAs
mXQfTgQ1zx9hMvud8Rvx2TM/P6fCDmwCvw3T8ab/f2OuUAvov26A6S+tzuIjr8A6
M9Fcx90xLZwZQAThBKGyCLRQENrc+qQPFK9XVReJ/hDxWpAW+csemm6wRblvU0UH
AIreOiipjCFKn31rnRbAThgRECFwM+NuYGRUyNPeHTdf7gSO6ph9WrpXHC46nrb6
5cUYzQSXdkPmMqm5yJSUWWITx8tlrV83JZNgLf6SxhX2ueyaWlxKykjsDD5tuNy9
KfCEfEQqawzFiQDUXXWNVyJ58rfjq2KYkLuEyFvC4E8YjVXJx92+77Sdw+IcSXdx
7Gnm1ZlQZxTKJVSGqKcZXT4cg/G67bjSURAiyqbQiWzwaBHAiR3T5030QXO6l4WK
6wp0HE7ui1Pbw3fZuGDyEV0x6kWhDHIoKGgRr4n4ybmy9scpEdai4ChBM6bO7Gwq
PwvVEjaaogBqLvlZwISxC0WURUwUrg5cBfQXFETmCQSpkiroiWsdSS0VaduPClsP
Qt0ewwAWluVjuU1LjIAYPbyxIHbLgwoM6zP4EDnelc0Iw8l5ZwsdFjIE0EUPdKVX
L2Dcc/HnTdBKruWp4IACdzlC5u56TyIVyBsXy050RfxOOSJ15eW9Q9tiI92RD3oB
0eclP2EXDgFBZgJy/v20cQP2JdI0/7jjSyXAJu1iBVhSyBW4OcWSDwBf8NkH+d5k
Vziit6f34VyNmBMXizy+BlAd5dSiJoqEToFeKox3sP3rp45lsZC1jPSQP/HdTACf
3LP+VZAhibjtFGQwZML523B1RUAyIUISYWLdd+CzFXZCmKQzEPItPY64IlsakEmS
nJuB4AAHiY6cl9jM65RWUP1UjkKnw608CiMddyri+PPmYWcp5+SlvYkbh3PXMupP
8kGD/nHgOLAc8SuaVPtpItBj8zlIzv9LArcu6N3GTARdUQSnAr5QCO1Uo+hCFzSu
0aCPCPwVxVHWZN5e8RhnIWrm/OOAiQjc2fAyHLPMyatQ7+or+wCEVRWcxsW4HcM4
gPafsE7GcaI5yzAmjM31oXrfU2ULNItEXRhu9tK1x+1qWXoZYRrZAc04t2fcRjQ4
0Lq2VDdpNLHHQ+6xcrQsQyOgSmWdxCyF62EJ7VWvGyx1x3svO7szNeE6ZNJeR+xM
d5Z1Wx78BuFNZlbdmsRjacVlryfR08c98J8NKV2uiknLJ59C17q43+MNsIfh4Zm+
AhhY3xHj+s/m1vkmH/ExNtrnk1L/FdTFqXcsFCAUXacy37tg7ov0S5E5qoRllec5
jATH9Z5BQeM8MFJ20vxEWbJEvZ5L2f2sNP0rlTBexRgBI5XzZxg/GBKzPvQ4q+bF
oAcGGwz0wJfpMNMhMmJ6A7y4pfiq3Qu0PLXjP0tgZ4I57EUv/Stu0u/IeLF6z0HQ
v/BWV1evj7CDlYEkpdxMW6CPNpwDGGlFo1LTg9VGlJoEJcvLkp58Nb5b2ag0nk73
Vnb/1lUfhoQtWMX+QBWBzb0cbZbiixZK9M2RqENMzOtujgmjQGcYpk/tdwtTpq+c
0SQ+ZhcKlwC/4ICsuFC+oaW3Ll6zCOSGq031GR95N/hELkV6ml/YQSuhQemwi1T1
xrLEo04RSTFm/vNyJl0D6gQNlzNqktCPHokpaOqtq/GT5qBc4xzU8k+dFAv9Zfdd
Y71AHt2smrMywy1/+2hfXmz2X4e/32i9qgpatRz1uLLTo4hfqQBUfquw0G1Nom9O
c00eG7Bs1cRe7DbX+GpIEfQnyeUDP2Lh8WMxKMVoqIiqujlPriEDYuL5eacCjDbE
ZDJXok5D0R8JqEZUqKKuse5kI8NuFeJcVhyrXuQ4OC89bATifTwKlsFwhDLcC2wH
cE9J69OBvPJvTJXtvPWqGj26j8kE0BmkTMVgze+kiHy7/Vi+bcJdA+d9455UTpMf
1yTpGX0IbO/2zgZacq0kZK0gysfQ3C1W4gjtASSB4hqluRs9jumVs6ils/iWvr8S
QmoMy5WRri1/cQ9uqJd2uci7hXUSwGBE6ehpJ44G5bEC6ninLmDuE2RptrRpBIak
16HTnsvl9G2mhNuM207yErbrWM5NHc593uZ0nqJblterX4Wotx6j+cFoA9W6+KOp
WQg2rId2ftErSWtIa/L+/ff8SgT7RM9VGwyn9kTdFdNqk+r0lNhgr7bEtMB1Oaqt
qDBdEkqPxy6RUahsJNrOS/6+9aX/ugA1YrEXW/1Vxg72JwfelWKOnVqNVWdDa60+
gRZgabaRDulzcerBAtkA3R6tHS58LvYObCFsVdOJO578GaM29AY2GMPE9diuSQKq
3mIBIGrQrst9n4jxc5Ip4XTWwBzU0VLHJxR50ElaXFwNASPa3fOoN2/cU+CWBlVp
eDwLSF6/reQbzEdyp8WDqlEjfwLKOVJNyyxTpV444mUujHU5v2uaqltJj65FO3CG
K7cClPfZCHzJP1FAxO3WHhDWhDPviaArcASAeP3s5HTUY2yNDe91NAY1zenxssjx
MYxIHWPEdef4VwAgEPEwyyKNtqQHs8hwQBMX5UIBrcEURUPwBoMGOwB+R18KsYLO
fe9N+VjEV2ft0QeFRgEDIEs2oij8nnDidRzfew4WZDRkfondDhQS+90GeyrtFI1o
SoIeBNzIgGjRWFB2r8Hi+zeEjmtVRaeawQ+cSwoqlJ2U5lCb4If135zjbRIhg2Ld
RG68Bp8yVJxPi5sarwPl0SN+FwrYx4P4tTkHQpi3+hfbqrrpNVIy56anKARGa2Gl
7y4B5yKcOapZYWURN7Nmm0vj/B61ectmFiwPBmALIEb/j9TxKjWAIGGHkLIYZ15w
oakQRiAw07cgEnxpmCBZBeCjGq6NqXsGgMC6A/N/IloL6aEs8VwG3tREN6JF4QV7
IIY7VpwSoxCr7UTMQq3qCOHo6YnVpumfu7Vm2PaEOJLwqL1AI3WQE+f2feKbvx7k
UPM/SuWIlo5hGZwROD77kpJlWkzeKcBbHNdV7B3CvuAKe2YNgQ2j5ACECQOXjiN+
EbZvJLpdyW9K1CmFR+GxpW+ngUqbqPTftcXBlBMpgIccCRluLOMh4eGsKjqZsa+c
AkvVSP4uibvf6SwlKr6L9dEZTXDQmVTemQIKTvZheV1rBCaRlILHBd1EIbaLyfrP
5ulJQjmoImk3cZYtxl/IuL+GZ5gUSux600lHOd9m11hderNvdpqPrlFj2fMX6Swy
OaLQ3iIZqhpsJK9+VQirVJPQD1nHJ8AfcjnEgy5Yc1NpClT8oiNZ6fGh/2s6Tv0z
WQj92OgCAhsQSEuBua+u+bc/jJTYSPPhh6rTMCGT+1aKYo56kOxdvV5VZ3uAVXA7
hM3fansjuGD7q2dsrSykfRt2qo4nEJ8qg+cJMgV+VOFfXFnjAHdxJHOmXWns7td1
A87fwAwmATsYIDjIYQVz9wCEuFnKs9BqDD16JmkIvjic0JMdb/T6nTh6WewPLNeQ
q/HFWaiZEI7W2VDHlrjGvi9mFoYbdpOTOxqdtL3Z2kXojTWhLL6UCf0WOnFaVOV8
PkYuWZR2R8IwwY+I7l+eNKgdzZjD1d1wR795ysNOorQivs8H2Ef1VJbxjCE/QXys
MznZ36v9Mmg+39KU+tq0Ip7drp0f0KWHSHWVq+EGJMPTIE92oLvwwSkYt4fBZvTA
K35eXZLC3eZvvPRVlp3UwpiFsHBMPAC/h8Lcfr0drbpMVe8W7a7f1v7rAdPb6sYx
6ggJocK39p86zJa0ASeZV0oS+H8BXXD76jv3xkW44WLZfJDkGnJqHZlJG1BkCxGe
M0RW4xvOOU+9cDaRCnxvN5Jh+OyKiycgeQt1yQiZpKNvTs1xc6sXZVMvoXt23xEJ
uc4Ixx52O//ms8rTxLfcqy7eEjjhApULdiy+5eTMTWdR/maecl0YY/Nv6NfCW0vG
0+xV+5SanES10H5I7ocVluIxp8stDEXvLlq1+2AF5Dotcwb7vXjB7F1g4m45ArYz
nANdyiC0EFPWCulJ/KFCCkPu5WOCYTOtjh1vxHPNuqL8rqw5yJJVDeIkhzBxPmS4
KtUmy9KXaTGvyRVdSC33GyHdWZTL/97IoRuQC/E7rY9XkkPVw2LXw9S1+0LJfWbh
HctX2cjcaLojzdRuPPTtAfUZdQvhsYE+hSZorjCG073+wbye/y9EfN3blczDa/aG
w74jNU5liexdWWhqmHaDd4Ot7O9fsfKgW8J5nc1ez0F2slzwcN9GAxm/jVpgNS5r
bE7ZiW1pBsXZ+s7uFZ8VR1M4SF9JeRc0Lyzk2c+zwz3xjKuaSGm/ZHJRjOruE+AZ
cyvU6vZZZF6knXXRqBofQkBJSi3CEuK+qIt9irCvl8EsjGYyrwXcKfmvYEtZJBW0
H1iurmAHwPLNAFO4w0+IVdgeg0PuBjCE20Nw1IKwM0ljgfuRphY8P17mu3QjID2w
yLCQ61DOLQa+Q/5zvGza6iBpo5WTi8LOnLZuFQRNYlZjTJskSamy7J5kCsi0dJsw
z9AcOj34/QWjYT8SJ3tDhvdL++FYaoRHU2i0A+TSMTmzlBQZ0KGvoK/CQsHakwIG
tPm1Rmnq9LZnAVAVW5JjX5liACeH2RsIk0S7AfdeFylWNXyDkxtYxiISj6iXeoKO
hJGPbeSlEQjzpoCG5CDhy71qSl4pza1sCwaV3wqcA4w8yuOtmS9093CqXzoZIkyR
j0R2mWbKO5k6LEvJCfJFqY1xsh1XAhp110mdO+newlWjibi1G7sonf5BqDftLi4D
yJm48vyl1nL1Wp/SEue1J72aD54WZ1WmbqRIs9aE/cdxmodkKQJBXMM3O4X0V2lr
lUpRL+Nwmwrp0i2LstxxuzuFiI5F0gAXR3zj4nkWVtO6HTS41zQ7kNtahhQK8UbG
jDGRXxNvFQ0UEcCaN/Liq94QeOyRBi56pRVZuCZ90IPTAjPtebDpv6KbUFRMNDFu
WKSfAWf8izLwB2CVHYhIM6FKrWL3DbCxZIMUCL2Nx0IzIigIlzWQO8cl2/LvdiE2
4sTFxYnOqSR0WiM0Rb0WfkUx93uQ+px/f55MfBu0G1tyr5YxJSXXh+5eH6rIccwB
ufBTfluWVnKnxkNfVvUeY7pfiTr4BoAGrepVM8JaxbjejgFseeajng202rmchGXP
iv5+0niWL9jttrkEDPfbM5rwM+BXSgRUSVIjLru9gh+5ek7/6I7Jln0IS7kKt0+w
Yyd4F3rAG3A/JjXGbeQGDPIoy1PG0gz1FQDcex7RvWsTY5JfYjZP6AiQulK1sUYv
ZGtYDHmQGTPwbCyR4+U8GOVPflSQH1UXuMh8oXS+pjnkVB2ScPjl1CuZkRLJpuzy
eRulvC2qNFW7y6wEL491rx3Dy3LIP4q5lFjQ4AWiuVEl1kovXI+d98Bd0wHgN+bZ
AXX0BuVtHFkwsRvRYWQ2+OjPkLimi9H/0Q+uj0s6atZNJimDWdUHLimIS5MM6lta
pyIthC7+k7IBTjSWv5TR5tL4X3QoAg9i8d5SZ7CCJKlrsb4o9Hn+blMhOX0VpBkZ
nSMyJGauy7YmbgjU5fbRDIcCmHO6rHDRGDXFS6CZniS6e6FEFN2EZ27SxIB+xCtc
J0PP7hQyRTClZivJ4dUQ9pzdCx/Miks9HP0OmnDHNVZj94oITgzSxfZrsVi3u2Nq
0FbeLfBcSzeRMZqYkOh+mnRA2BZbyTVjF/aQtn93n9Blkd96AxI98v1lab4xxV+1
+YqZMS3vZc1ZzaLYEoR78g2SGqdOLmTqdPtroTRazIbe28eDVhvMHY7X4rtuOdNy
zIpeTrpoAuuv1MSGpdvD61OdGZkt0ODAU+AXG/2dDpKGpuJMbYxganEz9YGHZhyp
fLOOwXlZC6Xq/C8uIc9uVFGI4RqHv8H4Sl38/EcVqW3P/zTBOUoW3G2G2H9+/8BA
mvlwMLbRSpGvQCf/xqul+Gyby3/L91sMtmqWStWBNnBt3u6GDCdQzTmQ+e4PqaM4
lkED8mmfY8ZEIqrxdGAzcRt4u96KdK1FuaqkOxQLvRRObl01VAfMvd+8eKAiekgT
zfw/t0Gs6jse8DJeSqNexFjaDbBzJm7wzSWmrtyJUFYj5dwBBKmKcdNuyyjaLRH/
UlbiSPlaS55hzneTo8X7FRypzKSzgodHnUVTO8POsWUdJGezfDZIXjXSXfuMnce8
BJPcvgnYjdMB2fWb+wT45/IAA8xUbG0aqVB0ZqW3E3P0UIfOUDMBErIOVehc0hzm
k5PqwlHKirwUkAc60BtQsLXNoq3FkhNnQQlVrnleXtIA8MV3EiOSFfGfx2fWEPZX
zFVO9tnGh78ZcnmCFf++pL5Bw0qZdSWjIlHz7gFE/twWJe22WYZ4J3Dap4bG5Wbe
z7M/Zc3OKu5HbC8x0sVDlJjnln48XZVZU1Z6LsGR9tHNj+CxBaCZJl5j6UywSvdy
bgIUdWodKZVW/PEkAkwY14fYdjOgQhoH5iH0IZ8Kd5a3ZOV6x7vHei8QeA1XndVX
ciawBhy9RfKq7pFkDkPrH51OY9+qp4uaUbH06q/xQsXSoA8PYh4TdQOlpYpxfsz8
68uJRgy3ZJa1snOYmFjk9fB0/G8GpmJaTVqbkYcoKSWQlvccXrwuTyDHvC2ePl/O
oG1mInqd50HzJ7gUcLLgc+aZNx5l1r3pYD8ZELpup+63mARwuRnFRKozEHJ+lGUA
i8aJZYQcN+9QJuh/fZ0i0jmYkQdR47jstPGlXzQnlF4rxR8k9Z1XwTLlbtFmFnHy
q7NXXecUExwD1RD0xALaOL2GwfaCvEcwFkPjfrenF0E0Q71tAqEWzGXDFUWQM7mS
XKX60OuW5Aqrast0WtKdUL8O3Ig7fjkT57mqXiSyCtTrAN93MPQeijhNVqU6UgI7
Ct6oeHdpr+pqLbYa/dtZYU8RizFpvgd3Rz4yhnjUSbsgAroVfL2z0I1vs/5bA1+Z
yM9tC2KIyEW0aFzPZazIAuLp8MDMO5j1Gh0XerRLrBcrlpuVStMmgIhLuxFfunsK
Mh05WwRf/j5qcy/aguSh1dEqFkrYwmU7IzZOGVLFJ4VNqxlOrueCpP1v3VPq3Q3e
KQ+7M3LiWhX2Zoydl6d7sReaTfY2a7VuSG6vSsIutqbr6bg5bvZ/Yi5GnDZb0l0m
Lt6m+XZPJkKyKWoyKMEaKow+nLcDZ7zcWY/ZVioNKS18ypnvwvJsmEKx+U3LXPiL
/9VAxI4z+SFgApTmEAa8uoROcfM77rAv4w/TutTedgjKfLEpdaHUL4bqSREyZdHN
HMF9eNpSqOwIP/VNLjuLYZZfe8gugq+NNB70Oe34WDv8woOC/s3PyORyqIyMqEPG
2kqj7Kk9ebkUSCCM2ExGlHTYm5Wr4+k77eZ0H4Y9/FURd4eRNqCzuOAwSk0qnis5
zIG/xs4/GLPeoxiTgcLBIF1t6rkS8jCGKE+/hesaOMJdSNbA8tcCyJ9wPqkM4dZ7
xXku6BbmbTYL+hlNsvei/56EddSFQMm+4ZgyWXl0RJYNjHInpAwqrHuxgxfP/1cw
QOqAgtNTYErdSUpAeF512VN5XSOk7w85knkJfcS+djoOEX9m4KugOeblkhWdH02p
Mr0xu2C9NKR9/AzfoFXWBqH+A1JiiCJp9xGQzsa2U9A8OD5G4TU+HwYMEys/q3PW
bgI7dY2BxRoPfQoIzbT/6E1TzroixeMuWG7GHMxMUOxBuk9nxs1UG0JFHPIO9K2z
LAh4nyG6Q6/VJ1U1SoLw5O9puazuQeqGAWIgBwmoLBmHK6fBKg5CowgFwT3RlL/g
FB+aBTAdftaZLVF+vg0OuuquUnV97Ts4phiX2DgLXIot6RR/2kzEPZUTZWdf3JcP
24gTsmlr28XAPcSiNlkKqqUJcexz9xEmuXHBchMuUO2KowUp6FZyX9te4UbqYn9G
fbpp3pAWxJNT8Jl9u4umFAxKRbx3Q8ooJyCoWvFwmJIXZmQ0QppDiVzRyNqjpA8E
OJp/I4ykPxXCQO7paor7Nu88zmlZ0bdUWB2PEuMFAkxyGptlEyWCU+WvB2UKGdc1
Zqw3OW33BlX0CgOkLrM2k6TEhdM8tkWfI/g3esYs2XffU17tWnPGxFoPUr6m6/NQ
3gM9DFqjpYxzScxjGI0tAcecBc0foEraXheYFYkvevRbKx+p6VFtVKjOqpkoaI/Q
rj+9xtOvpsdXaO7VkHDnEVmEUZ8GombPPprxoH4Wt5VJMFiSGz7QlU8xHR8Lb2TY
aJLsPUPt9KBzY6i29CR6oYVQHN38QMvdoEdYpXg3sQlN413bXhYleAU2fO+y4nuh
FJ7uo2f75ooPzhLonAT6leTMsJeXXgQv4B/3o19lGWgJLiD4qGwuPyrRc3zhomF2
YZ/JJoe9fQxPInVdI0zSf6jdDxy1Hnt5a3I3yNgaafCIB+gUUJ2nrdIecPmB0OGn
BtCCIT1oVxyXfoNzLLVY4Qx5mk3UmWD8VDI16z6Ntyaocx6sbUbqv3KjTeRT3RKh
1Fnebl43nuSDB6fq2XD1y9CKuh3H4qacHMyzmzmj+d11pw5k3VDF4ogZUF3ArY1L
pY5FpxCUbe0Pg/tgXIrW446cyCmVoqDjntvyhT47+F/YlDRkusAoXblSLF54FNyb
0/c/venrcsv8eaMqQq5Rcr7c5SQVpJXEhaFbujyDLFPYR77eeiDvD94XGiFeblk5
VxhpWRdD8ALzW6PqvUjnQxUnZjZPN7DUZBOrIT8Eg5xSrpvZFwww8PrfUNBt+fCt
kwM2ncD0r2mCKD0MBi5i45ZZaKkwQRKkm9I1DmSxQv0Vs4xA5uwwsvlh7YBIsKgx
+6b351CKDxjxLg0vMp7793xQePJy+7dNi6OjiCNL5s0pr3off0YMneOMc9PbHGqh
SpkG6Kv2nvNHMRth3ZwbFSrPrVAZQeBAw6hVwq5O2QFSrpbu3iVrs8mtrWmRyCIC
b8w8Urqe6zJRN9iZAzv6aHUcgWt3RML+xQwS1WeIYrQwixEN8jPBdnt46MpTbKrG
P/QYGaKWPZQnodhvyq0qKB0VVtQbks1RMQeMBtQPNKLZl9SnVvZTjXnuIlYbOeXo
erC7CE3+JxVKLP42ey+7g4rGnlM4pTbGZraV91Z0qMY/0PibwgCzESgkcvbLalSj
zX81rlOkbHVjrIzrGAQVwHnYkNxgJHcK2lUPR7UqAYuOHpZgSeCyrNFPmydvcaqG
rIsSTW/Fdactel6q+tgBZsBEPl5aEhnpSwjbHWKThsmGQvlVEDKdtnFMrj10bXYm
6rEhCpQ/B8SFFq+RT+4jM7pyfU9k2VqL1glsNSo2s62Nnlo9CLa6AT89oMfDWIt4
K8rPUPGIFtVcR+2tr4B5g+s3UCRwQfC9relkK1NP43w3QhvYoskfkEOe+EJX4NRb
TpKPKPJYfbq0XPrEMZI+Sc+zlVVapMVKzBXdI2st6nu4w64m4iiaAw4opCOfLB95
RuZqKizwmGfXZCnCsbV6DQcbojQpELwsM5B4ohFSlfS9u5D02BOrgByKbNU28JHW
L/NBFIa39WVUdxaY3y3Rnsy+zAMZgvtKBG0kfZt+HkVYabboIHDGDeP7Im1cZLhx
JeKNV8H6BJz7xYW/vQhpYMugw5AdQph0Cnl91V7RPv2Ob5TkC2W3uj/NwSfCnuwX
477WrvC9V0pqR7+eI+7N7GyhBVbVGDokm9Z3B0OCEPNUKBnPZVvxVo1jBSWr3UAf
cpFuahw1eWoXJc8tWGV6WyJ3tuwE5ZQfGFV2s061NDpGYfUmT65bbU1z6Spl+9YY
sOXSZOVlFtoaIt3B8zd/mpPE3mJX9qx4d8UlgZpOadiwJ3Rg13je6G2Wo1aWdaCR
AuE/V/L0lPWI/oXgiBVg0j6olM4T4erFO8dHWDiZm992ulJaDoFxpRYPCTCTu6kf
2noRm2w68C9QW2DEt3BZ9KMo+AtpZp+Q+Yhcm65J+fB66v+0cBE/AlGZSW+ROQjH
o5a9oqW1Uyd/tj7WbcFe8myxNBvu1hw2gvRDITukMzWjRd+1J4GlHWKsDUuqs5Sa
/rbC1TbJMARFR92syqnzQatLM71T5+X7Yy6T3bRNTIFKJ6c0HmNeExrvSEonUOoK
CpGL6KSZDB5djrqTjWWsbWnPDct2NkBVsNqBQNrJsb3eHx3Dmuc/O0JLEqC8J1w6
XT0hjYsl301c9AsuCetn/tOy8jd/lWyN7/B1QSEd9HDMoVZTB+lKhZS0kyTIp99V
5KNO7179BTWQRbEhH+e2QsmWpS/cc4I+RyrOn4V07GqODGPZVU9GK/qXPXz95sb7
8o8iRgS0tevukg8Ja3i+0FVtCdZFNQp+pqu4Msp7YMGbhTkV4tqiYV3j6VHzwS61
UK0ugSZhFJ78KcKTVTK9PP9peRizM81tDToXuOINyGDRE1EP5NdnGe9PggWcTSKe
wU+n1sJBKyDFshmBcPOAKROYdYufjVBbtzM9INBun9inE9VfgjaUZ0FOfSHvdKOk
e1BpsFoPwWj+Gpbu4WhoSf1D5bh1ny2ciOuoEMQKKkxGgrm5U6gSrLiXYgBPED9+
7QevWNmsnkLGoyyyQhHYQ5zKnzO70nR6g1kBRkcv/z0PzGVFscW1Wd6ToR+/NCMo
FnY/rMUTrSIgTQn6o5gipceZF11B97/A/T0kvRFD+ZVp6PNX6daCQn7rA6GbJv2T
0gQfEt89K8G6WRw4rDx8/Vj/9rXw5B2fd1FrFcvqVk9u8e4ATo2l6gR6LscDcywu
bhoWodLQQkKZl4QpiMKTt/lpmvV8miHSK35RrUE+0VqYMZtwunhbBOLmWkCcFS/B
qW7x/j9gKqQak5ve0zeJtW2hSyngpa7WUGdLALkkQwOLbh2HinxGAKBiF1i85Nea
Xt68YANANtk6kbpCzlMu33qkKOBE4P87lfgxLqf9suEnTxWqsxZmGsQ+n6x1sN4x
wV8FQwCh8La05qinB4XwkdrFC90yBTJ+u2OKyM35mEnQfQli+LxUOCCt4ExKUAY0
YT4cQob9+NSAjjodzkj3+FXytCnbSVPJh1oHaUsqDt44OfRDovSXlU/G/y4RDjrs
nH1IiWzuL4RgPMKFRG61zcixl4wKPd4N7T7uOiecZO9ipV+HEMXgNLfuBDCjPYna
X2yHcvJVcVlv87pfzGa39itrGFrOcFhRLq7SYPO0GFvGiQKPkNYVVwX878mpOYPk
zcoJNjXxTMh0Aduozgef7VXFfw14q+XtZUKy42wJpafet4AaHIG2dY/GAstLf0uE
md0isWzU94IEYyE5/saLbiA7VI8+5WVXhEAsjbqm+CvWrulYvAwlvJL3sikieov9
sW5iQwu3GInbV4+dreVlU69DrSeFD1u5VzvXt5bL+DCHVNYwQa97Smh9YyD5uvX7
S8anhh0huoFn9pTbSsE8Uz8Yd60uIuYW/efMkdHoXjW4ILZK6r7EzHsxJqj424p8
RtL6gPGi8VTS5kxq7E64Tig7A3YAPyB+VhOrdQ1b2PDkZVQBH808zqjrE9gEs8jG
ZU5A2VGa2Zz/mjptr8BZJZJ5/v8ynlORaSHPnXjFRpMlSUO/BNJ3zzbZxK7HYETg
8Gmguk2d8qCdQopfgrNfi4JEr1QoMio8bidiYHNY92Mxzalb3R4jR2nfv/acr3S9
Fsu3vumGRaYOaeUwG7LBfdyBWR615AS7Hd5sDNc4dUoDu4wtglaB7MPUgiqothLJ
9BHpLU/bdqtr3wMhx/rJMcXr1BwWHi2J0QEgkKPBkDyrL9RxrunNgzmgCGNTtHB7
jpOg90MVR1jcU5H4h1UJFt8kjuccIqLlqKOR3FvDsONarhgsMFS8E9Abg6JCQEBy
OElkUZh6TvEE/M+PqBqPoIiKj1yUlUuEkp2ClLsKtM8giO6/RCWyVHfSf4jnodv0
m5H1gci1VJmDYu2iyvEyfbb62LrxDHbvsPXq4MauLO5L4VMCru6dhyjoEGyZdcnz
6/jue6v2rebKlmUrtb7p0695Gg3m9kJhrVmvUOqPR1H6DnIndgF/2Uu7aPI5jJQk
oabWj1repqbGsgXx9FwosJDd1V95esA6s/Ubc126wApGBIu1GvdIfJgp14c5QuA2
XIdgG2+k/aE2x4IHrnO/K4RuwI2917c1KxofWfgNL7AnIOAipm3fL7obYMpNdTxK
9IyLZX60RgjKbCPnel3I2yLtCdKxqVaNbuJFemZOMPAPNfd8Z7HWSyklr9UXr5tR
Fcy+LxqdHcjM3ZCMG+HRldC3lHnIRZ0AWmXf5rMeARDE8UJc0C++YHgMQ5gIsFhr
HDL/HsWXvpVuczB1iuPHX+HtiusNNip90SEVYhHop7RpfS0SLR7VCFy9o1iWZTOP
+By4R6PAiECeSsDNjuRF8iVXxziGL9TTNP2d8XxDJ4YK1QDxaK8r28GqkixbLHhH
Zn0cK6caNmdeSL50MZSNU4MTFdpXVuhvxXq2YS4ewVnhlkX3ovM8PCTXNknv4DOW
uCu22XcwHG+7igxUhqBBHCpTaARVY155uv10SzgNxjsYDEu473QDUGyxuP+bOLbM
SRntUHNCoW5O5ffWLI9KjZfHoitLwJLIwn87kMoEYQwWEE4evkOk3DW0KQJQo86L
FU74yU+vLEauiJEOmefhIq5EeD0diUxR8tFnWjVToNF78TvDyYjizG4s6h/Z0IS2
7ezrtfT9+zB5rAl8QLMFmITnePP9HTifREpBNBU0HIfev5iySdeiErhQy+Ihzy0q
BYzZpLyx8nB8XQANz4Li+88XufgxPJug+goEWDunqNcSqqVdFsccDNSsKqa9rKGe
HtF0fEXcIwRzVc2rHbk++pqRpsghcCHTPu3/TUFlo0/AwHoToqmV+hQlONnRvizA
oLZJdq6bH9hAKbBBH3Ow6PjdJEY6oWhVw5N8x7XuLIVRJknUp7REP9qIB+xBT4df
6a1/ZYQtAejrga4qotoyytJuMiCK00QLkO4xuatekBxNPGGP5NBJAIS0KpEW6uM0
myhtANDQ/DRirSFc46Tt2vx0an9yik/vpKS5VUbJ8HdBIdAs+SxslLIgoltHQVzj
7RLqmfrtxYffIfUMMGQTILTxisRzjisU8qksvfa2wy18VxGoGa0Bt0AH/Ol0HJT5
Ybk6ybGfBPaB1IN5Mrg1oI061tUozuUE/BWtnkCddLHJ2f0SM+0dFZ2HuSTlCjPb
8I1X8qU+uhk4Qd5WbNnIbNTAqcMqkdEc5MFUw0mXpOq49O2R6pSrLqOwIhCkYieh
wsd+OdqGV4carDSYFkvBgzEmZDLMMnvS1iPCgu5Zmdg32SFVMe7mjfQAsT0UFrWQ
GFiBtoluXxjSmxNQqhmcwOyN4P0gWxKhOVxtG9Jhtc9PRK6xVKfjqeCWq/nSqxPn
VZFouwsUohuYd2z58lR9V5k8Aqkyccy1EU/fxpRjbQPGhMn7vNqoStX6piXjlj4a
kTOK5VN2HID2uuf1p1akNzdBf+LFoqTyD0PyJua0pH8lA72TTYcg4IV7g7pzn/Eo
mdDRvzr5/v9uNSwkFCjzwJywUDaocddWtxAR53yp5f5LMMdEIeG/Wh7YChgqLFTI
LeDthtxt8ctAWagBLZMZ8aAauvvW04Gm50zhFBauJ/MWptugZTFtAdO5cdI0ZypX
TlzGnKXI76mHWRImvdwi0UZlpT32UKTQ/XPfioG/XRNaTRga+gff1mV6TDVD1pq4
qaBAoYulSM+XyF0PxPdJgJ+cTVL29O+0pgjAe1B83MNyfNSHLJIe9sPTawytoaTe
iXqunsiL4RF6crnRBQDYTr+kHA+UfvfRGscwI/oU0YOCQKKELahK2FIj/0vjpvyW
svQxJvLOK348Nsu6wzZhb8X01RJB6rQyQRCNEm/T9BzdyLjaFSrgr6CSADFz+sql
d0v/yTqM2vE05FpIbRil6pRFiwJBTd8fIfyOdvT3WveSiMUNzQdvmon5bZ9KqNYk
B7J1DBW7ebgcoh9tRiiArL3seNi5W9icK5qwXU5Kw2roLKbBur0cSV5GOlPoXapv
k4ca2mL4FsUwtIxOPYQwjRvIF4lgKUqjh/jqwLSz4jraSHgNONojxQldl8V8KGIC
ry9Xff9phyVE+RHhoOUV1BwqeHGAhtHLPiEKKjqyF/sXH8IU47OvU+P0FLTdyrDM
J6a3KTAORTjbSkmJJyyVtSeboqK777LBS2/eAz6EtoKwsDklT0u3grgjGOGmF6z0
n2J13RaMeWCjk9kagdnvb6eAI4JdHhmsHnXUyiGHt3HNYk7tfb20ORCn7sHuOb9q
YLyELembVAVsJbhn9oXUmt2AXwnkxMHHhaC+V7TWP5huT5V+Xn+16xNEvknXniFp
kw7SM5BIGCq+gD9d30DJeOdfs708TZeVLTMcfV42USvdKkSyiDOd9/mT7ctTHUY/
V5ByVVOebjlEKk6wRxeXi2g05oxrzMcnBOGIU0BNdJaY5XHsnePgXZQ9B45juFAi
GXNyaX6RRJ4A39XrHsm8QnJlpk0ROYO5Z4oB8nc4BGpHP5hu45CVMOJHGci47O4S
COB2kvWiNLPRpgjQsXPnTlZb8c2/Lr+iJes4K6ODh2y9Y6tMKTYSfV2vGpTLAKF5
eMt0BzIDw1GzbocbtJUGPxq7pmQgkOTgT7s7AbPK7DwvFdTTBikORk1oZBUKRukA
+mFupUYmN00mc8kmbxBIdKaw9e9YqF3VaMjy0/yZmezqYKkVwyzqlhm9dXQdd4fJ
N19jxDowoBcetzxTIVNm/vUuluWcVN61oxjy9XACTSz512zRUcGMfk0pSJpeu0Oi
yPT6eSWZuBB20sXZW3qT8Ga8wtbWsVw/CFSM2UGXcGWnRv06Qjv8aXJBTWnQreOy
P2MwEadOS+KVsiu/u8rzN9bA6R14+Sit6DeuBwDlscy7np4PArYDbv8WE8dXXogy
4dP1JKiRccmQ+9DUn5SMjDXnBqaolHuYsYhFYaq+m0sGVKgN1X+09ZX08wBa1kMW
hYKotW4+ofxVJnidXo/3umvR5thSPwIiOKwFfk42etewMt/UKx/xVOqh1HWQJ08G
Ap3ePD3XuPLgXpF/7IJwO882tL2ggoqaHpGRYF42W1QheEOZFIcrg0SPox+SCayX
hGGhd4nlUO5F1iMgYyYqS6qF2PbIGIyDQCBKviD37hFmt7LgLaBWH6CSh0UZt7Oh
Q/NTRTBgigLZVgEn9toW7dSrJZYp8QcX6lRPY7j+7NzvpPZnsrt/Pxtw+3wnTFCT
Qpo8v4hH5ipCqTVXooN2NKH4bYmRqkE0SAnGhZCx6L1YXizZSZ6ivD5W/H2IX5pi
m9H+pia60QXa3roHajezkrUOcAk4RhM9vHpI6zrUc2WDcdFb2mkaxJ7IYGwmHUnp
mMbO/hOHVylI7NSHi9Xe94HzPFoqsX1gyGEfhHjzufdW4k/9K8iLAWVbVLpzq/IC
dbf7AmxkHMlCP+alCAoAOUhYTf3i3667ZiEqNk909LsjJI43jD+c0gqT+9ULJXS6
DLU8s4VjPDhtHYkre9iWy8FqHDYxCHYdN2624B9LzdjgkgKsMwCOx2474FKRg48P
kQjjEPlqXltJaPtfHTuIXvPs+zy7dzFgX+Kz/zzXQPKpxKmT/M/LQWqPrHXe7SSy
o9N35lubL4BadHNgU5sS2f9lmvWebct4JxzrRlRfXY9DwiKwImmeCUI4eoRQ7Tr3
Yz40Dx7edVSYE+zVKF3uLr+/of09q0zPZjNvfzyYZcLrG+qQeeQQyJH5OOsoO3un
OgnXIpN7NpoZR4EiH1ur3aU0IoEcpURztoOHju1+T9ntkJOMfA6l97q2Hw8LU+n3
0L7V7dtsbqKV+MADjIARX1hn784wwzj4WQVaXd9P00ab8Ca/JFhhB9m2TiC/e+3p
P91sWZpp6QKdaD/5izwT5NR8z9llLa8hNzOM5F7QLJupDBct/efp38FPAyO+IA3y
85UxdodjKZ6WRKdL3vB74eZMQmx5eIVjd5ObYMzvmRGFC0d8K0CLTgjoIfB/cxpL
EOte1E/hgEVQm0ViXExsEFi8fXGU1qvry/a2iN2mjtieCZaqJYbDdUxXe8J3PROG
xTSCy/B1nbTmwGqL5LEXFAuhGk6vZLTjieOhA2EWDxXL093IAjt4xs2ADF2P7ezs
ZvuqcsZVRisiSo7MXz6+c6550Gux+BZsTbV6PboDmDg0kyzYk5fc4yGG3AnZo6ck
UqqfNoAzn5vIhQWmyG86POUfCbmFuUauAv8BcCvSYpotrlGHczyRwOGH4a1ARLf1
uuznK2VkhuMA0zxWOfL/oRlRy/wBvs5nS1CM/udHC6qmbpuI0/JYtXmgW8PRX0P9
viO4S3gSvAMDN7Jhkn0lsUu6YtHFABVIQAcHnP07jNvd6Olg8c6yzUiPiedPrPH2
zIU9z1i0GHielZMfj+bMnNHUmjeoEI/BAH3OImzhDY9j84bgg1iFE8QYAhc+0Zo+
/xoYh+HOvdXoTlfdXQ0ExdcGFa87zhD9l9lkVn6R5bennzFJsb5I0aQgMplrEgGA
OAqTlG61Ivrz4A5i6cbIFsL+iDULqnK3bvvMQOUT02cckurcBaaggj8qNOC6lY2+
sT8Zq2rai5Yc15vC673qPVjt0zr83rNR2XeU8P07DCdxSZPRmHB1urIQvEsEn0Zg
36Mflmb5RJG1RXC0HSm0tQ6OsQmFXPR7PXOPBzEK1EgEW9tAqbUZh2T3xRHTmrCM
hluknFD4LFw5wUGQeRkAsqTyi3tQhd7csf4mrK10iYAqH/NAwfR+Co6saYgHAFoX
/havrcS9piaXDTejiBjCOXynJjBikcjDZNo2Kb2Dc+jT5rwiqAskz5e+jBqvF0Sv
hwTFRCKZamRRKovXDZrYk6632a+/pX1b1ThjrCxvqXnTaVcDR5APSzUrX5gyb2r8
91HjnWsIZF9VGWq6WbKi7F1eKW47cLzuKstBuHgB16Idi2KrUUHmryEujSvUyuSg
z23bg+99qMWR+Tt1HWYbcXQ96DnJ65lfVRsM4n3YsRq4YK60zs7vqWnmsnzlNc5R
vflUx6S4ezfW3s+N4dpMDgKQ9jjWeV+HKBYmAQa56bQXwVhSjyyZXVXx4J963e44
S3jahIiWK+xhw/sKYNb/z5BWcffmaioEPy2NfQwRigx1KIsZP1aqBoMuVeD/nGs0
VZRyo0FZ22ASdteFfv88G8iplhGCZRIXU9Rrbso02vei37cG+VpM1Vr05LZmodku
/4ZxrnUGkESnkSjVCCbKOZWL8KjjOHc10hnOpvPkI9bzmy8a5abVy+E8x71b6Lcj
M2WJ4SwMX4v0ZJPXPi/OhkdrOvodfYN83xifLsCBP6kNRTwPgVr0Ze30hBh7TSfb
p0FGQ4ealq8zsQTOH2Lb6VAYiCkCKoTuwOCMhiv/ZE9Fc8xgdxpVo7R30vB1oos8
n0zRWTAMcdpoaalhhdJ1F6Ba7nKdLQ6Y0SCxFgfk9j9Iisb+1zB5SjZ9WhTwuEi/
ZP4eiVrSVBdr7jRBhUTbfPQeiy/t5FD/kPv6PzNfFS3VFT/Hg1KJffo+MsnUQdWE
sykozx3Bnosi/5+IloeAl33rgBZosGLfOf6kTSVgsxbghPAAZwNzadZLeeYxUnZs
IvBok+zl3PPvsKkfcoS5yw8p5K8GZPlKrmwer3c2LGLgnlfDLi2PumM4fnZ/3Kj5
drdBEYvMO2lnJBRB7LLPAJg9fAnkzwrzZhNtde0wsl1tnGkZvHhIGBWtQjh0zpUe
yCV/mV+CRWVMXMJXzORioDmdlbCU48+QdHrD2Q7vA15b8/j4nXGiV0vqAmfcWaNc
ghlqs/IhNNZLE3rhP8MC7HWlFiMUAGBIbUO3+MDBNB3WsPFtxBub49CXoWL7tFtQ
rfUlGdpKle8CGCzrNFPBrVpX9Pn6ubspr6WauW+U1oxLa0/Dl9VmFOFUY9t4Hkh3
EdkxlCPnvAqwVdo3TN7nwfF7EU9+GSm4++ClME6eUAKNnDVHCncP0SqZLIDvzjrk
4+r6xcKEy3nlbFxfSr2TKYJX1KAdqq5mCHFXCmlzYSa0+DYl4GXWX1iqwZx1/t+p
a9D6Vs6Sxgst3qZyBAMyK8/PDeDUpTeRLmSS4+itudCBO9vHvZmLZghmZmgyuqnX
1UM73I5cG0V8p9bO/jH33LyKkx6unum05j+RmCF4mFmAgvlNluzegZrw0wiBti+e
v4X4qqDLMGJtWz8+HoaAA7qWpaFBAUjysv9kVMo3xqOLM3JmYNAFnVcNl/9DcB7U
plfQqc0iz+N0U+ZuByM03ZlhNzY06UwfxY5/EyRgvCBJWx++hc7g09X1euP/1vg0
sgFZz3y4r8OGqqJJKNGfefP7tSdTPGs1I3PmQoiDHfiIuFIq9ac111vpDk6WIgn3
HIBZO/l0RngN+RY0hewYdBhHBKxvLAgfecOvgaEaWBzX82mI4stkDR+BdGVvMlIo
L7WwGGOIXciIZm5RSaGDNil3oRI66yYN+qzVZVtJrUNnnBtuSncL/8+YE9QAycFY
AgHN2qDjrP5MqffqquNgViho4sw55bta0bt+0j05XkjhZGaK0pr0NUZbjGkWS4yy
N+I9Ihi9Oz9z8ZABTzPfgRsGU0jNdb9PHHZTI4L5K3B0p7Hml/emhstJVLaeNc7e
N6woUHR06ro+m2s4XggQQRMJCWKfUa5wTYDHf/LfO+WUoxo9kZHWP1FE4Q0SlVrR
SRpc8N7b3oou6BK7kIHuxAwyAUJj6oevcOt5GV7YqxzJDO20xAuLL/dBIEl5FHbZ
+oVRnMyngQT6PSdvjnBIEmVKqeNVp0stNeBIWu+7BEz8SviQWGJER7eLKPkj568T
N0l87ow25Xz+KQ+JeHxWk0VOEiUqlTXeGtsSZuEIniZc001mshke1X2y8wvk66kH
/S2GtgHTvA6xshpRvbJLo7MG8qQZmOQ5oE6MphSyDkSR3ILEjmxd7VNtwC6Zb3h/
P4RC27qFqfUnmQj0L/WqHkjY7Npbz+hRbUBmrnwNJEC6klSg1zVwATbmYW8tyVY4
cDzcTw+8+PS6z00YvRIqTt5nm6167pvmMZpWnujNK6ebJQB5a3WgN87m/XzpeXtg
u19eoYK06myEj2HLMbmRdBohzTd07Owvtj0D4FyylSyf6nEzlTKZlxMZahpiPGMc
Silb02HRpY/UICg9KIUh8ThUyx8CBJo3awmeS5kgNTvXkWSNkaQ0TzarztZsYpU7
lzGh2fheN1t84mL4+NWcfyoC3f2ZAH7JOHJjriixhxXvAgRl/5XMaNQIjq9yjmKM
zrnV6aEG0aOIDuz5ECvU3Wdk/g4gLM21l6b7QUde/48q0Fh1J/PVJUV39q/yHgRW
KZp05a1zaa1+260Rb95mWKiPaIi2MZzFbiUc9RHVExZJD97BLZkVNKipyf1cHnnT
SnTE+UgUwsPMhqkAuzGHbgegRNZHCZnTKaKbqpTXklH4fdFkpOcKQPS3Wg8vc1Aw
2/JRdonO9Hx/HMTNwyDgWivznC4E1naBykRYP1sMqezMf+mwl45B1z5kIXfnqYWX
AJbRxhYR/pJL/YuRt/uI+DA3b4kLh4KU7iaBdR9Q6eIturVXnXVLP3VaBU6bMIpr
XdPgRBNcWPys/ecBmQsQ51s2z9XlyT/fLmkfxUuLfgyeB1FivxFqToPFZm3sXGZi
LaTT19bzYXbikkiT/J+TQ+4VWqyXJ+FBtGpjA77eo3/U8cvNRH/8KzkW+mj4Tvff
Je9ZMAc1yvtLlqse12JsKsxwTOTWpQdkroLlnF51EL88jUlCNeB3nq24bng9TOY2
TjH1WGM/FBEV9/sIQDMujV4HJ7U2QJX3Mqb17eWkpiFJ69K/4C5h8CUFD84qRyct
+u69hkwNPNuMoDADD9a9Eq5VGdCCUtWy80fBQo5XQaTUOprSqZQ806MwjKzaO6FW
AnxI6WLrzhrOX+9lk1I7LbKZTDh47loj4SXh6AeOg6s1LIx0UUyVL7m86Ld49L4G
QJ4oNJuz05SrnRqatZW0WtCMHOtunvTwW3U/RPSOul1fICERPSo51/ezMdQ2Gkex
+xf0QiL/jRTxVcK+VoymQFlZrR1RrhNz8RA9fytOHPI62/rr/gDxmd2hvVxX1W2S
Dsy/B4NGI8JreKcq3UGmK64K7BnhFbkUcFmwEvXTaLzjZdJqFSmI3RWb9iAug2b8
rWb2/H739saD/yC3V6vugM0VJkJ377I7HyEL4EKJA2xI0AeK/90vrR5aSaIMbKGH
+yvX2N5zMBglwAUIJogNhTRBveklaQo1WUZXQIDBuN6Qp/P+rzHUKjAJjHWEUYNZ
ZmI1VMiWXeTOgO+ffujVcXhiDovS+5gMP2K03CWomeAsKkqEQJet3Y43JyCQZAF2
jG8TY6VgIPf2Yjd42LXmdPrk0osgtmeQjKcb0f5zJ3hlYx1s94C/rIodXZlxyRpO
QWdANNfFi4WPXHjvBhk0N5i8gIScr3lIpHcSXC/ZpJ6g1lG4lncFrmhxCQgpsE75
KeWqgDt01Bxaf90hptjxsJtNrDL97ydAGHQkRmhQ6AIvQXDoYrhSmF/lPuX4WZTC
jAPKqMKFs6KgyCaoiHGC36isZsAMILl8meVFd3YjIM+CYZeWTF1Drc0kq++Uf9sh
OmCCnVK4PGrov8MrZkzqYYcEVTcs5rDBZUxQxOf/HCoPw7aOkSdIoDNMqjVcSy68
WMwcmBsEfdWD/IOyf0Y1/Ou0ktdPRXDJaK/OxeQCtZcVKc4RPsKavLRLC3ueMkK1
P8YN/bIZkHXD5/0z6ooBKOh7ClIOTqu6QY4eoZhPitm66VBDc+L2stR/HKX94ewM
n11xRNG5uz2r/ZSqyg7zy4uKMIkhdCtK1Dmhthq1blBi3fSuKhBJ/Qcf6L4cgAj4
yTqKt1vjOeqIZYsGoqsDfKjokD+AyOldxbaA1gZN11fZkFuZkoCAh5RJpAiWMh2/
JbUlVjRJd8qQHBSZ2Gw7AMbHDv8cHpmofih2V8YG2LskWmgcoXMQektQliwwNdnL
xzRs831BuGmI429T8byUKZG15MgWuPCSUXmCbX6B+doEX5c2xuQeRFEDsxhKkZHL
m0D9J+7wJ2LHVmKOfiTWNQlgKGFNmNumuPI/2MM0ainUWLEdOBoDJ4Bohj8AjIsf
NxrllG8F9sUVGoQnpL0LKszZ6qBdbuqoYh3gFqL1Ja7H7drI2hUk4Yxqa2IGsfnw
U/qSBIg9GpP0B8iKkjGTV5joxz+exVXWkx4tH7MIUGtDHHYX2IKWvOSqPBQt7IjW
IjtubEm3zHYbgGZPZOhfI4iqgVG1skZHbwh8HX8tQ9tJT54qklm+MAHPWC7zZC7o
8Lx3KWLl+Xn4oRJMUkLK3GevWYpJEECjuWz625cBuI2cdUyKWjrA+raoeCXgEwHc
C/S1t4HoeU3ELHXwc8esTUrCUhoWPOsiI9dJzSWQ+oEQWo+u3N/e+mmv+VFiRtde
13SMxYRQg/mv2gbQEHVJZ0hMl4M66yf8MRLaBq0EBo94AJvSjrgFixXVqDyJXulw
GgUYs489uYcVORN4ULaqPwPHVd1AIEnWUGLnb002RD+uTM33vFmTfen8i29ADDlM
fCcP1i3HiE9wtsbzfd7mznBKAE2lHSYzj/rcU6HYmDOX5C/Q1kGkpCsqmMG5JDsk
37cussNvUde808WTT1lx14Kadyooa1QHhTBIkuROBQDByuMLsCUrGzPfW172/GDF
igCg0JxPdS7928tbvq8Fdn/aYSF30llbBRR7Fl0tMy3KKI0w6JQuSKB9MfAjrMyn
CBHvURsODcxPfMYjBqyBcs3DS7a0+wE85L4b6tVRIuAtrFxNTYI2znW6wm7l4Ndt
I+tUHgiYoxnfN0PC31AAlfc3QuCMqjQgo4L0aQN2s4ZzMKAPLldD/VAPrHx2qx4T
htVgk/ItPvvD0CGfN1alBvf44hgREAsvbHVYaKj32TP2x4IrLe3dhJLLIUTRrE6T
QorIaaDLpeATWnSev3bsPV0QKXPbKubojZm3nRarQ0felIRlr1yN8sTy8dZQUQAZ
atJx++FEq6u+yqVcqe/XKijtEUFTbC1W/tMsbAfKUVK+/8nUfy+qG0FLPORnXLWJ
eT2U6V0JFaQZWrxcwta0MSMgCm67qOPxDzDmQc6PdOAI4s720QSr5rMpSw8v3Vbe
Tv9JzLyLmE2/WY6wXMYuvxozfeV61R6weXtUKlQ01UhADq71RNId7Qv6jmbs6Hxz
lRtrr24KVGF8CBWfZMQTO/Gxn5jH22dBpV0U+qH5pUiz1IJQkPoA8i9V/Loh2Yt6
2DdlILqgYV+T7wWObkmD2mug8KSdBuuhqlA/HugxNWjwJUO1sDc2mRjMBF2PZ0BS
/EAntdwxqulubCDY8YQi/tSoDgvD2mLNGrxZbSBuozFzj4JRIfVhQcaDkbUJQE4G
8q/m1/xsPR+pWvFzv6oFE7h1RFQPqgL2dFePjgn0s2F7x2aaURecrqsW14DsBp2F
MhKWc1Uigzha0BKg+nHjkBIhsgKCLM8S4pQde12Wlzz8bi2TfpXkqYMdnpZT1d44
N9uqJ9ZRT3jWqRgn4+3op/U8VnqGIbF+WIWHk0TUa0vzarEjakM23l1PC80BM04z
moUdMmF/ou9zOwlnQ9bF9WLC8+1V9mcYnGP7fu6DwzMdA0Q+TjIi8IV8h1Dq/mMG
KCLmOPDBntAalMv4s/queTyKbCRsthm0yVHkQiroinStUJJXIQO+4W/JCrfEL/LH
eTx74IXOcCaRKsAr0E+UvYpRRX0Typo1E11TKpoFER6aQpbqsqBSKqxyo6AcmMT7
PVVxD+c0dZOWpcpL7Fjk8lrYeW4oGc1PKClGnV+dTwN4RevrJrBGgk22VH1qBw85
yTQVSjJd4sgVCsua72rQTknh2HtGXB0xLQwkZuWpCkmGK6eEzKNiOgnETLezw9ih
7lPxoqq2yFVLL1UHo81pt9LtjgJj4S0AKLFipfGorZ36BYNJAFk0ZuefQ6R8CNOa
PjSVr/J0GIqKrwdro6YFsbw6sNGimtk1EpmySMJf1CGJJ8ZBs8cSwcRBmz4p2+qV
qYsJTPRb4UfZjV9UiAIRJRqUkEIB8JvcregUB6rc0QAj8BZ9gpb8cUQBB4Xd8G4u
90qjN+aGTPZ/I+ZFXOPxNFPGOt4NP9g2NOoQKl33zofLx/u57pTIqZIwTTiXYr27
ePHOiQKMBNGAVxJ1tAHnQhltu9PhLZCZLA4DcXbJwcusZLDSMD3GLdm0oQSWqmJG
p3mc6YXEroL93RNzJ02IGezeDOx6Gg7hhwpLbcxHXRp1eb+iNZQvVHeZdf5HDoSj
sgP50lwx8X52pNqEy/MbFeeLVLMA2I91sekLhqTE27CMXimSCHmeSCvwzS91V/BC
FjSFdQ3/erTxscDFHgJqZIkPddoEcSe7BMOo4/1aTqJytvqN4ZQeYGGfMHXCXSfY
QlQfQiEE+8MfI0ZjS9sIEo7reGCZ2h6pq0SpaT3wAlZAhA9/UGdm3aEphVjGE+W7
pKXfWV4ah8wRnKmTNKS0pfQvmEjEC/TWo94X4sr1glhjWE3ju2ynigRHGCNNQTCv
LKaue5eFADUSxq2SmOCYlqzPo35hNRKCtH2Zb5MNYjH4b4psKBB95Tw2U0raq60Q
kEXDKCjBJXfsXH1mG7yvTyQ6+x6e/K4VjOWihYm4L7oL/eKKOPmewSUFEK685H8l
H10WL6nl+kc5OS/oIo0RVyJZjs3fKsv3feNPqoG7oSv+Ga9wjjk7S5DTZ2MhkE8v
WkF+zSwa2LPnGaXFktcH2eF/HKUntDPtRMI9QT/l0PQ5eOKULAoJmhafh9HFEJuD
Zvw/ycuuD+MjWwYrGeP1syZ1nREgyza7Mb7x6yq0QIfDD64na4qMsoBRuE0x/v9E
7pTDQnBueE4QilZaYkl1wFviQTUt6oi/oZaigf6fjvoREz3MQNndCQJlezdk+XM3
UoLULmatRYtXGQRJ7qGnKu0/p/rst1ovH+aHff7D6iesydAKSi4O58uAeT6A+j75
yNlIMz/oKHj9WtRcc8/GjOfPwfEnCOq3hsdMbzQY9hyd6tquHzhTpHlw2+jrdjj/
GTuAvz93SfnrdrR8b2Hn7aC+q5ymPlm/Qornmj2Cn/36yYWIzowSh0EyVZQSvI1Q
IcRCwbupIY5sNvtd08h1ZZ7SSNx+mFLIy5BH06A4efaR4zXgfubgTfG0wCLrdakH
UMD0+AZi3r5Sww47Z1XvnLT8mCq6ZcawEcJaFNrwsYLErr5HsKa9Nt2NrNqrASSD
95hAsdBheqNbEi109vM3v+n/yrMGY6qQSBh0sNc8kfsgMYaN53l2Rbj9hgT0o+sn
EWzRXKDa4FLHcDRfB5Aw0KHuOj58SG7vedsHPUW+mWU+35QgL7O7ixynCOcdAzUv
zIEsQ42hzr0yFcL6IbODhHeG4zifmyr9UMXZkW2VPYOhJTtz/zPoakJrgg9k71/q
J7aT8FytC3e6g4IxgynSmW1bLW/aS2L67R1s0as8RhhG9jG2yXxYo9g+Ev6NiMA9
vKr0vDduWkLG/5woVCcESabpIyOmZmh69WNL0wckKG05yuYf6LnWBXjiTbdNRIix
/Uwo0SX6SpGJ40lUpwlfBPCiMjpa3DGPFU0zQgoOzg6zW0xZcThh+6qL4FcKPFcQ
5WLRd1Y8u3s7z6KRBg8w0+d9HzvYiS1SuJsoF/LYPyB6Bg118N+Or50B14rFuERf
Ccuf5jd0FdiC3n8xkp+rFHO1i4KFmrMaJU5gS+gvAtGnA5G5EPYsdOR5vJ7uWGDL
6QaYh3swvhU/Z/Qk0SJwrgzI6RgjmRvsekTefZLtIK6YeOTknJGCJW82wFATqvS9
8VHP8ueHe3RKdbtOsJ6cFQi84D95aodXfwnlNoYrAkQyRC+/WI/cBgvAV+U7OuUs
L3Ads23ViZcpkMXNSnHKLkGjgKzmPW51H23a86ySrtFFi5cUhIW9vSF8XpRSzqGK
Ot5JB8w4wu/xGRbx8A5ryhnsgGFnNtmsiW/wAUp1FYFsTbl/OKTXBDyvaSRC9Ks7
0ZY+pNZcPg6tANxnwSUO/ieQRXOha6RNLVSaPGVIbJxkp5fYb94TJRWd4MfSwayE
D7pMl+kTIsjFNGe4jj9Vz/y/zAbQzn3UumxQgdEJNfYdHeNX9px2gAwxSPOlmZ3I
uJr07f7mE7O0rj+GAzApPucWoZ9bmG3TfLbHrCzRZUhDZeYxjQ4HwIPDZKLpbpJI
u/qspk7AY8SlRVm055fpdzowU8kPDQvML/o2VRdw4Pq7xrC8QB88CN0IUwD0ZXY7
W2ODb6FXOjlXzEkwNzkiLg3jziaNHrOPSfPbfCTGEFa9qF8742cuCqWt7QfbpgvW
455xxNdW+/rkcjg3a7nD+MAZGwRndsowsFpA2hvVqqlxf9hDWYqX2iVO2g8D8ax3
Cxpe7yRmndcIaEZ7s7U9pH1y7GhyOEK4dysBoTrucBznjMUeyMPE284Gzf7Hk8e6
T70FFUqC7nOMoLvO7myKO5BhjJmMsDbqg/hYYtfmIFnAUs0IaY2gexZ8JOxAhux4
poexSc6vq4sIi+cFXJpW84HdxVDaHlDKkkOgJKReW0GeOT/4TDqpVnrIdfL8xELF
Rrkk/d0B5XTAxFwNdlu7DbnaYlr+qYzt8BDpj6MnizXoq+UCg39P617WGISBl1e1
3GFFnDeQIbPCMy3R19T5044R+auvmoVn/fuqiyxHmFfw/matxhF94CCmQdYorqkT
7WSXJKSFVO9mc7pKJYQpWIcl1dzDFwd7OkirCjC02T7H80TaaAMsdkzJSo7XAvsD
U0S65jB9C1S8td6vcmWGr7ryoVdHD6XPb8llcr6SHEI8uS/Z2dyV7EpUtXbuzros
Myhq6ksyfhh8VakCh3B154nTV6mTmYvGOxr/ubHGciFHmfNu9/MskI694jJfX/ln
gSGt3GPm98Iev18f8cuaToUsaB8cC1Q5mgUb77PXm7ycdlP8R+Y0KXT2pSyLB1rC
fnP0i64TtRucl3IXHsv+W/T5hGy7++hraOkAaR1LDiMS3wLFOzxSMvmWtyuxCZRZ
wbczQuQP22GBSPZqPJOm1WS9Av4VeYaBwQbQoaHckMZWxN7kXxLHcqznk8T+FbKy
lY7SHYeLQTc+XN8O3OD4UAXkM0mCv5lOwcBMH0HR1nGvCWjmV2dk6POQD6au3DNM
lU0JvIv3tXGH3YdSHAxsr7VodIB0f1BGbC0I9Ubh9izpBdpQpxuzm8CXskYY8Quy
8RXmBa6tU+IuObwpMvQeHY0xV+HE3wvRpIanBtlChhElTp+iQGk3sXz1IXGwMjiZ
zul5FIgkgME3mxGByDeiD5tM9uHPYJFpuYY1eU8dfktRzfCsqzUXU1YU4SAWa9TL
UN3+3mWWtiEDdjtMybk7snC5A/ELLyVo42gBf/HKzEvNHL3nLvKrgK7LqqO8CzqC
3anazedippxhT4ZAYXr66PUqGseIQAwK3UD2XE+BR6Y0Q50+zbTzOdHNBCOMih0P
I5Ery388oLhItyV3oSSghMu19yMfDJ1zIDHtqJdMtbCYWLhc3k9OLE4rC473EYFb
zLwDUTxZTPLFIAuStTx1XV3EJgDxQ6vWf1C80EhNc/Uv6SnEu76M8NW22UFknmes
Vc7oc780t3jAe/p7gMzU6Qc4mn16cxYl98TMykfaY2SsFxlLjO9KIChSzXKlOlsO
eR+7G5s0oadq5DD5BWq1vfq4e19EUiJb45OTc2BvUK4up/vpfW/2dp8Wopj/lg6l
n+UYpkr5NmtQEqi8LVq1alq9dRu+M8maVqg2kxyvk/0iLuWS5or7kg+7rEIehLx0
yimlmHAY+16wYlNLZJH9KyC6oPsgqr5BsplTM0V80PY56yZ/SHf5scOecpUwtt/d
Z6AZn0FZgTKAfzpFrL2b1wZ9i4eaRZWAvHVcjUPtoYlthTiBcSRi/NTep1fUBxUX
pHCeZLJR8tHQq0XL0WD20vfpWlWJrAclEsSNNCie3lNestL1/yazqgT7zcGAV0Q9
zeykUnbpCg7+k6/nbD0G5IopXNZ2ggwBjpYWBdKPK3MSaTZIzrPUj9ntUjH8od+f
cNt048r1+SQgz8uKnPobM2/ZCnGY6dm9VWYZ4OqOPU45hW85E5CdAU1ftZRe5/aF
NR/0+gryzc5rc+inK/p9jqis4CukEdsK6Ubl/awTQM9/Y8VXCbiGWzjIX9LTiJHq
BCeT5+A6Y5VfOcalSwk16gsxYRNHWnuSzKBc+CZA+/SJu89LnU4tL3BxKbVdKvpq
6JeKeUeOAWZq6gszV3J2s2lSnXhNwSJYDtvpcpYTXf46U7vaW87mqCD4E3w91hhh
i1xzECSdvwsTsCISe0OKSPQS3fEFKL5aNhw9fXrstQqUJex7wShXNRZ/aj69hPpe
fEZVkAUZtXwqLzhTzNKsK4Qn3TtrgS/D6RXREBaC0NrslA/zeAJotFmM4tZs1RM5
1ntIeYLlzAc2/O/Kp9pXSiRJRY8QwYGo7l77xx4pMClbVN66VvxI3xHKtzDneIN6
x5Kc6K7UHm9tPoGwh690ci7gMBo1cWnDJGF9O5UYdWb+dJcK76IAwdjnWzMW7IBN
ppUSorStdHHaqpbfvYHBN2XlmvN7C9468zr07JrVmCFqRcbQZ6naCdGyDzz5CZWX
ktU6R1dJzxJReBCiCxvoavUjcpXKe63PxO9ZqjKJ61S1ahxcDEFROnrFny3/xt+U
L9c7jNCAJKdLtVcZQBJZk0GR5YEpnNMqRp7cbJB31m1LPrZ9CAeyv2BgOEoOYNkv
0pAhRmKsgrN5+admktJV94aJd3RoJzFSy1vpKErajscOprSvzCncdrZyIDKWdvee
3ZXDFUpxHtdjK7Bbise4AxiotXaUYJLNC5YxclQTuYqGP2OE3oc5a/i/sRki53zf
qCQRdWPor3brQM4KnskS+F/gd0ZEQcQKJyrOisVg168GBsggAgBosQliy7tZgDtQ
SOELo6dfcT3gMmYsenkGCWcPVXMWFqmTHo0542n2f+5P9XMul1tGWA32kq5UeGSh
d+DaOmeF0IA5vDmBgYfBiyhvH2UyL1pwhfn4FEF6eSa3Jm8LdI+KsSl7zbER4Uiq
mzSb4O/z2+vjW2go0JLJehjDl9Pwg/PFM6ysuZu/a2TXsLg4ulkG8ZfqWkVh3DIa
BlIfIdXhsYybMsSWwaGqE7Nh6aiZzOsItusbMwW6AOUnixDwsugVMl/Q2CFbxPnV
FW2EQA3BBt8AyuT2OnaztvEkbBogQJ7Zr1uJn+nKTBYssOcguerffOiiBYGf988Z
DBxhOK+wENkt4BY4bLkvdAJ5QxFtqYhaQdDROCthchnHa3Sp5J+A+dgVvLJXfWJK
TKukEKxP3Aj6rZdtK8I9wH2kvIYTrBRBiOoNdCbUPgah0LpV+eK4QGmxeAoQmla1
Z4xwPyJlX54GuL/a+/WOl9GLqpVH39RAzGDNp17aHJc4qjdn+ZgcLDhyF+GZu9/U
pl4pyJSZW+1r6rJawzq7BiAji8OI2DgzH9jYq5Yls6w4eYr8LpYQbu7lToskBnii
Q0lVTvM6Q8t0nqOIAVJ/c7j19NDS3o4UuYoYHPnGJZBoyRNXJ33t3ucx5EDCCRYa
Ut1kxKDnT/mFQInaolvjeqW3xVgVHu3ivtbAj+DHIpCZTPYOI5Ls/Y3jYqQQIUUH
JXlvurf6avoPgzOT7wy+nAzmgVP/KigYufpkToRLSZQ8f7KoT/9Hx9pgmf+iMfkW
mRf36HI+iOv86DFQ8U0c8FSuiOvdzqrMofBCBnA+xK7yG8LxGY5zAW++fnMFgBtl
zlaDSE6+GQ4XU5U5XEG7/ysQ4WUFTkRSggpZMjkYUljTz3m6b7TRzCGzG8hL3eB9
wwbMtdwhSHomesMdw/bQnmG8nwCIOhC9Hh8+JsKBvNm7pr20XlGaSLRPAavqoZne
eTqTiahFeEcvol7ZH7nVn0ibR3gWOK4Y/rKdExOUR1/dPMFj28xRIFig0yWFL+wp
s5rtkNEk+TtrVLPo/qYXHlq8VswFQdz3UuQzWaITibhuZ5CB5X3UuNvTzk/PLgcC
9+3pB21cNQZbSxJOkrPy+Rnvf06V6ksayi4uN0CyjV5MnTxR/GszsBixCvGMJuGp
4Qjbzuxl5YNRN8Yj5/dqaGylFdQ/L0CYo1KPfNgJXdGKrUA/VsWhdiyO2R2H5VG4
gsAib7+RIoMf78BJU++/ceZqlkTlRInjUZeZbloi3XIFq3U+J2mM9sz8VPGPW6JF
k7Ng1Q8bNYcddKnUspn5qafHCrVc5y8V6Vs5vJVH/r0PkbFQYSS5KBDIyoKiLwUu
RcDRzCI2yHrek9Rga/pPl1rGYdnRCMmQ8jnuGqeRPKvUcLJzlpIzJPqepP3nWo7o
6y2qVHyuVGIDh/TCzAP9EFDKZRKj6ZFnzka9P42U/qSDasjZPNCU8xTZ5JVwk3ft
PavqDs5Dhf/3sT/WszdVbq60d4bwVZKFDRrUajBweRIalkoLEe/Vc5Y41TKaTO/X
ijtKgHvLvs1KWPLqGGawL+9FN8eEpEIEFmxtGdFptzaqsNQSknRbHKlMKYMhR4CY
2PJ/YXuWtjS7JoKnBugPe0GKCJPAzRGsecS7uj41fTCFYd97lqGQMS4eJ+5tNwiO
9Ch5k1TjZGmFPvZtTbxePkp8EaNumH/2mqr471QUV/RzvoJYHr55S4bdaEY5KF6r
rBxBE0CiUDEAIUmp5ObMhektYO4vK9aN0tv7Egy8zvRY13zj7j1llERu3nGAjW+y
brwcvkBEB6rv+8v4fOqODXnLmOHmdvr3qDRpyV8ASVgEFW28kyiyAf4lFgMiEk7s
9P82zngEbHvZHMQDXIaoNpVeldUFEJzxOAv7LSBQfNVduTL3KqPq4AliuhH8xOoA
K3R+vyt1PtV+3skxWXK1x/wZlEMdCc+mAnxfzTMx6fOgHGvAOoe8LQADDgcE4nZQ
4m0o6wJTcs1WD6Fe7v6/JW8q3itbO+kPiuV0W1Wd8LpCHa1pz/uJmcooSb00JMQG
DAPdwWFhk7jgyzlIxA1aZTuIdzQqL7Di+6TWJywUXDf1RmZWyHOPAmE/6yPjiUhc
zYmZZ/ZTxx6F0NrhUf3l6EKe3UoXyeOQXFJQeh2nhTxZxPnawbX2ZtMfD8CaSH5g
1EfEr50F2oYzz2D7YzQRrFoy/ZnpkOnd8JMpbXMykXoG/bAvw+newead+xGfiFG7
yXKj5RV2ZfHqMZEavU2G/skT4j8QRtQ+hiZHm89EIt2rysoe4WGeHne5a0R35c8c
VSRHlLCFE6v3bhwyD/Lsmd67jCCEB7uas8K9TIAaPIdUdOi+rG/qQeL8z/idTmKP
lZvtaIDvPGt9FuhBgMtW0fYTu0j0PWdh2etZHjdmEXzH33+dqKAkuRDYT4lywVp/
dU9RZ6yOSkHyko7sRbWAxlaa+p8IXOeQ47/IswtvdhF9slDmzXU5OAlGK1oLk8Mo
d501qsswrssyoVnwrfXBQxJgcHq82IGnDKH4PxlNyZHIIjJYXiDjs44fMVMevpPs
Amlite9aVL7gkwURSff4fWDFUFpzhQXQUVbMG3g2Qb/LJKWZAgOVxLpt4aB/JCmE
W2Twwb/dVNbST1N1zQ0z5R2rmXIBdZD9Z6JBrIqeQUsGE4VZsKN+c6GyJ4RRnD4T
gJH6wIUCylVOLCUlBmb2GrxG0aurziKR3PTulrOdoqAxmAOQY70zlCdx767VqWL8
H59n/3UI+xbiClmf6Q7o/N4wkbcK67Bx9YEfd6StjyHrntOWLfWVfku2q4JRHmCU
qrA27+sFhNKQHhLJI3qojYh31qT8GjFx1Dy9hUgsg0P4IX6r+mgsUr9fxl7AnkD7
Mgc77hrSewrxLhs/THjlaT9oGtW9oA4zjgCFFo/TpNgji+9tHnZREXWsVMNUAzWI
LDVSWn939QaXlaHHfG4lKKkzNlWBsCQXhhyeNyc4xCPlhtlhIgD2CAcXt7LSbox0
WMTW6cG7Wasy14VaD6X+TukECc1AjGNWDdz5ws5mqOS79Tda1qnhr080zqCcWvdp
1rW6m0PmHdPQQcE8bYxVDdt/2vcTHgF6DQs9Ixzi+nvZnHemFn4hwwVMJqjezDxM
brT8aoLCVNYcIbHsmJqop3EGmTXvwyZ6eMwbZDv3SMhivCVHSeqjoDzR+308ywPz
wkWvL+yzSwwS+UbAxr4Fu/bEh2BrTCzXgoQKRe3ajZ/Vuf/jS+wx2Mq9rueYuWxa
BZaEi6bxk6or5RQobnngNZW4MFPgpRW8e/pfL/73miTb9XF+Wgm7aCkzGBFuxQE+
CWKy7MM4buOx+SiUau+tdqTsnX5yRR5eQmZC0QnpDwn8phG7h1WE2RBey1JBzlGZ
/lCwzwTyH0lxzCEpuN5ge4V8qpDojTmLLHrv1gb4dI7XhI75A0lXKGu3Y+UZH/Ai
Kwcrqo29N2HOM2u1W3eDuxZgpNdQ4xX4Fn9A58+n92npSmZzeXRNlOAZKPAnb5Hm
PoCm1mn9mk5DEBpwRYwc665NSq5eH77iXH+ser2irv5nSLtvgOIUgqrEw7vTZrlE
8n4NeKaN8O9vtkw23oXo7sFdzcB/xI9lFxoQUdMsvjEoG0qmau1gfi5I1nwXw/+h
6J7g6XsApZGtvFw3FZILGYFkm6PEpC/LcQzwGHB53bc0EfYJyyVK6pRUoyQAzzb5
04y+TBtdrCKGytKrgEVL4Lx3FhU6SIh6n+bZJa8aXnKrHnvpv9eX9i2nrrX/Odd1
KtZY3qFQHxiw7zyesiiFTBS+vtH0Izf+keQNFKOjINDyiQnhhy2pMOIZhA+1DcZg
nRzJnxoyWiQx0fOEN48Oz73kRqqUm9BpijBW0HQ0AoiyQp7YXYVMRQvFC38I67D+
vA26xFmvtz4/IIOZOdpXTkBaXVYxHyt0DbyhAvxxoVRGQCbOO7akFMzJq3eoeWwi
H/O+ME0yKztBqtBnuRe/g6gQ1y4SwZSdsKTcnf51mYpQJWgj+8YBLDUkmze9sdqF
UAm4y4JFv24+WlX6qZa8K51dm4uompY2GP7eN/9203wr4eIxRzRJxqgBiM7OkV9R
eECkEiTcxhvgX9ljW+rAdT5Zw74hpxBmaUY4SgnG1SajOY1LlUC7bZe5DJ6igDD+
XKyYcSiCb2oKFDjXrPMMYreSLPlClkpqDN46MjRtEo/8iWQCypTSI0/05ttenc8V
vRl29T0+rnUIvkGXcgScgR67DVNk+Ry9hr26kVeOpul/jkmgSp4oQ4Kpiy6aWMUv
DrC6w0LMpYIqa0TmMTSyY37WnbDIpbGz1BwVj4wO9girSWMk6RLY2frCadYGu9q0
FY0DqEC0AyLNd+jc7uBvM+JZESH409LfA44yeKW1VrEYGGyw5W/iUWn7zaxmLRrU
2+5M+3gPbqwCmzvsVd97sCezRdl2tTovkAf4rxyjx5aNP/HQoHWjULnHieK3Y8C2
+gVWvyEm4SXEzbIJ5IsUfJChddBCAPwDa3S9qKiDRsp9LuHCdHr57eq0gnIzN6Cq
OihL/LjYj4Qr0Aw2mZYhiO3UC9MWfs2bmgjnJkEL3ExqezdYxdWYQ6WGNziy0aaa
nVqlS8BYz1Yu/OTT7AmC22U8zHXrgquGxBVcKwJNYmX+mF3LLQoqnUGWMLcxg/FK
4mJsiy3biMprR/Kv95O7TCsB33E4HNqqnY8E95A2+GRkmUWoA5PFGnEZq10aZBpg
Y3purAYSm5y4xJi8e6nDv29ELiCvcb/YDnHzKQQ5HAm2b4KcGdHJT0OjThUuSFjr
EGdCmJpE3tn0RUuz6kAXfM8yAcanKa01d64eCCQZnWqLQ2AfXeX7ooEeWPAzAjea
/sysEjU4mEex65m0zWrxwLXEPen/p7F4QSjAE130mhlSbzh1WGx1SmALLXJ6VzlU
/uc94HlxjSIQCqy04IgC1QDQoiOICXhQDdgF0f25EblNBe3uLhwB4msf+yRAG0E9
Ls0d5CjyR0ct2/3YdVRppDF7jTTqs6WopJr26wqbKlCYoFsie9+mSG2TIB8EoNyy
Mrxusv1JDHx7PvNxosz3cL62k2J5x0XF+zu6ZfpCTRNmAo2sRbQzO+1o6lNVYj0A
5fUXI5OfHPZnHMgy66Qd1d/XTzc1/8z4crphgX996tGmNIQ8OZWODi4K0uOTT8aQ
Ce8Y4wo4XDLAinMizBTXBhikWHGY70tZln3mOrhuF8BlKonWRcWjDX6lGReKWZuV
xU9xgk0V84+1jIX8ai8m68FfGsSwQmLwHfGp025ELGQhRF+aGo+pFJfcHVi+QiD4
o95zaWVK8xNDR1ozGeZVsKw4HH2SqixRvQ4rePyNl5csZoP01ebEO9QPoadunbaV
nLjixX05tNPiMaeZ92rAFajfABZ9M7wPlhM5r/wnow1cVlEICuS0pxRSZ/IwQfpy
IMyPeJ4T6wScBkL8tKNXOs+5mxiYrjxyuilxG7PdqfaUhvEgCMehvEc6SnTy2fa1
M9xRIjw1o92+PtsTY+XGZff8dEPiTNJEFj2iCM6DrL+yBGsZC/Pg9VDZqETrr09t
sxsuYHg9rilWFzVPEHm2HPYf4+778u7jRwd0WxLfDsL02uL6zDUILvffisx5/MP6
Bf69ADtN9ATf9EL14XXWMVBrcIpWEcFeNx1xzURNN/vX9qAJrCbBXy+RcXg2llcq
OAI3wru95vwEscp/gsZN5P9FIJxJ6Y1bfPHREKSMggy1MQW8ftgVSF4494SIz12F
mBNeVc7sxYOqYrmyDYuBhNFXNIN84D9tDcPhtk1Ym9TMfvbm4ojWCJgiC6CxaIQs
oE+yeDvmBgkAuCHD6cbwEl3SBtkbMG4GGSLS6w+l5WuM7qgO4eUD18+2cJHgiZ/8
8muRWKBLb99js4/B8HLlYHHRVZ9xe182qfNoqX78bgxvRLdcdjBKaLPCNpc9zXMR
iYizgBDggQJmObx2QPi+anZusaIEs59KmKnIpbVN7jkQZAI6f5ne+v4/rrAad6zO
ppP02ZkqMC8vFVUOWLgUks9Kx10GF1hJ4wOHpFQ5eoDut+2/ODmGFcN2koLhFm0X
WKYEdBss3ecqis1BaOZJkLyNETLOOOy9FJsrgG3bsZxh0RtOr/12iKrY9DC1AnYB
ZG7qcdY08Ni9ZA5u7bNf6PECkdEBhTraiFB95hB7VCzGFGkS4epreyvxJ1hObWP5
gjvQXTm7wmWTg3X6b6D3DNCOM485XHeUKo7+cUqEDAxCj/jGhuw9odWMFy34JAhF
wyyAmDKhwdHc8s3zG4QbjGZwssgC5RsVmDPYh1mU3UWkb8J/6vs7Q00Y2GYx6hUw
USF7l75GqB3Z58kSVi6DsMRGwWjRQXx5XxvREFLLnB1xrCKqmF+eFlleUoj/bEVJ
DrhxwsvTTN5jU2AoPX8XWS7KNLzIuH/Z2UE27ptW9rz5MH7RTdTteG+7NHal2tMa
4nCmLNcgF/SLIRnzZs+yV2ozlDYsU3/iMoh8ONyA2QY53SMiQvhuHYSIqzaCGTCA
63lAmqRTRRqcZKY4LQVDUxnm6j2Ue1/5DpMYcro4VFM6Q/GLWlu/qgvMB6E2rVBr
OJz2rgjhO5G2wHWxz7I4E0vbRaEL3HJvyAL/rI4S+uAgQhGkMCfOCJoYXfFwxceP
CKoTr2sfjZlArTMyQTpGgwnU+9kh4j51lBsw+rWWNlSyMcK3oRRC14ht6VWwvK1c
sEaYIKPdqnNlpKB0/9xF4TwtgFHTjZKO25L0xDUXzduJcyk0w926irnZbsCwr99+
FYEXu3nbHx9ZkphYUHDxLFknr6tV1Xs6+ig+xRe8S5iO/gjeNr6QnolVPUcg/5f5
HWmo8fIxGXPHUJxVQLUv+zfY7H9ysCN+Tt3nQKLYE30ZVm7obGkDC5bQb6xP6a3H
fPv3QXpy5weyuhK/lRJnOkYNaJZRz9vs/tgOFU06nFcAZ9V17F6n+Vhslrl7Lnn5
s5720LRf1aYJDX+HsXqJf0BWdfzpZNPnODopyHFVcTc2hOiGFH7VEJ7CMY2bEIsY
19IRRNGKdsy36uoF4DuUpOhkD39FtSJeBKf4KlzHGgdhL5bOKzGjrPgKDWq73o8H
/lu3GgMj/vO/f5+mwVPev7oO6OjbL+nd88TsaKa/bdfrrAALwn4Y7n4KRs841uMg
UXzVThm16FpA9FceAqc9wCupT+LFZWt/rtsgiahHaEq+7+rbSUzKqVwVewgKFcCQ
znf8Rn4oag4df+Nm68SI8L8cZCu/sNO18qr8tvzcFeZDvckLKqgXMOWhaG4preUq
iu2LChAutnX7caf6IxLThV5nBM9XsIDej6tm7MccCj1RqLuMy0tMw0kY4IiiS47h
3W7/Jd3Iyb/kvjsYIbYE5p1qG+wFHLIqzEsxWkzNL5yI7tB7HRhAcgUEVAQRTmIo
pG/TuwtlNd4Uci85vQABLtAtdVFT9XnePdNj8mP3/4zgvMzEfXyITDaebc6e7toH
dMWDBLNaBbgbeqY5KG+sz2XEcp/Oe0Yt6M1v6qyJ0HWvvRIhQVS4QpN/aBd06mer
HD908o5WzOeaOJSj9Pbrc10FU8boc8By2q4AVZfFxe1G9Qyoo52xoQQ7tafDaHWc
G5zBH2po32BQE6Jlo8m3QuqUJMyAF3KqjBIvRaMF4G+Am9bSApsAL43fc5BqLmGU
8gtfyzG8JBir5g0rrwkDSQJFYf7m1HkY6pLdiVUj7HXgJieeh1HGNHaRuSmcIup7
ifJ+3x3ut/O6Oj6g8uVn43qml2+0/GCyX3XJ5yAj8YfwIFIIP/qThgn2nao2MqpN
rruAUo9no4/HWXh1EThLEgZ7k0QmfCol0yp01CznQPuSoEkl/m7FdgR9CiKvgaG+
8KC4kg7txPx3ckd73HTqVmtLpcpmgWD5EtUsycJDi3kzMkIi9pWJWAGPOTL0SRN8
I7CVn/Gu4Gfz3/nSCbuW/EbdbcvZwvnS/af2eD3wA3RUhkN6Rd+aXgGy76j8Tl9/
zFGET/2jLZfrdoqgVBDfcoE6bond1v2am1EE3TVLxk6FhIsVk73g/AQONtoI2nBs
uUThG0r83Nup+L+gWYGQnwMXHloK3awU9TArh//WPhbQVaFgyJFnBHTvFP/jWIkB
AN+52C4MVVSI4bQfxUh4ILrNgH0NNu3KiDLOZryVtfJWKG5vqYafwP3f2ahbD7s7
XdxCDiBCe92OxxTG9VQBOIr1p0FJQdfHlMSmPct8LV2UljX8s7hmS+ANuwzBSo8R
cA4xLaVnTZmPOnGK+76o2oTzldW1YC2v2lA30SSSFepfyCVkdaLAAvgw0bEs2MBJ
XIJ8N+3A7XwM4QjX7SlRhwiTbeqpyYm8+xZlIxVbDg1EhAtBNdTb8niJ4nPDYOzj
AX1fyAktRGApsK1xxngARTbMm2LYTNcA0cVAzhG1hEK2OBQBsEOdUtAaHoAOvbro
BKvw4cd7f4d83BpFHZTOE63RMzCZdE5j1t/wx4BdmpnNV6KudAoYBbHzkeE5l6pX
V7SPoxEyM47IH8L/HdfTsIPmjcSZEtpOmO/hmOBrNTOqo+cNy8o2XSiOXzxH8dBL
9oQLht1s623TdFyhRwu03dZLKYHWWyVSdwZ9eqhkCgbHgF7tlywbkalJmdx2I2Ol
5/i+V8EdkROlRcq1Th9VUSJMeJUSm9DRC8nf0AXBO1v7+U2nu9WBQwoZWaDYkCIS
0O43C0Tv/0TzSorG9jjxxj4fSKHM3BL8K6fbg4X12SBdiLIMJPFLduvgaAOwDofQ
WFZqJBW6WhWIKyjG2fs6xyZ74tte1hv6usePT1hPCpmj2jxy9I1qt1rlnFS/wIqQ
0noAb9OXWJzBDPstddjtFI4Y444SNAoQ1uDvvDeLpfxmBL7pyiFdJev6ncGzRDE8
nbNPJ49sq5gPSD2y9/uo9WoLVU22+j43ERNA+gzXbGKQGb0MnhAI3/Ud8PmH+FqP
nVVtrApXqGeXcEtJWpmMk96CW3xksFQhqEPcf54oU7hgEFvoWfWwzy1jHKoJNqiI
iGR8yLhYw4rdSB+08QwJWJLsBGmtzudXqQQn2mLMO0CoAb9KPtN7RuXECP6bTJhO
6JH+qz1XWyc1bg+82jiYIwqVGo852jwxDRPYlWVQD4xUCjzC4WSXvxvZxUIamfP4
t24yKYSGYHXM7bz+g2jvrT63d98rNbBgdI9G2t6Tql4pgMtrDqoU9kCo1aSH4ueY
zfg5DAYAapuRSQUaTkMxLZdmu3l7Mjzp+H6mGCY7rg+o20i9lXQ7XRga0yT9BbeU
HO3uZvqzH1posiS2vEn6d8pGeBSNnuuUrdt98be5VHNdejpgM6j6gIGk1TbNdMMJ
vLMzJa7Onq5eClLw8Lobd5/n5gWnjcsfkhiBrKX/Iu6zfqRRGIPBOMdwPYPGSnlt
09vTLZLEvPBSfSWwQp7YlIePJO195IxuKRzMwMJSWyuMjyFrw9dqetKQWcMRZ4PD
jT6vrDf9tzM20wqkB4pbOY+uESKQFcFdHxqMIsVt4TOy2+CoWhNUwQshJa7rKag9
ig9DS2rb3gKMKYwaHHSmjrH3QOvV88hyYAhHsNwjm9veR6+KhGmcQBey6ru6lzQK
GIr+k1xrcxmGcngKjFGNWndNDTFnCeUFAmJoL8Eg4dbX3eguVlO8276tUZTsLm4N
Kh06K3y7tTspLnvY6WyYp5QDF+Cgs3m2qS3Vmu0r6Li3U/YRi17IcxDM0bTHyEfC
jAPtDbAuVg0gXHe3J1bHZGvrk3BK2tNjObdQJDDO61asnYw6bJfgQVmmafvv6fXy
hJMolEBzrmroBSGG0dPR/eirUuvzMM9EArIK7t1+X2hima7kIuhP2uHR1QSLvHUK
KVtm/urnn/JbKiSJ2yGT+CnV834qY0HT3E9c6zKs73Yg+LgIqlM9KzLqCjPqkR2u
wtJQDLE6tE7mrkLVUiasqKATB2/Zrf28xNDIumtTxsMpKc1b1+NvoQPcYOMS/3F3
qjLAIW4XSZb8zCtY1pYTIRO8Vi7BE0R+ARKYM5gX93KUwylx+3YmuMS3vUB8a2hW
Gw/lVozsOO+ym/PAMwRtSA75gm0MWAKnqxLXELpZ3S92EjHv0YlTx0jw/soxYJeG
BopOda3zbtGRLf4V4V3axVPWR6l6Hn4zjXF4YWST+KungxpFfsBEhu03YAvngdBe
5tg9c8PtbjIhgPkmJj4cNPpToPlscC2UX18XimDDaFVDE/IippOyT7WVItekBVVs
a2ozuJ7vIqNoDFug65FnjgaQgEZxQSL4f6vpPfTE+BYPdzYcwi76vd/a5Tlrzdnx
qMSBINY1zzmqa3sGLHQqrvgNz3/v3RIdF3HMNMhc3jGzA1dTRWGUYnEWKVFOR40M
aiuDIvK11S4NTutaopnGP5BywgwaIH4bAMuFT9qVsT+xTg2QxN4dDPloF1iCnAPq
5ICqnMvmlI9eFLporw6/lx180iW9UO6LTGw+t9s1cd2b8u9ZLW+1YFNkjO10IqQl
MAfVuELM+ZB6FcqjS1xDSde3WKTd5mp/W67//+qQtNk4e4Yv+IhhhDSufixaDH+w
LtQ/mw704XKIMqn3MVE2jNnkEyOnfR++yvMXqxDmcyNMBbkTuAxRT1MNKw/nq7jy
6s5LBHoWbW9bZh5TJAqLEkjHFkOLzcaFM9sGR60pDKZd8K1Zt7i9nP+qsCWzcR1E
rY9BzvkOl74BMlA16yetMhyC3MzqNF7zM/gkNuHKcwgqmCv7TzJ68sX4aIGk0IpQ
mhHV/xL2S6qKSoav6AN644RxYCPR6Oa05hg7ofh+LRNUpgS2o1ICyGL07Qx1kOGx
2GtK5eCUhDCCXnTio7llWaM44XbmPqqcSuE0yK2sJhfO0K/elB/UdpMxm6pEJTlK
oZ//skGdPLmL8S2HFmf4e+idNmVbPt1mIq8bROTrz+6xVlgp7yJHitRn9Y9MLfxn
H9iKxT5KCiQBS24xc7TwD9mGOq4bQCdTqkdD4gG5geM/kBbp0TCwvRb8Y1NMrreL
jDgAYcmpb8GH/CdcNNcFO4tVtnxiGLYYWT+6L2ESgb24i65qDcQ/g0dH6nLLDpEd
Z8I4WrKjh9qJUfXr8AYy2aMaGCCWxHYinABFf6PQ7m4U/0AQuNhseFWd4wubxSwd
iqV6lxKykTdnswC/3XRVKkdgaW1ynu6caPKAxaVoD47mJLB0CkQoWssHIhsviJec
0aq/CkQgZw/9HHGHeSPZgxg0+1VVH2yKdcHixIUATFDOa/V2Xs5chv+JzWbJOy4L
MdsRDMvui2LUMXvRfdahFy1GgWH1xuy2YXl/xqiJqpt2U7aDBtbu/bMvg5eckCw2
akJtHplG+kNiEvpNlseFO5eoBNr9gR9MKAiuFV4egXEVCQBtre6+xR5at7JsVr1P
/nHi7PcPwkIcJLxFs38Jy/ubVYv3ZUf1suA6vinFMv7Cpi6soLWcjkyKYg8wG+Cm
mN6rQuEAMPR6hti1PrX590DQLdOELDHf7ceviq2PgzDAdfzGlbs20eCbf6E2jBu2
qmkPHIZKMG2srjj4aGjFaqOvZuqaC/bby+qYBKMVcf1PLZlg7UlpV+FotBQmHdXK
YKwtivnX14Wiohf2Hepctjwyimr/CkprO9U8yf6lj8Zo/VcsvwdXQHkmkbKQwyCG
ZBAX0mx6NJTASftcslhrbLF6o67BP1X5BcDe5hrlcmTMT//0T3ACGts2KUHR0s+6
B0IYJoYQatRjRjP66Aycd9Xt51EFwKZSK1K4iK8iUkTw/mR6qN7Kf5slzhcUPtLL
L2uVE4qP1TKSNDsnjbogkFEr7ToGEjOPI2/qbu3VBQk4w+j5BhDEbLYJI9uMFQe9
BSa2R5QTu9GNQZgZDJp/dC5Ru+D5UtfxV1Il98rSOQSqemJznx3Q7yrrNnBkp0wy
qiKvwAiEhkeOJNhYe9IdtLcn7GK78tHBHBupP1PFV3G7FqtDK0+P/v6Sk41UBzQ7
xANmdoAzQiHWR4Bq8j9yR63qquURAXXeW3CadZNf29CJOZwaYn3u9V9jRVrt+DcD
5KAmXARG0CGxorX4bUP8c9qxuXqxS6fH78amP7oTc1VyfCKI2xe2O2VJmKm1/Coe
/UBjE9qiiO/RD7oRmfD4tMk0r31PlS98cFgvwmEXv9h2pfsifFD5vZVnOA80r8s5
R+1wjzPDtNytS/lqa6GIET1TtbBbhQr8NRcnTcT3xJVIhm/PPoTCrkb9/FooLstw
2schg2yYmkj5XHiSmv7PhAB9/RF7g7gh1OU9T5mvDq9Ke/VHyXh9xvn3uVTjpVFx
sGz6pYAhHczJ5MElNWjbYBV6khoQe5TFx1+ziu3MZOr/nIN7qmelsKrPXyhcNKJD
EBHTnJzYNOglCU8Y28w1XDfFO4Jy6qFjP9Xi5XbEoUO2Z30J0iGeCmGHvCyGsYwS
0/PpLIOZWKyNgPTp3rxzIN95XwaQqzpp6YVa8Qm1o7LUPPQqPsJHjEsLy93qMBdW
UBXzfPdqAM87QDt0BymuJOWABhcPcnNyZqopvb0MezGPwQsb+5zJ+gP51EG/phK5
LdHnNJ/qnv9Fjs100xlB4PYroCDbRborV8uo3Z5XrMdgcxNkl2Kkd+BMAJCjIvG+
cUuqoAGBUTXy8pZm76fHkEU9q3R0LT/Ay4bDKpT8W2h0qlLHUtG7q+o//a7gPJYC
xwi+C5ruOSvkEsY8EnTGAvf58J9WBDiW2+E7Z2yezNsrBKgTu17pjFvAUuo7wb0Y
dI/2N92/XxdYftd826NHA+jP9lbUysXaI5opwbGDh3K7hjt/24lj6cDQu/MY68Hb
72nqwD57X5KIVwzK6wkpbjc5s2sQ5HVPwKmN/eGOJrvoFa6L+SI3UbTrLVZW5Wuz
5SmjpZs7fDarCmLJcwPjRPzcmYEQaYPUc5VOfqjQqMNoLWVNtSAnzZdZJ5GAahxL
eedSQ4cXpPxMtrf15Qj8BO5wDKq6lDiDXcBV46kjqmwTtUjCSff7qgD5TzVXkbNH
TIadfEOIXZ4zyrVoGRiacmQT8ciGtCIJ1Lh7mrEbhO+VeZksNC4cUp6EkAfAoffa
nTUWszzL4OcRC4v0kMsxUrT//iN9JXiWc+algNCNwsXAGzu6OgAAd1BGN9T+NoRl
w9PgziPCTl2XoOpbBmbdQuFCvzltJvvpZHSj2bnRJs1uO2UADc+B//pmKxqgqOuy
HGcw/ZjtkOHJQapV8xWEW8XzP9neYScmoAejw797p26mZfA11It4nIjnDe9mU1xh
wkMg68GGmkVWEDQtWbPOs2ilbym7OQxExmTefXP1NUmSRB+noGRWSACkfyx/M/xa
pVRSkhz1TtVMdihSvjxXdOev2TBW6BflTc2gXLsc/fuzByGnT610JNOHYCf2Zdt7
LVHGw1wlhShCJizQVzfii3oPSGajjHnK7tFRoiq6meH8XopiMAED7tZAaYNwIA7+
/HppFXqFfFln/FeScuPuO1K6rkMaMpZqCahM/g/IVabEJcoYYOKRLBGW03j0Pu1Q
Hj1axcW3k7zt7v+TH/kIW9ua2aMYScNvd1ffNF51gTcy5p2hK959LgZN/0DHSZsI
Pp8BG5iX1MgCQKgqu8PuRPPI123MdiqcDE8zaQCL17rl3x51sEB6/1iYAX2chXDr
Y8EJdW1JSpPiC65yWxf9FHEUZfzTDuwGIugczkHsptNOHsP+Yv8pOCs7V5pVi8Cj
W3zGKSzvROXfSuDCsbqrcVZFYg3q8pOoVTorqagQfupCqz0ZEVbGd4AHoEzK1Q6n
/YpDJQNBoSjYcwJtikp7tVTqWAu3mSbGo8zmtLOckGv2nm41IqnChw0yo0bLVFCS
Vv4fUsxGE4LFO6QH9CLdSJZgrUEnnL5WDAhLqYH2x+CLZeW24Totwf4Cg/uHe7l0
/OWXQdSAgZsL8y+/xcLppCXJ30lk0yvtDtzMtA2IwQaSTDo2j707mhXoQlqKj1c8
4bWMinW8qr9TIHjDnvh4Otvve53ResWV6TtGmt5+vqJYQBkM7Grk8b+3EuQ/IYjO
hB8fdvQAPwYuLI9RsjTQtC63o2Ln2soJKSJb1hWvIyGGynH6y53uxE08BeANJf8N
o9TLpeuBI+lh/vDG41bhbnIYcOk56mQbQanv1t3vNZX7ZOYM0a/yTOf5PQDua6xN
wNbzEIUIahvbvJFTriy79AJgaBK4/wrnIDCP9cI1Q30aLqDMz7zoisHeqnueYJh4
UNV99SD3ksq9NL0/rs5kP187LaMJcggLDJxuyhr3lj1a0ZFusS/9ctdYrKUad9CS
akuNb66SDsxB2Muq7JhF7hvzdgVeD6DX11iL9umUZ+7SDuq/7aly7jy5L2OKlv4Y
7TgErBSsooeB1bUjLabEE8f8+msy9rzV8jx41NAZeRqZGvZklj8POenNvy7GEDCj
3aVAr5UZnezOwUH9MJyDrdmr5b+Y13Az3jq0IUqmuDYQHUZDY7qj1sNZB3Wb/fUK
PtzWFmsL2TKBlSaCL/HYiTQwb6trntRgLhrTZ2HSIrlFJDkgQR8KUSg6Ka3YB49V
IzMvpdcsnjn56Q7vkm66cCijxZFnFoEFIa/jYojNz6mc/u/xBqoFyaBrEuJ+fEc+
3ZsZxNEk5yDAZs4Zl2sGMwP0qIE02QNy9f2WAn3mL+HhWd9G7Feafz+rR+HWBzW0
29+YkoI4WtLVS9PK3kD5TPv76enFRixqUhb9q8voNXhI4cX7AsX2hZ//5xjFtkMa
F+KfBWAwLkncTeCVdB65HkaJxPG+iz9RsDRbGccQCwbEzz8bW0MtsVdW6Hbcm7DJ
MV/acsqnknQEJAK+EiM4JKnGwj168yj091AvaBFoB5RyYzoxO4SOwHe2fqMzVDBr
ozJsIYNv/o9yxwBhF+3IRkTqCwUdNkn/dYkE7Yq9DYHBRgcDtqcxmkZbyAJzpEmA
+m72p9sqL2j6S7p0BnOJrRwmMati2I1i+Hpxdzsoh+s6qnqHzkA8q4T5fK50qxRd
KQPNEzrrlCHkeo5aUMHVnyey81N4q851SJg/7PaXtIs9XIJZy2BC28B3kflkiNzq
FwZQBvZMd7Y6bwtpjIIZ7NF7IID0uS356PXUsDEw1l3+CnArZUnJRFPsEAPQ6GGd
R+ubFnXFwW3/sUmnUpXAEmV2pkuERDnfcsnFCpN619FmXo52Y7CXDggrm1L2jvTd
HGavFfDbN413hDDFRy0DBlTYWxewZv8fWQDVcNqYc7fn/DComQwTTL7Cb3h5zE/u
6kbdMPtveeRf+w2B8eREen3isPex+UKlC+w+PXSy2me71bd3+8QQdh3sWU2zbPLr
yDvV2/u4OIjS5hz6QQ+MNjsdkCJJBmzGnpA/HZgHRR5cDW2QAyYEXG5uXMKCKkNy
VnsZQpylA1x4dK+0YtatLqGghLJ0aBfPU9b8eVf3ZkoHNDmYtCjFnUNp6jq/9nTB
55qLB6S4B2QopliG/lRSD+xk0ikQ7UIjDNOPtSMt4mwW6htLNFSO5LpniqK8jtNn
SyAJWIp8UGd8leOVUDEjNlFsJTceDKc9yhZtotrM1gFTlrIocgno84Gd4kde1TtV
VO12tqpsoKSVTBaLhjZacNj23VZxH79ilSfmkbGzOf7MyPkVETaAb5Ntk5VL71gT
JSB1ek9DsA1CjCDvODl/I5SbxQuQWD4CqEnG2o65UcJZHRpeC4K/VcSnNQssD0md
Ql4T8KiiellC20XLqIATutgTl2qff9xRrn/cvTSR09XW7/S6o3u+/09oIqkdK5I4
pwSoKYHIlWAFdRXbc4OkBRTovWQQj7uVRkUDIEe3i103ljYBm5Yfkok1jpV3JiTi
kAtzFZy860ikVPsU7Nxu/ANyVNHDAmfB1Wt325+sgeGzCGzY6t88EA08JbtsRQ1+
/SPm/9rw+58DXaAMQ/H+Ze2FF//18t5vQvoL894Rs3QSP/reTt3YGVERrNYO/kfy
n8ucjrb4k6NPRc48608PrqdpRM+I6rsbPmXPLbNuvZ7cM81DWRcyEnvWwZlsXC4N
S8PYnXZUwgdUTegNScbPABPdVYZmb60eRxWXi6rNgAWE+e9MXfHQnlaEdd+kZGz2
JAwA0v+c/2CmHvlEXTvSaYOyybtdWrCeCzv92xVywmjUBYn4X+HQMBJeFbkYZ+SK
DmFsexWvYxf4qN1mwZiKjC37KPI1jMEpt4VOChIENpHm2pAV+UNuYdiIAeXwmrMP
DZtFUkqmF3ZZVpRKbO0YKCFg1zix/ZXpI6ljQ4u+kQUlKY1ZOCNNdKT5D9Km6mSM
EXXfVcJE2Bu4wD1djfS1/u5/IFyCmWNzN8Zi84kKeHQbjb6F5WHoSKrt+abOUejf
Dq+6prxh08Ym/5LLOIXdWjep52b+iES51+2/MICD6kjgG++8RDXpd545ghJfXYxM
8GraM3I6WN1BNSXaf3KgU6kjcrv3Er1Tj16NIHh+unF4i55Y1Z01hsVr2F3QeIBZ
Hw7zzTkL9oxqSdZfdVT4IHUMxy2YukAf5O7f+8ESeKLvfYSsIvE+UlLMDn265d9D
Lk2XYIADz/uLxEsmMaxc+SmceXh1+wieK5Zu5ldE0l4nlBhjjGjJogBTfzxPxWLI
3uN4pEYPPT7ooUeJBAmhaCxSpLmlNsK/hBeVX1Y4hSCRjull9QWr8UVbZAU1zpSa
DfEOMVV3043eRXrOnvJylgtYhSJlY5CgaTaOri5UmeYS5gQIZrhBXjUPntqoOUOD
ZBbBOJCfk2eGa22mJrrYR8o71kGQJ8cabtQPTv9wFC4QzVr3WOdlXXLM7RDAswFR
WAbOd+0ODZpWdB/xpluzuntP5txMVhDmsAyIiA+QA0GZ/SB1RNpysqBhN1tsEqvo
cxZNV/m+Tpu2EqsxV128W0nGtMD5OKwDIJ7R02nTLxmN6NCJtpZ/rW1C5XMZjzWj
2xIHjKOS5GaBm5FjbGoVXuKp9veN0TnPFMhn2RHgKQnnkG3juNZ5paeobqniBKc/
RShAz89VvHhUSkaofg7WirSkAGF8x0XB9QW2cUqMcV7d0i090hvusCr5E15/WUVU
m+jGZgP8D5gZcNOedQssosBEFuTZXQfajOW+XEtW1xXH6Mz2kpB2NXpxoJS6p0c9
xPCKfBK8G9ZJMWU929B7RQlbzGSDVkBtHVddU6xL/gpkvz1p1uZ7HpdiL/ELdXOF
732DKehl4K28resSozv6M3imVHbXzjtzey0RCt2ORMlvU2fI0I8ANO6CzwgT1+6W
ONJuiOQIrVKFSV9JK2X2ObWJLLQaM+H7cITacMHtD26+lq5XezYbW80nNV1CGWWG
KnK4KKY3K/ai75bRj61YZMfzAoc3dkRUDfsJaf3fAHpsA0+6KMD5BjXQ4VvnIvGX
nFtAAOE+5U5P4lpil7IqyueUesVOKJxs8n8gyWnlfQV/5L/39+PyrxFs/WLyYPF7
VBL5ZYH205t7x/5xFzrGIy2LEISRUKcEN8DKpUJ25okm7UcqAYf6hWxgoREHvNwC
qXFSnvZYf967eVqGUjFPp4ol2g/NNJLr0JNlgXlEoODwbReCcIRXZPt23aDjgwxT
O1yEDbObSmTLphk+U0WJy0MT4E8cfdsGzgp8xsaSioDwvj1QqnEubFGQH6+ut8xU
J9NeNGU4lwaWA+JvM0dnVA4ys+xX4QVGnc0RpSJDN42QrXOyUo/VaoL2hFwYtbnK
KA17LcuPFpcK6lCYYLAnfohhRt3i6Ot5mUMaOUQPEgxffo2cboD/jbibUj2yKTmH
tN/1NuYjrDIkGpkOe7ZhUgznfRY3fT4exRkxyyJHWZYGoF3QJnjnXe+YZgPE0+9Y
JoN6OnYUiLcROj73YdBcz8XOG+f7vb4hU7Cwu8CXCtdGLgTN4hPiLLmFtdR0LRa7
Ufv2X7pBA++YgI2G7cK0SHZQ2GZLS3EXtduphjCSAIVwFDjnHQguKeDq8+H82RzH
64Hm9y//W7fOdB3LT4bpG6Sg530jXo/tKIzmuoT2lTIr66aLyu1MHIoeTtMINlPx
C9A1sQVk2w2I3ISNlbpa2RzejRyT+vUTHJNqkWFvvpSl6Jj7a9si8W0xVienN06G
iFAmse82H+1+/j3mFT1+bv36Wz95zIQXaCul+N3J/E2rItt54Ry8GwN+hxZUpW5i
YThBAtXeUX+jBBKdoC1VttjfaIkQmXnCkh/hG+630SD5wjHULNaTaGLiZqEEU6Nb
iwGBdtzb6HjrDMLcLOIW7Gp+FL3zYNV3U6VsJulKGqwliFkQ0m2U3lKicjbHzMUx
uIZAR3CXTPfrGIcZwyYsYsfl7ByALozqD4/ZPX53mPDr9REqmnfRxtTlWR00qngb
bTWLB8dqZqOjoJdALZLf85P1a7MwiPVM2nzikzlZwYdaAtq7tD092X9Vp4z3COM2
eKRpSYxB9pFx5lycD3SadoIdzX08beAgz/QwUJkBt17922v2aNVAvS57uMcrcIdj
4UGQ2ppx1+URbIgwjIiplSuozQkdUuONkhdzKlTOXUUAsCJ3bHCqaki2O52qt8w6
eVNy+83/pN/V4QxzihDytXeT49hqje95qBDXqFBoWI2lnLyaYt13mwpTOXFmDRAW
aN3pXRySj8a358FqSrYmxIhAGr2fQfgG8IwsDkpL0G7IDIIWnyg0hBMdDksWoBf9
ak4J8OaBzeqR8ILq9UoIiQLCxCjywfS+NzZpdwTxvg8rs/xC6emHr07M7luswcHk
nRcgBYm0jl+KWKfJrA9tC7v38mplUxdgJhpi3NIqnR8pJrl8xqEIhXTAeZCUqOlt
qQ1Rk8TgC734wZo8he/alokMtwcajDuFKldfT5qtYH2VoB4rrgYtMqwcC6xNRxnI
H/TATDosma7BC7opaWfrrHDosP7DiHUERsRfsiFNHBMMkUZ0m4xBb3FF+4gx2N23
jsN0o93f1So6FKwmZfc7lzW1XHvtbpOZnwz4B0faa/a3qqMjbPprpeM+tjA6aJkm
bK4hgnEZSw0a2CdchxCPee7LrGaUHDbzyN/GAXq2Dg1dn5lciSJ3a/PobMBGnYr1
n1lT79d0FFoIxHxUFxjBwhnBsnRkGYEm8KOw6hf4agxQSFPE0NQE547E/MqKSCI9
LX9e4X8yT3My7CtGHgTgIUxkxlFQqnaVq13zTiyhvMXLRtQcyM5O0QNcVcH1InAc
H+ipRaeAWoZk4/pABmJHUUgl8a+QGndzw42Z9ok24VkEDimc7P2M5tAZjKou+Sw2
ATc2Cb3+3wrnYFrdCNf9JtQIH3mmacGgPQndgVmeK2Dku+UH82502zvLK45gmeOZ
V+cgodZeyEbg/vswTqSINXyE6cagrLsw/t2QjgWdsAtbF9VPUMnOjJHVWiDltiZ5
PE3lLm7FUfyrpUWEu+oYDUcpNkYVdejkbxuwLhbGB8Ss7uIdxJQe60cXPWWxB5sB
s20araqmIQYPAW9COv+2w9g++kP0CS7wdvzEJAw3R8q2nhvbNMbx3SO55hmjORjb
zDWB82b/EZBPlV7sKd87RQd4HtuxLvm+1vxSbDIHTjsiI5q7bt8VEkOmIiRcSh0o
zUVfxr3F69eOEjOLhIVBFtNuBZaQz7pRMSyGa91bbU3kDZAz+1FYzn+vH+wxHyR0
qmJIpGS1q3xCdJmgU9Qqq8tSsiVdCUd/l21CGNMW5H/miOgzRXZ13o4wDTYaZKfe
mC8WSCQiSYi0IJAxlW/C1WbjvrBldF7qJ1MAs2mmYyfK1H8JtNQrHY0ic/xjkBpJ
SAAMG2zJtYThPpTKbuAeEx6/zI8kbr0N4ZvhCov1CBXUFw5gLDsIjZv9tg05t1LB
wbNzzZha8V8Nk1eBropsAonqPMtB6Db51/JX8c3I/ehEhchGQAyN71H0ISZdB3Rf
8WIR5o8kEdiKVPsR6z/H/UO2EHgtD6BSGNTeRXIwUxFHDGIBxsoO+z2poKq03xTL
jKlEL3KQKSjDPVHZFiw6UK0SvCQViyq6CLsHvXy+eSpezLxi221cbA0knQyjEbcz
7AmIumh8XqPBfwfOQGOLPcMkU2i/fqU8O8yqI3PGe+Lg+YZg3UPvHbV/mJnckSxQ
q9ptbOPWXPCpKLye8FsN6CaoSAMvJXbFGTbliJsTMkVnW8FhAcjOcDkENcfANxOh
YBYZUJY7kP0sWz1CLi1L1kn6otyEi8xj2tfOq//jPe8G4b3qi5Wa2VJjEJDG1v5d
MaxITg1BI1zEfCMbo2u6I0E6LFui+S5eHwKQOzzBlu+SXJugIWkseabPjHM+GmnC
gF0tcPPQl38Wl6LpCuQgCwJF7kn61sDM6Q9WMQsbXP1Q/QKVpldOw41qYZGdt/S0
uvuV4AcI4zVsVTYjzrrdDqidzdglDLOiEiOv5RrFcwUM0s79nE4+X+K7UuIrgofG
S3ZJbhhm9nV2jIZlCltyfvIF5yJz1924VfutUNg93ZhYuP3A7jYAJG3WqkMNHFXt
UcM3ohdls4fMs9ucnMRlNThK06le3AiWsezZuMKLo+pxmf9JzfugOIqtTNeKsyqw
y1+kjvaHgUUakMa44d1vuNZjouu6w/FqMbLY69wlr3UZI2uIRKjWc+dI79ik1KwU
IHTPWMPYyLRDkZNYV7fOwNZ38avqOJ3vT6Hcek4hAx6/09EaSYindzBsKD7/70J1
XaR5jGQ5RYLgMuBNS58XTJb9xnVoNvTrGMZ6PQn/VkMOMa+wvYe2hV6NXNCP76+A
Wo77gza2U81j065MlsakQ0mvp7R1v0I2O8kR3U6eKlok1caPI3P2JSBLHvDZ5Wkn
hWwwFipqoJT8NOO3ETnAmIqLcU0fUk68/DON3xcbQkU9DGfPIfgknY+xgVuWSWYu
nZKQL4q8RDWOfnnL67/GEnlskEDl8uj/c/rzfTpdc6Co4vaRbX0tBapcbz/CZhNj
O8a7uV7/knVjamfcJeHVYm7IuJ1Q1crbsxSUjugPZpMlcVR4FA4e5ksgLITmLWBJ
4nD2LTLsON8IArfGeVlae9QMKwhynMuG8QRdgJIExdC+lwriHjHwCl5bNJm/y3f7
3wrGqWSI098nOvsbUDBoMl0xer7NP+vAl2pw4XdOU0waTWF4dIWh9f1ofM13sTBS
dsmbuOArL03dcdMSNCz43GmcbM3m0mWeRiNGDhzxQ1Z0iBLyqjhCDbdz9cMXEhTe
80xvHbQkYuvIVGFD6NNwCPjlsD+BTk8F3MB3UTfX/Qwtef7nXndQqzbV0xugL0eS
WuKnC7+1Tdj92y0cZcKIZhqsLLfs/6TojP3pB/lx3naW5vJiUA3o/jxO+SeK9jac
TnCLZkM49nCKWacM5hAvwxf1MZq2mU9P8ALz3An0N9cOxou+1EB7Auan+XT7KqBI
bjJ+MNXu9GWApmQUsTEDy5jcAKt+RdRSCj5THzJmC11dNOgeUg98+ryHZxmrjiSO
1M2k46Gvd1XFaPNRb2SRPfjRMPww5IHlTq+HWoiJ+psWJ76jzvicyPykrA4sOFw9
x1RRMEpySlVuraNms8rzKlW77eRkW0BXzX/del3LwHIdASpJY+3xg8GapzlE9EJh
rVyubpir4ojwQyuReCAadGwT8ioNE5VHhYZ+SlagL3k8dtr/XmQXfjZRmgC6fL/g
cSf8qedU4ujntdNMlRqwusYu6bQ10vV0kKl2EkZ3QIIoGbjnlfnbUIJ+JnhcO48U
2hvI1LuuG2ysOt6vJR+pnZ72uhGO6hWyWbQjUI10YDFJOt2N1MKMOPogS8r3VWeT
6JtCMA89uOKj4ahtY0CsssEmZURdvH0bmE601PpIwxLajdoCjOTbiMj8UvrCYSyr
len/Xb36Sp9tF6bayr9gfS8Y3pp1GVBV1PfyrZ9G5rgunywg2iU33cKabl2a9CWO
6SBJ2qY8KoMwIvYHkjdiLAU5nzn5/BbJRW3dTPhpn3D2FvqO7p8h2s94nzlclJPa
EPSd0Swvs89fKLBiegWTi/pQp4pBV6Ys/Hg+26yeniIMTxM3faiXW1q/JdTT/ftb
4VWm81nyIAykfGL9+UqqUBA7NKCN/3QPLG7hoXdlkmeqCXfGQ0uEoPALNH3chXga
2wcvQRij/iYBtlXa3NCzofOYvZu2qNMXrvacj6fPDQFmd+xzDPHZp6eodwXwukgu
N61O3Zve9BNczakCZfL+8nudtKFXGBRiTYzluuXuW40tKeWYJWSY0v0pZKCtpwVD
cBsmF0CEJsdqUT+Xlx45wXhxFnYqbrhKflQ6I5sBQeZk3tXbzESSrKrtNoXb5gl6
FP2uwX9w1d0VN0JLBK9U77t0BClhqWNXSwKdBJNKuJYRgjm+KIq56Q6thHVk5NxF
H0gsiBmn3EGHBZS3ZpTU0rz4NnJQfxLJfBhoreQW8/NArMkgFsz0ItI8M9iXahXN
DmJvRI9obVhIFB+1yb1MzFCciYMJgUAuAiepn2YZODWY7omwegPsiXxr3FbKKgl1
2UO7/IzFfyGYzhOxuCSuZLyXhc3j7+WlkwfdoBgeXW7caaNerkhw0Gco5Lb1H3PH
Phal2qDcQ1w8DHAM+rYsBhXs3meFHZipWibQzgexs3FBitEK0pr/GQmao2R/f8uk
NfPqKJjpb7J0Rn98UZAgJ6RG1TO8Wgn4yedRH0dA/bLoct9dSPAkRUrgOBx+DRuv
wfJgqFAlCRpfnZdXiMh5aow0BSKztDdLG1IDcI8eJE4wGJO8dY17ebgwdLivu9wE
qJzzLn6wt60bz3cl57+8QM+howDAHccNjGTRqieAQZ176hmm/F+rZmqDSqCYuA7J
WwLH3e6OVzGCKTr1n0MXjcanD3kuJ3L0AD2kOMs7Fnp11f+CTIEGmX6AXF5InpsK
pWHqVHkSUYgNgJ48Ox+nwrqmAM0McX4ECcj6RpsYp74m5AhGdfsyVH+TvHi5c8ZX
K3W85tSAi0BgHRcGAdDQrcB3/I6OGsFQLsMW1JdPeQXFRy4RkD/a6Tv1ikIDo7t7
eE6oJCohUHAYAVRu1xwodb6XQcivL0Vl7YEzn/nJvR0xFZjHRYK78E8B1+wPoGx0
yHPpVL4pZMUpwZD3kYWMh4ACyzB7hAJTb74JzMZD3JsWOnb9fES2pyNXUJNH51nS
8gF3i3xiKYGki6rz7rRRRRIrUvjjNJZv2SOf6ImHqaSaId4X/0lEjIyCOFpaBWAj
sUZDJZlpVRQQwpYYwMs+zsNB5YfxD6/I3sHlN6eVuowoKoxkJZR2rf2iW4Bna1Pb
Ml8w/hEXX899+tGN+kWduMwraqtvmZkRN9Djt2jGWzA8inYOdHx++yxpvRHWGyfM
mSFPQIuWd21iT99vlJ2soNdWGM+WXGVKt5nYw5vZD3BoWhXfTAxewQztzYwEcTlW
R3j9iJcr+ClG0TUwErRBbSkkKDl77yn7v5Fm4NP3vzjr8z610UXEpUa/l6OxxDZk
B5WRhE1vEd+eVx++O25hMh/zQmcWqDeX0alO944x/UIGthv0YCWKo0GsR2ts7mus
k6MlA1d+N531KUROVIrQXGckb9l8d2c/GXvaUKVNKvXhs/BFTm2LMKgtB81MJU0Q
CLYy8z31t5zN7K8wdtdkUTiSn8VN8r8AiU3mjqRz8Efj4BY+LmQuUhszbRStZEpv
lZXP5ePZwrcFZtwyp4lYv9AUJ2NbD++DH9glX7Y4qtcbLx57VcllRV/WTtFjZLWL
LHUguPav8VOj4i322vipMC/ywCgTX3XmafoMujePoJ3CiRgClQacnoNbPp2LeAYp
Oa0SxYgbHyAAaDa8m6vs9Kh79xnM8uenS51spD1x4GSl2FJQ4J3Xyk1JFmkdWqFy
xo8SWro90gXMIqqk//0JLQ/Sk5hF3O/F1W7PHUt0EpBAoBYloIsV20lA16pVY23i
itrWXXgIFjAPQiB1kKfeSwf7TvXlOzfuboinI6T924Zy0BPpvm/XWOnsB5L+Na8U
e6oGDYB6tuJVwVCYqdr9Pe1cLaToV/KhgBprMo/gK/S9JDKXw8oa/IrMi7VZsqM7
k5yliUrm86N7d9ykY6Cdjdzrxa/ZoGpm7YAgKl66xMQvOyrBfKhOCleZYquKhq61
YsZzPMt0Y83+GDBRlHk/8+frWSN+F3dspFKW03BkmbWWsllxfY/nAyXWnYHlKEeu
u0UKI7sx7qf48ImFjlV1skqHiUAH64Pcabj+jIz24ev3W0jOpOj+cBfk/1tps/lZ
Vhxf+51/AGGgcKFr0pUwLcQND9Jbs1EbOv8p3ZX3kG5gCixIGaz5nKC923qIj0bC
3gseZXaIiJfm3DgBUc9+Q39KTirLG4nj/7QKG9wPihXNWbzvwTrYiSdpEeTlVNTK
MBJQRB1aY+dUTwMV6I9Qx2RAew7OJVqX1kEr6rA29CWQLRpoS9N3R2Q6iTOj8wkf
tMJygo+c+xKpYnYPhn4ftLKefzoLt+oof+KDk9SzP7V78HMFtIHpeD+a1qEY8mCV
OMy/KBitQD44YUK3VZdP9vIHyvAxzWou/up15L9b41HttCJBgIV/A5vqM5ZXt9Kc
1THDpeEljAugQb05ouQ6Uwqv0j4Xd0EDL+woJJFxFXrSs3qbh6/2GoWDMsP8lsDF
YBUCKMIot7v6wK15ZlVnUVXwjdL1fbL/sbIecvXAYS+k4kRMelElw5XS2E7dkeVM
DYy73MwRoGmTLB1dQx5ShKizVG+OMtr/N0SO9yt8xlzQryIdTZJHM/I2VOk9cR0T
f7vndRmy8P1vQOUsLF7oL1aXSPu3VFwPSYxyw2WFffC9J2+WxZFHzYNVbrAYb8+F
xSrhlQxGe5/xJNrua4Fn1wZuWxaBCnJurQ7ay3QZvyew4Bd75QraIj3j2OCIVrHX
96Ad8KD2iqcXs8GtQDJ/4kGw1DxUHcGgnAOeWn4UNvGZhKLKdh6oV/23boaj5r2f
lr02JNcaUEb8DBgEz4ZXtUuLaBP9ShFxM6BrBbsXDwc5lFGDgdZrKWq9rpvvdjlW
OR7kQBNEVLLZAyc6bcd4G4AZ3RWRGjWL2jm8sBs/4nJJ8ohcJ0GByRu67N+tJdwL
tKbRpAH95PWJC0bY/cpLmnbQkqp48l6MMAHi4wdHet8QTokTkJpknKZoftpRAbwG
Y25LNGsg37XlPQJVT4q4Kga6xpPxza5LcgNlr0bmJfp3tlU5/XMJOtM8AxQzaSxx
1r9kfXykwMur85KBE/tpsAKpyelzv58DsaxNQW0w9Lsyr7YPcV24TqRK3ib1Ybs4
8A60oUsooyA0zxL5yJ7F+cfHDzELUbVwYzwXPT/Cx2cjL+lO3xt+Kh5p7iJmfrp7
u/51JobZaDekInFcRNJqJUjnj/CTHT3dQ9tjLPiG8uDdZ5L2APdfIOgz0ZpBwdnW
Ikmv6OslmctNeRsm8q/zxRmFmNuslVnFsLjBos/Po5EtSiXxlXE0HTHVN6XPGxzx
/LRtzfZeqj/uYhnrTA6Nn9Xq5EYSqrxr5Djn9+jb9d1FyRL5DP8mOxz8OIHd03eS
qNFqhwE13Hohk5+gWzSdNERFmyen7/cjL7lI6ilmy3cFgXfVhfOOjt/t9qSP2s41
JuYNUxNzwFyEcClGbObXssoI7BPwCYAEpugjNGlccyQw+Kcbmiyl4QI/waAw7bGU
ydzBEE8ttMDpWBxeoucPAznEE5X7QehUeJ1yCnskGTqGaq1gYjPZtlpqsesB28bk
PDVN4VgMnWm8/eebrn5ohNRDzeIMndJUmZmTx4J/KwGkNrqi0tYAqJrEdt+jqrha
vqqbhakkxxMMn3p04ndWWlSVCQUQrDL2JT4g3c22N/7+r6YgVMPvwn8j5NF7udA8
Bac1Jq53RGB9O2Tv4LRJ79FutfdoYW+ozhtHu8AA7ptnFSQqA+fKtgpF8FKioEum
bwZWYEdoI2+gbXMgsQekxC0TOJNgDd9sNrJ69hU6MhbCBYypJTjLWWUH9/+HvjaH
oXJPK8qAzcc86AlPUxxgbuYDf4vY2vH1qAL8Shbadpt16+QoJx0jRn1T+aNZexp2
/8DF0k1oyuXgCSGZf+SdwxXdkRvmvU8Wz58ZrtSpXXtkZgFhHBmVLD2v8FmVmhFN
KdLx+HMuDcxU337NcwhxnlRiUohgGKeAy0lFZ+GWXZ+ar5DH4Badjki5uYoqFoJo
f7TlX3GjLUIAgj59p2DhoqESf94FdqpgZBShdGiCjlipOBH3yVcucFAcf7lS71oJ
SRHiD68kd5h5i2/Vk0jAuayrgAuEeOA8TY5HmA4/aRU7UXRw+u1yhU95uwe7dJWe
n2rPFlQTSfsqUjIzHvey70IIRXLqwl4PFPqdXfO6e/A725i/tIyeXgydn7g95IA0
BXyAXXXUg4On2Sy1kk6ZdEtTgC8SxnW0v+egXPuxt5fhzg8BcxlepWhxSuHqZqSR
ZFXR1kJEijoAqq932T0Ek41mXQwcMsewJ6RY9mSxWMmMZsNnm45H+enx+ZwxCOec
DIzYeIEYH1oX+Bn+jBjapUmgsEi4NXhWYn+DriwHXPMDKJwpKDFHNecz6NvSzphp
lxngR6ub0KP9wQXvYcHi9lRfhZDXayjQ3BAOCLded1pzXN8lFtGvOPcmCetgN7Sw
8P08HQV/0poza+Q0DcJHyc3zWHq0nK6CpfbM344NHBcZDb13RBIZQpLRLTtnWum2
AytHoh/gqBdUDiYbP3mewPh5qoJgh2SC9BNmK0ezFCFy5v5FehROLuQ8QtXxrX90
wE5xszoZgA973Ixs/Xf7gAxOISEGCzcT0ciPec3baxq46US2laI3NvfD2vhOW54b
bZ6JBz4aD4bJBv03XPg4DwBWvh278oWdsNFzKJERJavtnkd+05mFn8rmg0XS2tUy
grw0JKZ8hYITupeyKWw9OnOQw2MTM+FqBMhAFG4crCplYkiTPNL8Xf7R6j9ahS1F
VYqkCipGFHC15SmH3PQIDJkq5whWHKFfKlmiSy11wJJ8HY/BivfN6JakPTlNzGZW
iGdd1C19JatHiQlgl3ahl2CtqIzqR9R1dWstoU0hmtfrttwgBzipsf9pu3phwktL
WzT6SmfXmHo1A+L630RfQNxseH/kA40M31gJut+3ID/wrYcnyfL0/tUQElORkeDa
xvOf3Jbrb0yrYutFHaMArGqZgne5eEezBMgv4HKtMNXLyHUtdYnu7Kxg1HHLkz04
hxs6is8cmHYfV2j+qEM34vBZMygDDGg+03mQAe6tNVGYu4oenP6eoUiiFNjGBohA
5GZnwHzSEQciQ/zzAosPCry3Lh0v+XiLJGGz+1MYM18EL6INcxVsFOEKTissAi1a
W8ikdD4CPm6wEa5KVgKuyBrHTzOuSNJExZfhTgId0WonO+eGVzL/8Dmr9U93GaZi
FQdCs4L8jJYUsNK1IFMq1724u9FmSJtyX20L1eTOpr4yQA9JjcQDeomysMX2/j8+
5YgzPPZQVrWj3gtowdYn3nruOlxDC4+B/oUr94ZdOIEwhcchZ3AXNLlSDylb/y4d
Ro5J72mIZ3AHf2jBZ7qXckNWDYNfsGqd4arnDox1RI/QpiaaZNBiuxgXdvY78Yn6
XZU3Cqb7Bsvqi1HGTTFzjMAS6wXlI+IT6K6kiQnM4xisUxhKXzQoufYwuECopon1
8eziDD0s3/m0ytEfDhIZ70YlDCdxqC6bteF6l28cDnkKH57YNtKmpxiP4/zMBQmK
BQwNsYJGCjTOkVgzA/xAhs6b1RP1Tqe5A62UVcGfnjADdhDWphTz6DTt8EM07CZl
CQ+UFEGjkdec7vdsOWE3sD2PShKyNGzTbPtBlVMvvStgLbRkG7pWf0EM+rOsk7b5
rdL8b5tf5y66JTvYN8BYodwXbxdxZEwHrsh7g1CXEOTnHv8Av40P6u5oDnu2BmnS
u2/wGDULORaDviO9dDlPMXGOJJ7Pj6cbEQ+95arm8Trlzy5lISdPg2ojQ3/+9CmI
OnK+HgaOgRm0ipgxq+sGQ8X2UQPGCBzluiyBKSX5MMIg76/qqmX8Y9JkqdfvcfW4
GM3J/EAvhmogk4NPyAx/+rAapMFVZRpCD5iBk5sJ139NltIP7V61JDp3mIToEzcn
9wHhFD5nYcXRsIYmp3j4fuqz5CzvKQijFvd8TS0LMrTi7g/Pdq9JQfbq+ehbgn+d
r2sUDYaPfZlrzbjSIQir2fSUiymSgeKydQJq4p8oYFalL9h1N+JKDYl0wcJ4O1VI
1537rhwkCshHv3N4vBzrjO2RXo33jjlf97upZDpKVYXC72y4voeCRJqy7ft3lK5E
5SSERL+zxnacsuuuKCTjQSql4i6t4hQCuC9XCGwv/LA3UwzMJxseogEBv5Xcfny0
6+dHoRRIpI8iQJzLEJPdmfWaupeEuqNVzApd2fidYmFrEnLLjPb7xos7IE24c8hZ
sJ6sQneelyUqy4+/Kl25eKikKVZWsfNfxyWCR44YVyKtJyv0Qw4UJg7/nEv25H2M
0ctQaDEf7vEd6PXCUIAckfUzuo+aq22vEh6w8rrJWnDuaHC4FYvUbpc7c9bMPJxd
TT12/lX+RMvQVRXa0UHRubuQnLxv0ycO5912rfzLD2pUJ6pP8TDoMUkz74pYvJW3
skP8vmzC4EfAIf852c1Fth5qIbx8Zv111lTcTq/WfqZoMkQ4v5U6yVs/hpA+VQWi
dDm0BfBKcxQDb7v5wefp/LRW2fkIaidm254GIndEUyaG9rof7H5IuLNY/q6kDB/S
FOZ6Mi6aakeSE/G6zoMMZxMGlQMa85BBISkMCloBNSpQUqBLhT+fwWtYWsChaik/
V3fimri83DspCl005U3EDwDZgBuyBoNcWHXNGwHwNnwsLfRxgQ4FOuxZ9wvpQkLY
klHvXh311Sfk5+lUf9dtkZvxOTl63hmApaJouydRqRoTdRzcj0Fpf6r94N4JOxuy
cgz3soSG0Nxyd6OuNBZ3qi1OXeCmJlyEkBj6yo8PeAmzq7Jj/SNUoQ13HHN8xYGg
iCnOKD5JvknrJF0hIvviVmu60j0IgYvlmA1Ep5T+/G0VlcrxNicDc43mNlMWaCNY
G9cWAuoIyW7fCBs0/48FlNp47ZdvgL/JOcAlmSQJHe7wNAnHdVLUBILGL3YNiLr4
iRJHCr8PgMReQGCLtD+IMSl0cl5AY2ZJ3d7R920fL7MWQSngapoyAR/MQAbPV4fR
5Fv4Fk96xXt2iugkuuKanGljoXGbdERsMibbcTLYF9Vu+ECwfrPNcPwoMyK1ZQxB
A16B2JbVv5XMbFhaNApoeOkJdScbQPkbGBgHOx5J6ubdv06wCiFUZa6todxoNoh3
+yCsmrZIZwctOR4Ui6ifJEr8WzG48APR4A8YPTMsbxNjMkJGhakN94B5ryyrsMNE
SDx32ruAOifEP0cQhyiHiBIgXZVPtWMa56RVdL4aN7D0wtwN6cCUqwewK5PPnGwp
LF6m4T4TJEuU0NXY9dYL3VE04VNE02+ASc8mYJKjWZPHaG6uF+B5TTCRIJcGhcaU
cd6REKGH4dvsQCVQ7SKVhkIHy7DWuVjpnr5Yc9MeVtEPZOq98qyattLqfR+UiORL
0ljj4V2IR2PJdtlaqckbiq9b4f520iqvJbThSp3tnrIG0RATb8p2IKCsi9qYxiWX
2ioozuL+kEO1pBioyzVfeeDux8Xce32AlcrVDri/NaLvAWBdPstpJsPawdj9U54C
S1MKqcdbcuJQ3Slqsl2rBmoLXLa0USH9O4jbYWKhyifXeGar7CtDu5kApMnzGf4w
LDgW2KWYcvjlYtGm80QTgV91hsTxvJsBij2BfGSHykOxjp9h8wK26a2F8kH123n+
iGZzWKOx4xL8a/L5f1J2RtP+fCbfPTqMrHrSGT+9+kN1KpT5AWM/D3z3ibUswPEo
jraC9H9LnOmG3bWDJ9YvXhj1a3G8lQzXUvNTIpjoJPtoBQzcn1A1WEeFWIe0kWTE
n24BLIrzQmoTB1wVPDwfMY5oajeGzWeRZZQ17L2IV2bfu3sXo5T7BFqCRE/+nkSI
Nn91o6YgE9cfAFGdqsUgv4emz5DvdkoCZBQnNDQ2+r9CetV+F9KO5Yi4plXu6Z63
1h3Zq16XvSDsDkxOTxUgjt6tWolCazQ3Wm+7pHqn5p+aTmADLtfz8cL9a1hhcLrp
W7O3b92F8bYACOv2D6rea8RSc6h57Axpq90iWQgHw50IUQnLFyUi62kRH9eDcdJq
HjG+pPiXdV5yPcht2uu49D4h4yXnm7j7ievfjqBzYY93Jc3QSjQaxMvuXZu4LUr8
4IElEvzHTFJWczTst7yF2FqXtAcQo5vzIWyzTWW6UdWETZGgQqAXN21L3ZMbCS6H
eFmSbHWtjfF2/04hp7kljvzK/CrCrFzzB9t9qL4sufpu/zAM2+aslD+StTy55bjX
Nw7ITtStn/p/5mI8gBlN4KkGyoOJX4izun0TSiBAyFYzzCpxnE+g7HPJvtW8c29J
qtQwJmz2OHeVSNBtbvLC0fOcL+FhIko08TmOZYXe0Pq5uab9DdIKrKSYe5FxgrfM
pkkFtu7aLopm6AgIahrWqGLk4+53s0HokHVzr9Hi0u/YugOYXWMJtGDgrFQpcn06
RYTsWNAEkO9k7vy/cE2AAL23ZsMr7vnZFQdIwouOZnm+N+edqAtZENaCkW/EVRtD
a5gp5aR97aB/js+jNPxuL4/12fJZi4rcJQBbXnX1N5QIJ2IQI+V078rrijkFZrO1
F39lOGkGqKHAbRPidwPegtUGdLnh31rVBvumfHaXGOizXzIAmR6E0Yk7ZYcQfJbA
TbnAYacABNOW5EFPBEnAJ3A0SoVCVCRDXxMcwxyDuUX9nUZILfVAlJJNfKrhnJjh
gqDJwn7m64UmMVnHYB/OVOyChmsLG7tJuLqVOHswAfQFodcSG9DTSr2u6K6+JPzj
J7YmF/0sD7LogZpetmVa+aoiAIzta/7PEnTmibULvGQjnhKQ1JgQIcrqeqxWZY02
a/x+AUlCsq+ZRj6c5wXG8M1KsVQRtgnGFGyBVcaSM9D7I2WS7d/NZC+ZdHJmTKHa
elkVyYompDnbOi3cM0L7e8iPTHNkm0AbMLSHmh6uGCK7R5+u5t3eHg1M+aKsOq73
aSHentsXD4ldnaFX1CjJDlJWmZnAKwXAO+nbfbuE13HRKmgPLeXYKpXwaN6Qq5JA
cFU9/oSucrzrUkRSfQNDxCWQYwR8VIahvROGLmsZtepoO1+db+PNEUz6zCjehIHq
OUHHeq/J2z9D2B3ztlBbnwXFEBoou5vWH4+14lRtXRylTUW8Y7jNRjFv5WyFT3eh
nztF4943Nfr84y9SFd+rciD60KwuAmXTOxCvoi5dcdIoby7ciYnji3wootnbpZRq
GiIkINd8e1NDi4ugrYq9Xot3c8Wy+nqCplJOI/Rq/PF4Zo7JNbGJ3YWUG6rcWMbh
sDm0JnvFIFjjpUhiRHBLkyjP7MrMabv7ShW2KNwkN5ycBrNIi+SPX5I6EOvCKMen
rT673VTUhBEsXDBTZNYVgWa+mqNJgS/EttwdJ0QydZZl876qL2H6ib8lBOY0Tq9U
avY2WZdbyLEgWI1LJimyCVpGX+gQdL/oIJhrVx/+TUw4nq3cOjlDqoJSikdiMgFZ
SNQ9Xgol+pQ2+2NIp+p+npy6odrY/7fX/17pXcSVges42R5bKNA9vp30UCiMA8a7
mIlFZ3X9MZ6VKNie4BQ05LVlLkeoc14An4LmXB4gxvol0tl/lA7QKDvcpVFmj7x8
w8QtaNxLm7GAVbvq0SaggGuRjo0WMQsSVixgoDf0FZxayiUH1lChEw/BSlq5aSOR
e465n9idbvxrVbX8cOzdr/2McI4js9lG4z0kKwwDUxRKD+9D4ZjjTAHpFVXo6MvI
U0A8nVBR6Vxybm85NStTsxthYSI5ha4ahwXB3hVy33JaprzvW6/yyOGxh5wuD+1z
r8lXqdmyWsDl/JHkR8RGq0QOB9yJmQ1zr9crIy4zZlFMmlprpVo42olNTfjwZBk8
AEf5q5CMVES9oyEWzN+Qre7ClJBoxzpLl2PNQoXWiacf5JW5hHMp6oVNJJvvoUZ8
VdrvglkF4nOc+Y2y2TjkUdxDk/fl/BuaVnGjE6496RWrbmfFlVp8IFddTMeUVlFc
2rDL5LJhArLR5DD1Dqr783G+tllBXGpQRONxhhvJ5u7NXGsNYM1XEHCjN1wFlTZ/
44NtTYpwwGGAId3J9YfmbTR1rXFP+TYSxiIVefww8UdNQUkg0tIQMLGRLlFBH3LE
4Ey58oCBH46cKRlOpGVJ+LifgDM9M4Wwfl3e/CMXiBgQMRE1gRFUp71/rd9n4i/9
92e7jNugKX9UdzEUoabOF6t2DJmfx2nUKKU618HPP3SJg9ybl0Fecq85msVCJ11g
V4udYQw81OOUiRGi1FKsmGz5K3GhZ59eF77hKzkrjnCQ99G/HdFmqdvyKzv5/F1d
ArA8FxnYssBCsdA7g79HEFi908kbMw60GidrdfSRXIpT2nRTahD9IdPeMRMBfmLb
qjgNjSYsnsRqV3QDgD0aXSyaT9VD1EGEzlj4ZBcg7hzn6nNrUTiB+x/DB12RE/Vz
U1wJdjVt7jB7HlAAZRk6umAOKKMj+GhwsthilEmV8UcZCjN6dwT1/J1su6BU6Z9G
fw0eVnL5ny6idMLw0DHgWewuNVY54D6c+eTy1OvnWP4/Rz3ERi0Qnnuri4wA9Cfg
XwBi11hdM2gjsESAdszz31Ov+ZiMXAc2g0Y2jQah0vtu1tjVyipazv0MFrikY8ng
vzVOaik6T/KvXTmV4Myor3JfR54QqB39Deq4GVP00bjbQwZlg36qH6AO2+BeZsnm
cZpPXw/Gu/SeK0a6IBN5PJ2hUFaiPzWLnoObQiaLjDlvtdpeRu9OPZqNzeH08aYQ
ZwbiVUnVZzR7Od8r1Fs2aAJSysR5AXQmZhgCjPUbaH8QFoK0nN553en0EcN2nh1c
/phPd2Xw3vImPdptFPxJsgmCmqdFmwEC3R1aozc3A4X23vnWO4dJSlPQI0ppa0nM
x5b5+C7VATARLuA8j07vGMtvi0zsAl9Jt8cwHp6KgL5k/c1JB4RlN57X5BBBptIG
YUwdVE1FmQCW064SrhLCqyxK1GTxTgvUutRT3ve15oaztYMYrdxzM+tlHzEphq+C
rIZhK/KawVquMshTvP8xB1CIzqKnrjBPzSE166pmgWvLII0ACv7MNQ1kO9StsQaA
iJT1Z9r/ZAOKpgrBvc0fh4Qa3GJfiR2jo9JTFWYUiR7Fe+5kQ8nQl+/hw3lnO8gi
fLC2yWtJrn7ue+oHSsmtcciFcMupr3zcNifwUUCO0cM+0+CJolHE/zr5SZR4+nky
6hluAByrnRgfvMPDfzuuAWCrWJRipt+XAvWfESK3qm2aR7Ju9ARx0EStXfeVlt48
x1vL0ZQhEBH/XPPGWvZS1aNbQKu6wV90V0ZXukVXBIPzudaKT2YoOGpjIog0AHDh
d/WPK33LirPN7GuQKhDhKwxGuE7noIbX/RKhrfiMT85UhySBgXjWTsGUwky2ByCs
1CNJRJ+5jp/KyphwJtV8xIx1CEco40+IRPBXzWPthhb9QhI+/m7+gz8cIPfKCLG6
t9wmQB6DqEwTVvaHmOXIl6RVUVtOa+yEjI4352Gi4jscuhlI+mTmPC2mehXNaE+C
ktk5tRIIWublQhA9xHNTNhqqjpi1UU8YZCnroCh63X/J2A6FVd7dxUjoCUGhE4R+
Iv5Mib7uQ22j6oehCNqT0cHqrSKZTIWdNqRspyOOZ35UZiD42TNQrWdJ/EPTFxfD
J1uXaZ3iuJ58WTAzOv3wtayVkiwxDkXOKLvZ/VSR5UvzW/lR5sJWtfFueJHtR+tl
rVB/YzazEWAApKZ1mr9LrtStLuq89QgAoqnzzQIA3dkN1CtCKhrGi+OumDR+HPAG
gVSga425TmAiSk5r88f2Xiz21TmDwXnLrBxLw1h4S1jmgv+mfpihltxx2ufFefci
+TMKG5uIqqV/BKl6WM4rSzFAtyovNTIJd1gUaKOcwrZxlgCfacokgNLL3EuunHfg
kM0JWR30dtULr2ruRmFenU6kHh8P2rO88VXwWFpe7iYpAwNmT65KTjFg2aw9rFPN
EfBZPCfD5TGLQHcnaDhOMholEoZQAYZ5Eqpr0Q3D710lYzhVqzuE8iTPeDGefjl7
REDuv863AZZpxJR3+u1FkZfas/ZV6ioK/HCib60pYbkJ8ZwMF3ZReAtuK7K5K8yl
Vk9B32dycz+1ev16XTM3UFD+fzahbx0392BACiuq5tqcR+kSYhgYuYiPB544mbVP
6uFybZi9SzqD9zq8abjJgnf2iyjRvZ3KsQyvBEwrW7AEZmY+xENbryAH7f+xDCPQ
1oWp1L7s91iOatERyI9xFx0Kk9RSW6tc+N10SGuorMpRC4Vq+GVnl2t5eu2JP6bS
8w7VH38OKPS1TPzCzouoteTN3UTQDUGqiCEq/KZ7bL7jRDphNPH8v/mRwdvAlahS
Zo3GSXGK4NNVUovEZNAQXMwKY40xlL7vUHq3AgTJvRk+1p4XoiMXMJlX+9lWjcJg
Zlv1CK8udXqprVlWAFJOVCUrLwMTdlPqISQDcsIowlCJkFGisid6TuEe6zGDifNE
nqzVAsB3MFvyOyziEQLIthi3IG/rFte6kA2YZS93qDaGk8fsndH8aPEGNFdHbXU0
4Bkzif3RrM3DAomIKErhc6ZyMJgYSSj08VIbXFivD8fIRzQkRx2nMqAsF0YUY4EG
VaZY30TiS9D7DWXevuiIoWIs3QBl0BpClojqaw6kaZ+SbsfOdiWrRulFwXSbNCwg
aaIcXWI+abMivQaFb45yw/gzguhJYTjw9Qum5cZAXY1Co/db9TFXfSA0YLH3qiJA
TiqvnbJeLdN1PRpl/1shstbE07l/pE6mMNiOBXVmelB8PjHZrlZahX6VjHmc1yDZ
indT0f5hxRV80T3qzy/xxU/kVDwbMrwHuzGUQSVV884xn9119rkQVtws7zZ4ke+N
e5dR/fscUSYrh687UfeTv3ZUr4e/ZpyI2ukK+Fa6ca46tUAJUYioOCB0qbQ0EQOY
WhEnTVYTYTCjEKUu8PQcrX6XtA+Mb6ysOkvWQkBodsx9TFMTG82j2kQx+DPlarZG
K4kafKrFkukVXUpqdy5un1D79sXDurkTFTqGbtsHkqbhRuEsAtdZ0A/FAYapqiHR
ur/9Lk5+c5UOwKSVFo85c4dwI98zJbTwtmE4JIIFbFhfEmxJuAIloGf5f51TaQKT
MMN7Pl1+9I0bxbcCUg19+RVxUgPPCxFbMUi2hlRgVuPuz6WXa6RdHEvOVwcsN1xh
WLeGrstvow4ftDu6LmhaJkrCsza+naKUjFaRE36owXBEBIzpqca5CsByBKzbApGu
upLFHQTKHrEcnB5o1WwLqNubOeAAyqwmVSCmynW8jwZ54u0DDHeyvjEgsOxMSDXO
gFcDTh+ff3GaumEdg7F1e2SzVAnTf97dJ9EqPJC362N9ttX04KoD8vKSxPT35rN6
wq0qvflxnUa0QimsHRvHXkl6EDh/UmMvrpkku1khDgKwN7Nu+M/KlDCKz4W4kXce
aRWBN/UnFlRI8DG8SPOAZTvnZ5uAUeEgG4DgTbj1Mz/aZg9rMK7VTzBO1/nIpOnD
e0/JBG9gigaZDQtVfZR0jKDuMPd+ZY0lSsGwJs4UZxdl/3Xv3mhT/5Dtli1wIMdV
c/gfGRfWgKatzXGTMnKociS2JZG1fLIzZEjI4EBgqoHGr0+R/AD6Tp4QRzaFVNEB
xNp+tAlkoMh+8HX7FxnDEIw6cyDFMjCs6m5/NIhZPDqQpyEmyE2IOJN7jhb+CEWO
EFitieJB+ZcapmWpacVYQwiJcRhxGP2jS1P2YeLq07kyOy/0CPN9BozRgAYADtpf
SJ5VWbbAGkl2oflpuZZwvEclbKTXZ9y11s+qLXbdcxtaQwKWJKWgHMDM4hNPPUXU
xipYSaTuSUjpZWCwv2TrrnGl8tPLdDwQPvl/VIgkOqQWzUqMh1YXlH02Y565yqEa
ntpdaOK7wTh9pTDg2llAw88VICpXhTrJHOh/CEltjVn15+RLEhpiJyuRJtRip93y
IkLUGpzz+1/YUkw9V1MOXFE0ThUnVWMonI29Sek22dOzd2DBcoEXkSrrOWfVXGfy
AOTMlZF+58d07nUxDIkWEe4PLfYlxM3tjeehprJOGuX6gIllbWyjPGbWW5+OxFya
EJq5KRuIhLRgwCTQJT7ELb2U8x5ghRs2ugMX3EjeItRRHq+l78+DUre035HACeln
UGzsePSYKuccUeu2GZDQSChwcVg3+oKkHJq0H6cPIoBWygHusbvQ7WbXlsdVC5aJ
1Sb+8/d73lBQ2x0QqHq2djRS0FrsbrM/Tq6XxODCpQA7HP/U6v0j/xMtSx9tES68
wTv9lbsWB6DYNfjt5eo8bJLJL6JAGCzBudFwEJc+tq+ul/J7fiCol8VNLhh7s06x
gOlg82FrA2ivaXZNfYDazod0pAvhjZuOpxUn1m1KG6TmfI2QC2blRBxVDio0hNRt
ztEKvgYFhYuv5ZV+SUmw33imLcrTfhiEIs+8/A/9VWJB3JlGgDOYMlbd5A9vBo4+
NZ4YT8Z4jH1OcFO3tWVdpDDQHj+TvfH42o+4JughaPvhRMx4GX6cpszusg1ah9fY
wfZjyfAC/7PwiYbY2GXdcNEieAqNx7QOLm5wWJd6msTZIcx5KlpuH7g38Zc+iC/1
RNQuYYrTCoqAQx6bfLk3YASKDU/kiiht0gaolO7mn/2WJAZmtUmSf0eoInuuLLEd
MvzaebnQVSjIU3SZ3oHeisBHG5ss2NINvvkI5O9/5e4cgycFfFa9+WS5dYJqha32
5sBplNA0tYPJt5nmNVnWt8Yo7KmS9oMZk2Pz+crlXrsXRx0ky/ZrW7gELcIrENja
B1s7FtilnLMlNbr28DPH+mycPG9fdQ9vTjzrQyxu1eRs/Cw9yiBDJ7B7ac3/VPt4
5wgVy2+DqjiGI6GBssMhFoeZfN7RVUQLiSrI6aefJsV4q3gkW8ANP6FKvNkS6G9h
WmhwZT9hE/uY2OCMDE6ucZpaYEPq9RGvEjR/PFabOgwfYTSiLZebkbkWbrtOZu+e
Z6JKzqkqQ3h2/5HGIidrR1JTqkSR27ivm2Mg5kmrG4GLoLfL2fJPSA/uMZ9YCfFx
RWCmTLREM6aYorfEYRxXu2MTN8j8CW2Ei7QwtsPEzriikPImUsle0A8Gn3TVihst
cFBy4Fjgbx/0Kpaga0P1Tz2BeUzEqH4JvmqIlQB08CzUUpn3Mv/eP/g1SNoHbdgf
qJ3imYeRYAi1AONwYPtzv+Uo7RX+eRQtUN0zCOIqXFVEIgeVg5ENkoSS+aNoCw7v
OEr3wXlVcWX1Xx2x9qIlv8K+8vs+YREisNPEhDb/YHhdfOS6fMsgXE8XIbL1BKyk
NlkCbo2UWmxKROTxieNH7dFBRB2IjFIeksUuqPShp7DA3924X/hS1WcFCgMolaeN
GUa9s4/YDHWAxScBLIlComq89kzTdcNw4E732+7RebUphxPZ5t4qxfnx6fvZcGXh
xTyHeNdUigx6ftUe69ekMCn5P5K89ab1MS+zGWzgiLXQHEcNyiQjz7ZJTXm1ehS/
gHPzQ+QO9+qg4lqvzU/flLH7PjTEEQIxef8w0vIB5ise9wN6qf2pnQMAGwAo4Eai
PN673XVjyc4dc+Pvk2iJCQEVHVfvraFdE5/tB7hj4Vhb3E4eA9lZZDjlbzjSUIox
u9pP0kNQP95dLbGH4fOIsUT4ZdEroppOrAZw35GOZAs10DwFiTlL/U1itR/Ydysy
qE9CIAdE41+CMYjPeoPdL5dn2oZCPnBE/cxY653vgIFbzQy0GYRieYgc8tRviE6z
mbQ205lINobiEQLbJmUcb7Y5HOvzBTfl9SxPE6eOCnY/fvjbTf3SjWP+s+Lq0CV+
El0wtZwiyXVY8Bqq7o8HFZIaMe2H9CRXDWPXOjQ/5GmWGqDqN0DMKDkVGzW8BrLy
Y3luq51POcsFjgmweXHgy/ohHVYXkpttiwyeL/6mJeLIEqNcVex6SRR+5474bFZN
BU/erhwOpjy2/0tj/n+o10yGm/xCFbw7vt2jwrQp+CYkTt34/9sxnR50OWOqVh+H
N6q5EpxNq+xNxV6JsoetkgHIxJdMgOL2yEnr1gbGp0w4EzY/draTaUGtW2CpN1iN
keZUwij96AEtsI1CWgFkKGlAQ1a4IzUOl5nJtvDGvjDiyXVkuAQTOrQl6uIsfAtd
tYKgN53AMfyfCZkmzHO5dS1+UTTe4DpZLGtRE3MlmXkySMx24MoZQgCITHpkMT8c
N9zV0O7tKlkGe0tM9hZNGAAe34pRfnfjbM4E6WKW67VU7Rg01RiUWyvZ/RqZXAoC
Ewj9vo2reygW9ebxE/NTJP6yhRjJ4btbxwa56p5NEX/XOE7cmgdKNaFc6OfJUhBB
/2BsUSxR5tzIyaBk2gp+mzCueG6AlNj/BIw8L2cYjPsVnBETD/CE0FXpewiUuafJ
wjxNVkiTKwV2j4b3cWvc9iPYjFYVZfBTOdgTbvdYiFtVSZQO21rql+4hT5pMPc3i
nx1L4SCnJsmkQZ7I81Bd9sPwwwE0IM1DEuz+8z4b90FQUvvg8+yS4pnRqNccfzJC
yWj9PTINWR1/Uo/kqULDY2Qdt1BWHWe8cqcYtybYojhU8CP+lbgPgG1tiN78rbvH
DE+lDnj+4UlDbrutFX8/7EOnlLtre3vFbnrxCerpyb6j0Zrtls5fIlVazPSQbSYx
AvfS20Tfxr1cA/1rJGOWvUG6kaUjiXqbq/ecYSw85fHfLXl0NaJ2n/oWKDUwUrhs
0qXalwz4LED+50Q+VqamCHKjKUqTXJ160rFxKfLCHgJHnc3wWsBHq5ULZdFoWrlS
KVJdXbry0NN96BO1QKCyuj39SB7Scko3Z5WImwJKaOggOcGxVMOVC9q/psVtZCrl
iwJgkJo3pJ0hcAtIZH8uXFVRZ6gRtuI6xIp/uscCN9ANPCCHKmGWpVK1ORn/W9ld
l5yIDSDipAMYe4Ez3kL9NMs2tM+iZhtbLxJO4H0btGduTB/JnQ9NPgF7xBkQXhRA
K5KqKmgg/b3k+/WW//XXg46J3IDo+4zwFi2l9132MszP2X5YAS+zUQ6RXmr9/IsR
zGEnAQ+sUD4mj74S//TI+leQhdJOOZec3J8cTicX3G3z0tAVuP8OcKb7VNnvIj1e
D6JMxNOWioEPTKlW3HZqEH0wguV4fq654/IJFdOroACWGzT6dqQ4Dmuk96aapM1C
ZeFSxeDZAFeGvhdKMFnS8Rrd+24eNwooZj1LEmlyTAp1OdbhSOY1Q6sD6emUSOAM
xuoRm44VVGhzvqFg92ZZIBIKDnmtRn7YEgzskNrlh2E9WklYVU1IMyjdQV2qu7DS
6lhrABnSA7BVVtAeD/useyLgKaWrm01HmInQMxZE6/O4QEZyBdK8gN/WxX8XtqVD
KL7AiJQCbAdUIGptxSFUDvBGb15ccYm8Z4R92PSfWcylxwIGrtFkdKMTe74HUJb8
w3YNUWox3s1SUr/NIOXVRLRjrYKR2tJ2lrOD1dhNwgYev6OJSD4trkbJgxG5Pne8
5O32vusGcSUakJ6fOrGPqMb+4wCcEp58eT1xbM5JTX9reX634CCe1ld6l7KzEFY8
DWKCZ8SrJS738/mIg9ulicUEug8eq7CA6datv7IJ5zf6UaA6gMUmSzNhkbGD4oqK
Oycoy28igFsd3V9WvpbMl0PEyT2ylaOn1y3xGf8qBtQDQursPa0FE6X5UumUxE6V
9jd5Uvni6hrTDvhs+MYeXKhqItFw2wSpKwIS9YbcxC5Rpb0P9QZdwkaeDQtSoaPH
wDZFc3dJ9YNcBTDLSOMw0R/UoTOQmaseEZ0S31V50QcrZ+N5WneS8k6HtpXeuaGA
4vKTwcVmkVZkQbXh73KFiR2gLcs1ETIxS8C1sMT2oALm4YA9kdOBtQL6/p8zB+ZQ
JV0j0xjP3aixonaXQwLqjFeXBOr/7cCAFBphk5tztLCDAXsKqas07jPoUyyrXobN
epQYLgThh1cPvbRxEsth/U4aKAcZVnFfmJGQSD2VWa9d0QXU7t0LB4FlaqFpx7Cl
ukTsv6WoXZUl72IXM7N2rgSJwo2xrlo4W9VxgMhfKSXLm1m18WWVLRvLCob/jS0z
B9L+cD9gfcW7AL1WuU0uxvRwB9pDXNAXRQaIn9wZWV3qqVY3gXaJ7kYKoBxDBRBs
lm7tIb21peMNZSqoRU+H4IkMfD1KAj9QcTbtsJN/euhJzALb7CKEjUP5mmUzVoKe
OrZffOIkDNm9j+BpB+SSuZS3H+taTcBasUngmhTfcrzjtg7xhSEJNITiOApyxqy5
KqHg6kWtMQtjxbENOLX64aO5mQcO64vOlo066weLk2o+wE7ZEctb0DLIxfAjb6/s
iZ/suIwomEwS3/cw3vSdgHS+YAuRAJi3C8NaH6zC7/j6B9WGNjGLBQYEGGbEtg1x
HJrs5fe+wWjMpvVY3yLr7TOGXqNmbhGXgOVDyhgq+GkMCJsg3gJ8utl3mhQHfHQN
Zejgj7Vdq0Nvhp2a4SSq9o3mdZ9UoHrBcO3kS8nUVXh/Sp6sUQvYHe94RpShTt/g
5+jpeF1d+g6WLcLTcWmuvB1PIodrz8BhK3C95EJUHiSEUYnBGJPNpomVynAzH400
uFK8DDF6417J3T/KJEPlbX9GxGrHpdYc5lG66alccvU9Whaa5lLhvf3CHladiF3U
IVERe5i0B51ClgRYB81B7RcOJLxjSKjxOHEBDOJ09WwRNI6DToEAzs2WiyiZTg/H
cJvgS8pkTxi3vhKwO7kqNB6ePiRQshdDsvq0G++PwkZkEY8GQWxp07KDNb3h8tha
yW+tRKUv6ctjWaJmKVZA8ZzShHKa6a7LN7hOFa1n65AL7Ehw/djV0CgtnNruFFPU
xsApcNybK1xDbsWwQwXxbZCHvj3Vew/Eild43DSksnmSXu+7j3xG+ycbIOVcWYz/
uhcelR5U268D9pxOJWaQo2lQBC7BDyHEyv4cp6unFMzF2q8X/KlNd+sVwMYgVac6
bhwsjJ6M7CwREYx/1RIcyAm3odflrJfnCHEKIHPf/GK9v+1xtDJ7QUqMatDicplN
qAQhHsW64MuD0G2AtmHgdgJ9koPz9XJIt6u5CRSYUPGxpnOzJaD2T19Z/3dMb77Z
9NUaMyZouzVyBmgGESLLcbTRFq0bLsOX48QSBBL6Q+8wenPouKaUr4CqPbBOfuvc
+etadCjmx3o+R/DbA3aUxuhIpOJTh8MerySbYcEkJEmKPCaJyvPFq7PI5lmZbd7J
t/6dckJFrgB2BRL5dx8H4RXg9gcdspHeJmw3U4GUJ9ruN5ekgAPucCb+2DEhmLmY
GzZtd8U9H1y/iqvBfkOCy0+7Qthyjxgy2TcjkqR2prJJZqW/SqNR37vI7RHGQyN3
jVbrfs2d3mSzjeMtxGNPs6b68dJdxrIvbKwTsLUZcnsL/dbizmm0jqQJT0vsy4cz
pA5wkrGbEVqIgXGiWQ03D/D0men273Wu/OsUHso/3l/u6lB5uIhi5ygTipml3cGa
pkFquARBf30u3wvO1/xzlg0V2Cu1KOGzC+sBIZGLMrMZ7+QlqJqi7cGEji9AqwU5
FctoBDzTHFfH4/LrcG/fjrT3xrNGFM49qHL6L3Vqorna6Ib4SRI4thJdN6Uu0C09
KNs7g2GJNqfpzBXLFweLEhwJvnLt3eb6owCkPNNCHyzlxBQ0AtHCtwjHDdp8Hcz9
Ha0vxazuIhGzXEvmbs4nYjE0tM85ZTXVzUIIx/hbtpxKpszDPTB3Sqiy+9Dukvre
0gzSciXlF777c0dqMSK/a/E/xm+AwRvnx1E1bl+ZmJgFYGXQs50w1s9mXcbxhrrI
CfqxVEAPc6sNS07h/IsouK+TfTUqGwsnvDGY9wBHfX5N2iyWo09wd47w0Y87NtYa
1+CxAtNu9MdkOF75tVpYppE0MjH1bbgn25PltfSiTcNIGO/nh6IqCgmmUrbSJYzS
YatwU8XYROtMpTzxkK7bxvbhDlGHRxzY13kkL8WQ9oDrMZr5wAJtxoAnVBiPu7lU
Y6a8BkAdCdvJTjRKW78K8p9cDK3K9sPnuADGWcM0iwO/mxw9gekViRUfkWo3XOTI
DIEbLQBsUgAkVcffxzo2HwVpCJ4CjlXEMxoTbIKVzOKtgjQgFbDFyhnh1RkDJ0oH
IzZNn/WrokwENKyPrJvC6jNLuYTwAIgYt5g8hJ++Spm/tZwa/OgEnNRySZ1HeUki
l/u92Iq7ZkE6Iql3mrJ4p8eDSrUfLt/1ElIq7HvSyjxaCNevznAfBAohrLIjRRlw
Vzuidq7hgJsIPIYXDNgY/Qa+Qe9ZRKDhrHneS5NZE4lm6bzoplUQ6n3aVZy/By/o
J6lqmext2dAjeKscqT0MxddE18EcKIzVf9g07Hp2lrcsY7ADMN3GwO5axbNsHsFV
V/Is1i4p0PA/dZwpTniJpeu2+9GW/afdMsdEuDkuZ2KaFbdh9o6B/9M0aiQtbBYR
zpCGaT/Da4V5bAGhn2p6GOIkUtgC1g/IiwbeToxKTQi3j0YRAj9pCTLM7OtmB+jM
V6h+cBPxqfxaRCQEh68wxp5/mGX6ilYZMFcCNd6AkumlhYPr9dUkj9yHgUCXy3Fu
56kBvL1YK25esOl3FLwKlJ2SggCZxjuIaUPH0hE6uLf71mhzcYwb9OTy04R2YPR4
b7Nro27KWsL+IfkRLsCH+Mh9FrORc8X1Lbj8t9FZ/RKsXvCttiesiuE91oAOgLUi
ARFPVlJbYRiUdXRwvG2CeUh+IrjYVR9RNwK8WAwk/DpyjESHGGIohmXbjnC5ab+D
3drVNv/Uav9NsIS1ysphrHjmurbOeo1VYW1eivB+Mg8xgFs0og/74EBjkaYmWpCP
rqOVH/3XYZcDPVhRxmIFb9eYZ4xoItXPN3AcqBcxAqQQRxJUiCrfOEJSlGxTk+A/
p2fRk/FeGMcZ5y0UwpILM/NdiCoKMryHvNEKN962RCZ00VQJGYtcuPBkIoyU7kXm
xIR0WqBH5WpEfcEBezAfz4GpCH0UvWKMM4B4EHKTgwdi2TPrHQZtPVAQ5oUUJu+m
f+mD9sqCE50A10SZfoPrU935dQw742W8BeqEAWkf+TmbnMEaSYbQ+/r3PCOVroRZ
xNwXqnPnzL4diY8b5jNhDBnkpL0LvVRGvy1FAQVBmmzX362cwjuYFnqypBmuag6s
p2+c96p9MiXwEP2+jMsDBp/VzKUP+yJ/Ex/fNRRWvcFOOG9la6O1nhbBNujvvlZf
OHrE5BmDM9r05Ba9G9gTM61dYWQnbBDTW8+yzLp64NGTvb29tzCG7BGdV4FG0LeJ
95wbiq9IbMIdcgZC9yIddHYkSmU+AgujUONiMK4TCsRRYzcW4FNgJrNdwbXdcm/g
hoHL5/va4FcCKaya/SXRoYA2DD0Hea5kZvVqjGnID0QiY9GBMqyFsT68/eRf6RJy
9HC8L3phVIRFUdGIVfq75LiIJ71DyT51tmX3Rs6lxMeOD/Z3/2vCASDKwYj6BQU8
iaVW0ym3m/PISZGRCiIN7y1yFOw7y0TNZl2Zw+gJDsQzeyzNTmAM+uq8MCdJOUCC
3GAeoLp0FWuUWRR6An29FkVER6o84Rimnw9UazLVNITqumiKfsU02qLU84fYxt5K
SNVaXscYKZu8z+Pk2z/zm1EKMyAAUg3M95759g3koGwLWJVOuEsQO9tWQCmWozFP
vH8qnluyBW2jCwVABx2LBKaPZxn+wJZRlX0srvB94D5Cto7lVWA7cPKoj3fB8U4P
70z8vbUBGpvEj7REfjDOeBVeDTBRfmA3FlTHg+2+2XL08uWdckZQ22Tgodknkoel
a+bCSevL2+aPEMUwnwoNYFwGwv7ESdxV93nHhAPQdlNz2+yn2XIo342XuBhbJAIv
L6LM7F08x/9UoEfVeCSkN/fbd3ItU2lk14i0co9Koa3n4dwowq7vQAE85PeFBvaM
8dnW1EQjZwMvW6vGTA07LQfLxM2OoSyfLXwkWUH4SKDI2SGWALT0WFWU7znCeDpx
zrhrRHCDtYYFlhj+w3cULeyEw8gQ8UsZswM4vMiv3KAJBleYq6v3sXytx88NnYZQ
s4IddAiugf9zwfPDd9c6/6jl4TAE9ektxY2Qra1KQEMlnpfODNFsOMWlrQ1CEtNb
I8uYK07QEOprRxxiSODoeNP5YNseRHCQ7L6Vj8x0tvF6j0HfpyEs3n71I2vA2/VF
Qoo0OtfHGe8FSu2bhxMUrcYY7Ub3Np6tkMebvWvtTuEKcC2CQClQWTgIpMM7G9g/
zpnTSBLdE0Kmxd1114A/6MKi2DnwEbnSst+CzHBtcyd6B5G6J+VEUZyacKTI0dZV
6IcdOL95Yk1/7CDeSYvLHBt8FN4y7aAjL4+BPIhGpU8sOVbVdTXqdBst26SE/b+w
ZzHD13ktv9Bhj5Pxv9DX8i/+UscciS6hNSD9Z0+Y/Ftiy9mXAgmgo9/P+djpO15A
Jq6Fz1wE+8vPST6Gm/e+oukbUTfKwTuAKdRSHG1AH8JEKV2gspDSBNQ5DX9nL0kq
dd4CC/bJfQf3x724zcReluwQQZvU/KuZVZoJtndsCmNBVuJS3UaQ37NKG595KPkm
vRQFqWFDzqOJC9Xc3r5HYPaw2YvVJ8yKL4a3tux6hbYiwESRiGT+iHJQr0Ll7b+k
1twi2mQpAmlj1OThaFoCHJhqyf6n5ieVz269YZQ6duiv3PL+HyEwIoLIWX9SoFJK
0XoYQLgjjzUk2z3sp7K6w1At81L7qfWUPvv4fO14W//VecrtsmesNyTDwhfQm7uA
+e7SUyGhd/n+oYarz5MTQ41P/CP7uAVXPM/eGGfUtuZylm9p5zFMLkPdO4TPLVcZ
9auZMisVPQLE0tfx2+TiBr4DnbZmfDiywmIQ/lk+qc4NOEbLZkxntve9pbrSxNKW
wA9eVVBHcOvq8ysXfUklRvNq1/v8pD0AcFGL0M4mrK7qG0udloUQvwqS9lEQ4Fcc
xu2F6QnkgAB5HLcf8WBWqqpZvZWhsCj1q5mcZgbtq3aEYAq+OwSi2i/UMdpObCkm
0YfmuSzDXEn/l7XgbhJPLQnPYjrbinnmF3AYkPVug2XOBzzUnaTSXwfymVHghYc+
LQPaG7v7qt7cQLKo66abPPVSti2lH3sDvfKuPPs8pJbywdEgykN32LmO3XMUlXOg
sLGMqHw6NIjZo//pn/vTtT8u66paxD43R3woTELJjDZua6slD1Q7UyQ72Cai0i20
WUAYSoZB/NX65zOywHxvA6lUB0dxB5TmMN9LrzG/5RxhiDDLvQBdVRhF+9eUmmfx
nZ72grRcUFm+oMjClfpuOZAJe7p7XBF4RwwOcxhEGglsVH5kWSg3KZVZiJuh+saU
6Vp1Owh8zkSY2ZigLw4euRQj4InW89yZOe9mB3zaifd9guZ35lxyoo7dSGsTK+jx
CrULOHiX6XpSqN7Qz2iWtpaMEKtk3fkGJIgRVSKcsZlMyP3adUf/bWavPghi7p2A
aA4NbOF3UtcO9Rh6mrKiLjA/eQZmk69G8HFq5mHmcuaFQlnNg6EZadqiyq61vzUR
msnOselqph/2M8St27xYgELicDTIHsDlrDcxMUbVMuxu5DVtI7RYOqrvl25u4fH6
M36LBBVGj+h+hjP/xfvNXNG3YTXT7MsbnlF7cYStDbPnbhfr3ld8myFBSauwEvOC
/CFdE8q0h0GjNdHf9v8PlEGoDTybUlf03QC73eqNEB1lcv4Pai/z3SWcxIm5Uje+
Z2w9voMPJlWB5J81J4dw5TgKg0f7n+lgOAdejH8GHFxxy9dcK/qP6Zf0Dw3hPOz4
aYYDXYoSz5qyNRbUa5aF3YigqpW7BghyFC3FvDF/9o7vg5xHMj66LFFbYygwzYld
ArHpFClWuzl9pXQ/nigUlcSsNVrDj013s3f5Oi+EOjvGmAjtOyERZ9AZ18VtKcnz
4mSU4h8i2mIpgUa9S9c3ffvLip5PebUeiCeHohm5qwGxcwoTfNFe4DsvCHLU51aQ
789+jly2cd7ef8MSoOLBYRidzmulmrsXVe1zrMk2svvREOpuxbKi3vMf1p0liIw2
U2pElwaK6vP85o9UosNO8U9B34jy04OPllTI3aJH73f2uh+ul/x1Xv30kSiuw7Ou
5cm5YntAjGdfk/ucv3TcVK1C2tO/CeNbpatCRy0RssRNa0u8MUCprLkA1t3E4gVJ
ng1zpHbXI1KOVCXGcI05lWQgmHPr4qZIeJvU905Mq0Ms73xuxLJ+pzou2XH4TvSm
zq+J6nvg+JGJwbfg1G8fWPhTLyE7QqvnUmiyzuex1T+rp67+Ejh7BAc4uOsJQkjK
B9KuRUwpzT1ks+Tb+DQSMz1+EiInxcHsqqTK29ult630xBJRQYh5nlWEWiNHpjP1
HZLydilbksU5MDrWt4AeVREsNxBMm2tyrQakZsS6qtdUY+9g9JzMxsnrRXwXoCKz
Y8nFD0KOVYzO1N4DIiZKECm0TQq9APjpntCk9WS+/QKZugp8WMBa3rafryqKivsd
IShKYhK+2OvFzzD9wvqXdj1B08OOzee8Z/BfUCEx6YcpX/ioV890sRyGE5F5hmP+
iBwqIbqly4uc652O4som2s+LlHa0dQk0CZRp5BD4PRKxzf+AHGtogYMl3o/7RZxM
gr4SZnuvw9traRAEDjj9/TQafBuD9GaArgiqeCfdxU9XbIs0BMux5nr4Wt0StEyr
+aLOs2YXOqs4CCyoo4bGRY4wEO+WxboGtv40KO1WfC/O/29685uNjx8hIQbOZrPg
qVPM6nzgW/JIuxXT+2lPUTMgPKtgPsvL1wzsXcxNCMz8ljk/ZvswSKXc5GzJZu0o
xnn7pXkKUoHZ9j1trqLsiD1WUkVsR+u5sNs9rwVLtUnS6qHg7MDPBpyV2Lqeaiwo
+IGLJ/OzxDYZPfjUGCWP0f0FLxkoRMG+hzFGzzu9ppsqg4JEnbWu+lIIBblAV4QV
PqStDZrYXg50E9KjsiXugnczRgDpDCdQ3xfSI5bQSB9I5Xbq7eHEnXmn0xtgvljO
RlaEuunc3Ry8+Aprn4Y6cOO3E8JgUuqPAthjkMnsIen8/TzwjDqDAz9ea1fX0zf4
XYqqODZccz/BqC1xV5cA3x9tG3cOPk8W0ohb5jPF+5IW0nJ1bqI4YxbRXahmkiwk
E2jS/RUHgLv4a0jDq5037jD080/QrFpFH2kSH9WfC+Py83Az/RXl1tlmEjSSNKcO
R7I6lpSVQwY+SvkHDcmgcfAGJJq230/sx1cu+/YZq05jv/SZ00VcmQ9GZCndGUmW
ulK9Ys1Jo1Uxy4YpfVKs0jtvSqApezCftLcqtJfK0pBv8zCSWG0W3yktruT8D2jT
libkMxjg5yEiN1OcL/ZAlCtROcSosQmXRcOzcywBZ1nKWLOHN20CGU8Jt00/8e1S
3p79cQ2jHsTfXLeUl8hJB682BYkre6hDQW8zYVX3G0hZ5XGfkC1LP76Ok2GuPwwI
Q1L/V5+tRUJ91RepRdrbSXyZod9fB+mCX1tpzk5tytqCCrzLUzlBgeZixveHNZVb
kmOQdKi7pcaK8hvZ7GuBNehkK9Wet2h+qHszqmL2Bwdt+SoZ3JwdInYuQD6RD/zJ
2ds9ijetKxcrr/UYs6FIkOGVjDqVePBlYKhPnKpYhsylx0AfthX7lXAmOjIdHOfC
3NBJ7PSKrC9EN+xV4nOKbUG0WoYVrUMBIhA5i44cc4H7chfiw+yzAYTT0D/JEMFr
8BGPowucP6/Bs/ITiCBdVZsT+xBJWLh5qCuifw8IeLCMntD4fZUc2wKZ2J5p650D
EH+EjTvTBdn+7IqoqIEQ+xlUiSLYR18RsQ0pMDAI2loOVKzbppFUlz5JBIqLBLqJ
EDz4Cx6WR0Zv66tCE2Qj+eg0iLfCOss/NVQUAOhXClR0ghA/jrHOu96mV+IfAJRb
5Nwp3tV+00AMnigzjsxFD1dREPJwquVCVZR/REkVFmZzp5owgqdTIPG2LU3A6r4O
mqURTJBEcqjcnz3M738uPefxBu2miOrcY05kNS7dxgmU6g3HyQVJTMpMVggScGg8
gdkGoc5qAzsq+HRRfHL81s2ME280ZS443yO5PEZ4mBtNW6baO/z1h12BYTx++C25
INMKDZRA22q9OQv8euH+CdcjulEwbNVCr6rJeg2qSVbvuDmXRgDl2P0hdDm3HA43
2kwy4K/YqQ6HyGXb0TOwBkTTAm7ef+3Uyf2+6tjZXp9FWd8oKcXSc3k+TpeAQoBv
9JiRUOBS1aoYFNxgoXYSW+aWRzP6IhsO5wDpXk6Air16/hfAAD7MAvvDX2TrymNL
OSRhGiaWrypwgd7Jw43wvj7AvDleYb4vlFQiDbgHjdNBhtCc3zut9wiM8i3JQj2E
SVOmg0bs60p7Mj3zIPIRYVILqFe47S7yjYahXE0r4/0rcJCgxquCYHpfkUPPJQ5m
smj5OIiLo0X0iic1jaEjmP/UvLlRLxV8vsAFM5JRO20h5hicTNBPdJiE7k9S07Ei
/1xGW6G/bhSk2K4ckPRXj/PagLlWNkmAp0gTHDCHgWeOaEyfOSfmq3FKJ8yILfNA
+noqc5Hz3ELgdu2X9CwJObDPUHmZHCGdROdJPnKNEcr+KCAC1Gr9LWCNObXmlaGq
QcEyxEfK4BFnmgZex08OseuyKPgkjYCiq88iQsV7FdNfdOxkiDppXa3eNxNFwbgP
u9PP+smRJBbDZkl4Ol3aQGoE6XRKMlp8aBsyiJOSEWf9uCMi5F5YBjtisCEqasnf
zX38KW6HuzxcTdFoM6l4Bb5Zjh34ZBUaGLQIO7dfP3bgQCYUPo6XRreMe1BE4jtB
wNGt28or/uAiaKdU8WjNjA+MwfnUAGmWh6TSSsQknSE2QUIHQGnWAsfy4MwGr3Pr
y/kJlXVtJFxncS2nkpKqjIYiWtWPncGWLB0nQSZWgbybdMj1Qdr444ng9FkNpUlN
nbr97XRPp0OO/7SgNXS2GNCOVpWTvcY+arDEtM2EURKqhcd5XGMoT5ZSlfE9zwl3
PkuCae9hwvyrWuzzM7uwqJwoQ1nVhLMwKPG+Lmq2T5LbLHmwRYXWpicov1t5nl47
zexyizsxzxCJRIZt/T/DQ8A1ohRg9ms0Rzy4E0k9YnllYCeKiZXWV0jZwbcQR5V1
nPlmxiCrgLHpY98WSLMQkDrts2h+X8igIpwTYu4bXw5jzP1eEjCzfg4gJRVE5Uxu
UmeTM46VEloBMglbAW2UqhHYl4Y8I7F6kdbhYomVYzr0oEMBg/uOuA9K7nZQNHzl
ft/BvuMCVYzKbjlKTj7eMwaFXV1x+QmV0MrjljVPdTKLYw//8BwK7Wvui7nm0yIm
mKG0+DDfCU1MbViqz9A+UeccnFhZ2jTRazVmDcC0xknrXJSaZyoaG1YRA2a6Aauf
1QXtpXcYkqLl0H6JoH4oJJBzOBWv31bKSjZWyxe5JtJyCUm8NBbwykjwE7OzyVXF
ePmuT44M42alDhcbMs0jEMmfy1CUauflpRHDdLSf8N/jfRCDqtD88YbpwKJyB6Nv
ufaXrmHKtbwd2f/O+RutaDgx9+kwEK3tweo3npzTsNoWj5IKC8APS+OrGMya/TiX
MTM+AWPwyEyCopk+rE12pRTeOz7IVG1cm3uIvboIFbNS2R67Q1fqFh2Xx+qsMUiF
VG7cMCMR7XtGjfVwsXBMRblfVUk/y3+L+aGwCxuKzU3BS+VqdPH96USXz94Kzyoo
mLbNOYajOkySXYBp4duVEsgnOR51+NMqBpxDMjd2e2loLUWWYjnDQIhvSb+0J/y9
1Y/aitWo8L4sOyVUKNqzK9dBSadHwHKUCQKZZP8oJ1edxD/hSPHaMUgogTIhQ9ub
LloW+XBeWXroulW1rSOfdNyu/S0Bk9iLFBcQcWWb4+E2bZrgCndhFvDjFCSodM1W
mw/3lis7gDGihRkn0N3EVwcx6a5943WofR611lIj7cKr7j7mVpQ1qdzgela0wFrw
S0u+8xtEP2d4lsxXN6ZyXyGTHjaDmadaTriAPuWSThhFnqeBY4WDcbJ5RqGwZFDr
o3RjaOLLfdyxnDY/18mGCRUsN0H62zEmf9nASsNCBGqZw7bJtIzbv/8tTqlpP5WL
yziXapiRvXh+cgVB1QSHZw5CZB7Dl5JpjqKgSPBi2/w+VxbDcYomf7FLU+y90QnL
BhgBdgvf4uGwvp1C1tuuaxWvftQoJ2Yc9/MK2d3bgyNWjldn/iyPUGt3Qm4uW8zY
MosaQsRYr2WDaTHux7YVeA1ZsTTzfD6okCAFdwLsKgikZvQxFSb0q89bkS9N5RaL
EE1Kp6LV9xWMSelzUBg+kOmJemjd7X/5doWQErYhRC54jMprx1fIgf9BjDqENyJX
57deWzA7VELate11bvohrhQVXguohoarSrvAnxcyZVxGLlStip1biKgpgmOvUrPv
8xvAJxsGxXyAEaNglTxPNbAgp4Mhf7dV5rge8RxofOHAbIfLhY08W+4fnavTLa+L
IwROq0Xtavhbgy+SdFqfcEC42FO6z8kzFMjHeaBFQ+zQAdrRePIdfmPOcGrmDfja
pWVu5ny5K7i4KRT8POGCQLFiZLMSg73udvvBmHp0yHyTafrHWa8pnSJUwXZpfkgg
6mdWIfM5QuGxcb6bBu9S+Z7Y/GXijCBVZhwJxl7oPBSstbBVefQZ0Cce5TScZ/hK
buJI0tIHhBf/uD4xSRlLIeOJ7+/WHd3IXTjWVRd/jxSG/p2MbDrVabz2h3xapys2
Eqkr9Gc/aG7GU276TG+qAkKaH4iTw7a3F+7lt8qCZempI/seuNDWKwLIWJeoMCYz
ZL3PZkGYnMOVCPYj/Qxb8VH8U5GaR81/r8AIH7NTr54csTwIRNRW76+9oQGt210u
fNgXTCfIFZv7a5MglqOFYqkKm85A6WudeiSJ1qN7BLNVua4KabIAyLYgupDK1T2A
gxyjlQUZhQCyW22Cs0RbOz31qhGFjbFfHUUrwpVwTRtIMPavH/PEFCBXeENN2wkP
ES1UBzOShtuboVxWsDHJDngHB52JDwcYfwHa5pwzQkkzVN/h9ljo0GqOP3MLb6Bg
zQDRKwxsyynsdcUnXWTfjYVk9K8f/tj0OYNEkjQTIO63yKuptuPgrj/8witXNLmu
F+C7WnX3x/FuFyssNluCAt2++2EsyMjhyT+UtGkUPU13C43WEkRYBRpFEZTmRVJG
DSuQUezT3w1bE90cxdj5YXKfyeXLnganSfYVSczgfibizRM6i+DuwnUZR0p733IA
gNGdlYRmAJS6CXRn7aHsuH0yrwH4rNbJQN8/byC6fzn12hRYSlE8MMEhZ/eRlRia
IcVtVqACVH7zl9sH0cbI9VyMIkBoiJcVg9JcEuCPwFRoa/wUMTZ5FN+9PfPXtdPL
AajPsMA09wFjzVXqDJcT22E+9DfjGTg/iQ3J+O5B6tukSKTwLz2pogS9v7qgcfVJ
nF+CK9ZQK26KQ5MykEBM0VqxjgpUH8B6gBBpPQW7TRV5kj/xzY2El9VzN5EMgwBN
DaYJ3rfuO2czfcuBQ9shoAFevx6fCQYHG7tZJ+ZZjcHqQPfwYaaiOVHiaYTfXmmh
J4u2cXvQATdPqMTH8nGxKDFYOBTpKFsdzjuWpaiQ9xvyBWCEocLXlqqukXnK2d5p
NufDyNijLGoje25ng1JeSuskNBlFA1D7dHZ82bRj8u7lzxUGnJCiRsUyZx4TC9zQ
UR38BsfppyH7uZOsUncw+WqQPWV4Fd+82UqwmvxUVUpzKJG3yopXrqYAO42aY+XE
3HFXj6W9Ur9CM8Y/SDqPBLyg9i6YpJ++XqffMkBmWTErNSVOnTmRY7LRx48Xs+iu
vKFSMl8tt2lVnoyf5PJdgb8khA8hRNR8wq5+dWo4vBjEAIY94tsxtNYk6mVIg9EQ
4T3+D6Sa9zwnqKMJX7YvPjY9qYwoSDYaxKg5XXRskVgPPEppz/ykFue7e+nm9ien
PttS+o62zGL1vTp2+dNrMR0aGHlQZ1sbmdogoIGUDyfS+ErtbuXO2yAYWwFRUIIB
zXiB9zacBw/8ypraC5XPhI43rCeIpdvP0LKQ50aoRpuR4Mq3f4VrMAosj2FfZObT
KICm9u2rVpO6t2f0QLBrVte+s/LEwtFJa8hKgr3k/Cic3pktg9PntUuLR6+AtF0z
L9LCToFe56XTptJWD3qgCxki6OtjNlNcBWf+HRJ+ixOHloh5UbpoyxPmHff7LuQl
1U93q3wCUcN3UooFfs7PsFI+SY6IM7y6EDh7mMFFD3iNRowwaNx+lfFAduogkm02
kG2J8yFMYwFwP7kJ4yyDoNR0RvNRpIbF41eUirmhojELRJdIXlzmDgx+zcoKJXqZ
/Z3aMTDka9c+qDFYsX0bHopwKBCaysdJN2ET44gZn5z/thkJn8duaZKh+sfDqX+S
ix01UEAhP2r4LEtg3MgvuYzpsoFLUmzW4VAsXIdGh7YqHuEzTYE4Ueg02FyUzHIe
4hUupB/OsaMvf96KVY5eKWSUYj7F+OHhQdwAD3m9pKK5RnB318kp9RIpRIPlZ07o
3zjttwZrLug4JRBM1hG9lCVhP2NUtvJPpAtHT+nHCztt++HgZwX3w/ZKqQdZcS7g
znMqFngjCaW1eC55a6nQ6swbmNC5TNeJvLH0SesksuvaqClcNaDYz+oEjZNUEWwB
QkCBahCIFJJNhoGVVo9ozAtWXbXfwE8bbuIrxZ4t/Q8ITWh57zrJeqxwkBu80tWK
D+Ft5IfU/Ocg4ALrUof/y06srYM2nIFeweYBqpck6qmHhsUoXhQFD5+rJAWsykV1
Pv8hjUOz/qHmBMZKresMTHsYXITD50nvE/nkGRWyASsZTNaTdqOCmp/Bn16gIcuy
u6ecNwGi5GViW9j1DB3kPTMaKBfhMQuFgtZ6tKX+fgCL+yn4vYzq9ATOUnlhgczj
iizcpIgp2iESkeZBosJhEmw5XztBz2Hs22cOhEo8ELCGFUmfZ6cZSHZ1VRpm4/Ox
us/uS2X2g/CbwA1xRRFsqvyFfvRvGzN2POpPdxTxw0iNeReCcgGTZEYOtbisHvs8
lISvqvZjY/ZYtsdul5sAJlaZk/61dJ2Gd0zQqR2GvuXKCv+Q8H0QeQZe1GAAUHuo
l0VQLhd5TR3nLupnNBxpxnkaLiF4RWrop4HzBFDWP7Jk5++zbbBI8qiTW9vojpru
xg5vG6B/1ZrYMZJ8gQVTl0ebL3tlvZJ6ZNpxSrzcoKJ9PWaVOxtI5rVgpjE1TlhN
n+WlKWC2o183ynWV6DIZAGgy6c+3j+nISbTqT9YSg4fJB4SNtKBXtFAg/T25PLG4
Jawj1lcjWkNtTTmT4UK5VPKkQMuyHOW8IM46D+SmBS+MzjC2mz4hjcFGhrke/e5h
yVEicDLBNHSIllzgzoQh6AaAMnJ67qrpM354vJRrNYUPBetzCQXI0QVjRod6P3Q2
4iu7Biv8mvZRt3JjemkD0d0n+KhKFaQwVmDSN2B9Pnj3TGMj9ry0NqRyOxK7oPUV
8dacF9Skoe0lSG/f6o/IVWraK3OYNrpDTy86M2fHcn95UqkY/00K5RdciJPFSkEO
LRSLuHqssEy/FQz9lkvYh/eay9FTQmAAp0PKvyEDvgfcfA2tueOmP+fYhkpTCzwQ
wbRzqLTOm5K5tJbIyoKto5Xf/gJg5mwwDUShTA6UYoAtS8VN6bj7APc12k3h2fig
p5zPzd6EoVVT9iqBL2ItJF9Xm9kE9pMbjd2+ZVdoDzf7ac9/c1SoUZ2Pujcx17Nn
XPQ4ljaYalWzM2KXwOwmx1dg8QXsZ2JUTxxM8I4tmx1rNwL63ElPb6J1De7bKt3/
/fh382/QUhbKIMNn2LcuKZ/UNtWg+PX3txvl9+6McrgWwjmPXEUQaOhEM6iOgiwC
PYE8kjyHC1a7NVDsXyQU9ndjU1WIOgBwKJMqA0ztTLpGEA0DGN7hgfZ4szWhKO0e
Ce7hqhjgTEC8Ek9CDtIXTY2YB7KY+mdWyJ0xGKYhTqFjj3iOe1GWX1+HnahUoaWo
kgcydJhWMcvN13XvLe1XMnmWYdBvLjKTc0Iw/TCZk0WYOwpaKX0UmI+Vquwh518G
Bar0JZLZMtSBjKQXsg4FoWvhTTg+6iXcUexdoUmYKk4pIeoiv5oqkYpVi6WELH9h
+HVo3ZEQPLkIOwiRWdCdvYRx5cCK43cbWnYRNukXlVav+GA+c3JJgXoEUXCPZYU2
kKnGjp4vX6WB+UvPzgHUJOy2lscwf5PnOU6gL/iLs4wJuqJsgjLI6neGFeh4MIYc
zL/lz1oc4soqzfnKOy4DfMM4SH0wdVnAu8TVe7fQWoxkUin3vIw2B2LDqWfhrxkL
48ieGoNjUfsqA+E13cF6DI83AIt6ARHlUeRG+SJHk+Dv47so2kvQchQPG2sUF1jP
iwE1pa/T3s2OHMJS00vGSumxEwqbWsMF63UtO8T9HOSwewxrA3Z21f92YVPiBF+i
CA0BWKbiQUINxlxm1aXBMGiu/wiDtAL8rpucnG9we8lDU5pH+YhMCGyT1ydZOSIr
44pwHBEtLNr6nxlU25UcABlRAP8xv0h4ki02E3FTXwU0WmemtQuD/7QfXZ7e1imO
o4+26vo85A4FhyheBVtMJ+wC0TzRv6mQGo85pMUrwFaQ27IIAV5mf3wTFsFNqie8
Vv3tYC55CA8LMWI4Smk4qKmAwvil43yrTqnJgxM2c1bp9QWiGG6Cjn5sYHyFMJ61
aANBtx9po7GJKehstniVIsm0Vls+GHuD1ynE9Nvvl9P+1eTQ7lNAN6+ug8j1MsV4
DCu+xcQneSXgr2UBOL4wtjaMEqAa7LJ0VXdDO/x0KMVusvRtcW0CZ7xl4YJXORgy
//8rHwEKTTBYGzoV5t0HQtcRNA9D8t1epXIN5D3c6kcMPb5T4xW/EHD9AsFw5qNQ
4RGQk2/+r/pX+fzRREs6dbDUG0Zi4ih9J3ctkFgmXUMSa+DphRAg9S2n0+pO4PQS
xACw/tz7K4b0GUmSDbWU97y//9I4MP6SpqvRUYqdU/uosALG4lFV7cOusvbPeAVV
R+2RBg5oquYSMqnoGAgrzTzIeWRWkVZmAzG5w60Jsi9g0QwTgCiy4xsuWI6eQgPe
wrsQLN3Upkhq0C5eRmR5iGsZs9y5+y94v4dKKn4ST8I1u/GVhPok8NlLV+GqV/BE
T825zH7/7vyAajQ5LUX79rJEHC4rayd2zyl64tp9p28CdflPWk58o+eHA5rIX96b
fBGqvj+wXWlX39rus7pHQvOOSZUjBpmHfhHTFadY1QtrdTI3twYFQ8NmMCP6T27L
A6e8ty2cEwUXJsIVNFggTau1YpMspdJcK5ZSCnaSnwICuZ2epDFmWx35IhgtXynn
DUuicYHQHzU7MSxQ3qY2a0dbLqtWKSG4r/2BO/yoi43xCrH7hBzVkXI4ET4kHePO
CNIOoNhYvRdnxDpQyuNqYimgG8r+hC+bEbFya57cAbmfNYVjK1cJYkuulJWj3VUm
SPymcIILblAAPte+H6XF5ZTXswQircJtczrXdmybQ3NZswDsbsRpJwXlpHCxtb3a
+MOOkwf2Tuc4RNZTbWdo/mMPiQZRnXKD5An2i2v+5NbVHW7O53dWIQJGwfDZ9VCI
izGg6Dqc/Lj5OxU9sm9rHod7c6Nmh0DSfNFld7znj82dVEN+ehePhY03wi4xEkyB
ksUOsPUP1HpmtChFfbjdQTLWSm0Z9+e3kEdrtdCZD7/PhQdM7t+5aRRoHkTc3g6/
i7uexrpRb5+MK+ca/8ZFl2qN8HvmcWKDUDDC2P+buAnq2PJnr5YgXjnV5K4nayh3
MZ6ApRhaDdpfr3+XJRdwM86xm2POjIGJLqpaIbA8wWyk6PflAzy981dH9LiYG+u9
QHYx59pISgIaW7DLbLh+74OFXepbucCerTXhYs816Iq+4E+43pLvs88x5RKeQfSq
9McRwzHtj8rX56s9gzlbF+EyHSvLsslUE/1O9nhcUt5/GQsRsoZd2Kk6JMSAKCp+
F7LN9OJbPMVguuQlC1b+Oy5xf2D7/YZZpAXsVtRtGzk0At5lvHwZsrA6swN6sI8L
deW2gusWPVuvIvDYkJYMVSRwiJB5sCwK+WGvYuR8UWHbTtsO5aSuDU3Os95CsPC9
IuviG9j5zWmXlspALRxnO5d8X8v2u3kHBXC4+NZVCOJaNUNVQ49agxokpwNaY2hr
MI24TUMvQlPwQkSveogPpXI6UDv3DS5ltNP4eBhNNF9rg77SLhsFB7aKMDPRFj7A
Of4MyLVClopAF3QM8u3GRgZqLhsCB/qYUSppY8cFDgpx0vWYFI4f6uru9F8b5KHG
yWUXokfhZDJUe0mXLUNfNx8WfUO4fd4xhr+9XAeOThUywmimpssjWED7Lex2N6Rc
z4K2i6SHDflA1qQqyYntdOMlMxi+Lx9OfudN1FIj/8EocahciUO9NOyScb9Vvryn
6snXGurde4pfdvBcxCwAzj3yruadua77y1jCb3QpEHQ4L0m7SCBf3D/z9Dpr6fRb
pEqNHkcmwWHyGOlUBA+uVbbD9F3smVgeA8pA2vUZfZDpMosDVLa4tDGG6i7dhjWP
CCjgxWN2tuPQpvvLm25ue2ulBCSPPJaqGwcMJmK1EOFzN0UFOAl1rwJCeioNfxi1
S+kmmi5v6IYuHFNHmKu1GqOZLcv0U07pmAyUB7d3BWvpj4ofrCKtM0NqJ1py3wzM
BmgH2faJ0JENOearoCh9XXZbUlz0mABm2rzaqSjPl/QTZ6okw9o50VEZ00/CNN5+
oFEJ0zb45OQcS6O9VdjklvK/WqJVoRw2GRfSVMrNfxsdhQKMW3DZ4MarsKG2/UpS
2Ly/mT3Ey7cLsrDyXN5NxJkaJFw2A+Sk2ZRX66h5BZ8ZCVrM2cKXmrHOZWwNxWbN
18/0cFGq0gmSaeNi+wKxqJJZs+S9+tpycAZYl1hTZ4UekvPEHdifHQ6wt7JsMHUY
bAwCFK3zpbnxkl4nrnytCxeJApUsXCl778FTV2d2NPU0B5ll/TEyn2rf1U/M26Zh
ia1X0wCaXyl2Ok2e8n64gJFnQkQjQ5YX2zCl0vsd4ETn8NEsvrmau2Pypvo8oHzR
4+V8n7Oe4sl0HP5uvCggUI/NZn4ZeDhkoF5pB4zTPL1DrzunPOh6FuNJHt1pTeyi
Cqt+joAWTGdDD/eEWSuIZVuqzZhEVbpFO88cN1Y5SkrdNPJYDBI4Shxf1jAfNX2U
CZQhvAf02WmQDNdwrdRaVTmK8jyV5oIacld8YWUScmvoBawZtAHdM4YH4ecNSmg2
vqliLt3/nhzDR1BrqEKWl3BDY69gXKM45kZprJ0knzxwTYAh/VFcUuoheYsLKYPQ
26sxB1QR+jWIWDK18mPAwLPhPF2chKBQPb61I9xH1ixStnSSv5Y7h3b4z9jJLW5V
QcDARHyHdcQw1Vhr8FEhYzYqWw5iswN956UibTHlCpPrchv76tUHGyiR/+AfGZ29
qEguvuWOiBxCtsh5RpCM4YsZUBe/hnNKRp7i3WFdmG8QDGb5q3CY17UIo8cxZPkW
nL3d1REy4DDt+MwXNDzLX5cK++bhFlF/kLcw+FGN7FrXzF6kJRokJcMdWnqALuaY
P5XFWR7bVQDRZLjjW186hkCFs1XquzKZo1V+8EUFk5Ll5ibPmKZFyFcMFLWj2BQP
A2Tx9+IqTWT/cpa0flnfobic5liE00tMKWxHJAxrjPSytWC50sjCRmIUaoc840bS
4pOnKfTn8pYIN0kVAXVTz6PWvH9ZDEOUOAY8xmx1t1XKxpwxerVtH99doUbh3mlq
jOVvZJLD/rkFCqtTgvG85aQd2up+ciszxc5231fSYODspKrnOyv0GFx+3P0b/dyF
CEvnyV5Pdiwe5TFlgtZtQ8MUG7emc2ZRKA+5XxLUjNUAuEfq3eEcZ0NwsmOmZnm/
2kBJLO3HcY2AE9fzXjqnvtVF4DBa2VtpFXO9PlW3x9Xam6m9J1uMfbyeq9JjvXW/
UEPDEN+38E5jHmVf7bN1kbqGBsxjFxbt7QN+HVAZ/1fG6JMG+gX5rR2HsMxWZ9Ld
rKqFMw7t5mfc51ei6xQeeQ7hIZAMs54D0Yl5OibvSwQUJn9ISTfxgzT+517RpZ3F
50VPURlzD3PLQ0iKqFSK6Oqfps3QYaRpgLfpOwsqEiTOwQgz7+6JU1V8lfLOp4Tn
TM/pryFhQE3iTY+oJSB86nP3FcRLpLVUUleVrFX02VhF3eemFFNvwTtuDN+QX9LC
9STJ6X458Q28UC0YODo624qXSjV8/kwgVYO96oHcNAb0MQtLCrx2i+2QTPAKsuRo
TSZZuDNy3KzxYDf9GLeIQqGG4FvDizSleYfnfsKzvHsLS7BBUea7ZOscjRqJUoby
rSbzUqq+i9gOk5bfgCjjEaoS1kjfE7nEf84gA3FA0ohsRx7hX0n9+DqrMdn8xqw0
hoYm+mroGVPSTkU6Ex8BbmhuryGzuRUaXZfSjftmYx4mnA/G82H4LsDXOo6j8J7t
4dw+5NaKBesWvwYbWxypjDXkdKY8eSvlFiPY6v3SQHEGUnpyPqo+GSSgm3uiQvv3
s35QbqSaSZmWdb1JN0hRRgKbdvmzxjvS1+HSTgO1aq5JSKXGhGWSdmL+rH5HeTBj
cfBNMcjcXDaQa8Oj4gbMmaQbuOqLHeXdK41+034Ik8LWVBAP9HCOH52ibi+NyHNv
mQetEMpS5QH4gz5zA+n3WD0vnmRbRe5u9AVSc+uyerSQeoxvP3jZevQwSarxhQsE
XqLxuMo1cW5kQLW2oOOl6/pS3RHjzUIoC9Mnm86ruF07uWFarcJRBIfjFQkHyt3Z
UwUGPGJZ9BoMfNApVI/lumd0Hjk+1z9mbRH3FSmWAlTt56a9dqod7o+NK2mv+1nb
Sox6O1tjqJD554U0mc7iXKMAXpTCOx7IZEEIAhYh5HfqBO0cRUUFCdBxMRDDT5XN
qqaDB8qVi/SADG0Ssv3v+doddOIotnkFvzsHt+ZmOj8iEasUcvTXwNo1MEva/bcm
7nvWtWtUedMQlYC41lxv7hgJc7jqjl5iIcuK8FyvF4gieu+tNOVWBMlouo8blJXj
Bwt5kORYp/xg7Hl/RVjVQ43+6IDccD9Hq7FXUOokiWxZmGdn9KbFNLKXKuD4PpGP
E0ahFoWKxYmq9Da1Q9N17riUutsoGgcbnzkJZudHVEFxNTB/1b7suXERZHRsvgge
m8y+7dJnaS8qCkqGi3oDKszAZkn7QakSR/KHZvoXH/gP3nwtO/TaIOErXi3ZvdVd
DPtwrozgzUToGrVZC2fAPRiTlXDEHyZpoz8cNY5zqjfO8i2V9rhsVLs4r3q6Myg1
NIDbg5WdTwM9ZAGenHEiX9F7/B/l4fcv9cnwXa1jcrTz/F7FElElCkdY9Cqow+4T
GIGKOF2IZw7LEcHVOzi/cYzjJCm3beOFSkYQgUBvJ1KMTGbThUSwQ7fUnuU6wDrM
XOPlRF4Vhq+M9zlkW2E409D7I3UE+siST0jOBOKcH6JxLtL8YhZQRD6JjBMAH52o
9ptY9TyLml/Yhg2rj1rER/dVppfmDAmnlHYVeq4BBKnZGMBlWg4kc9aXtc4geIYy
yqRYzFF0LtVKnUsqxu3BUJhM9BzcwhJFZRAnsDCnZW++ctKXdelDcI/LbE0IqfzE
ay4QbwhOaZxfrl4Fwr15u+MkaHVEJkjxssxBuosNB5Kv09xqEdEhPj4+AvQeuko0
uw9MEqH7HK5OCqpBhms1v/k4TRIuTMnw201pprxk4pVxE4/i5SX9OhLR/YSYWkzj
AStEYWkuEUFuTd4nbDeQJWcE+D/43bY/WbDCcYl8SZrQr5QE5yORZsFC7atcgwja
zShEZ44qA5tQyrPH80uYSmVtGRzv+QoWw7k+81sEg3xJBU+fgHqkdshYLq0oqXOI
p+LSlV1DBO5o8Lh5nSpUX+N98Aviy6dyWbGHFI/ZIiI4gRcw/+TFYZ0222m2J1Ms
Cd0hzA0Gw1MH4i4+pvwqojc4plU1QsC74sCJW+CSXDpaq2P1+ES0M8oKm4r+ufHV
Qiw/SoUg+BwBIKuFnInoIgaTTF8BqgwjL0ZqqCS+f20NBJVV9Km5QjEzy2g3YuP2
d6HnPTWrpoBPF+bViRjv5ptTzcY0NHmos3t7KI7NuZJjQTO3Rf8xRz2guCYOvFVS
+boV9XNVizkxtURRyjkOssUc2jQ7+eDQJ0TvdijfZ0wMArx160xxd+TQ1RmU4a97
TGEUf0cnDqU2O3WwjJo8Fj9KLI+5y/o29P2PbCSzmJJzW5xEF9mBbWvvCdNk/cNB
+kavAXxOXkfygTEP59qRwKIgUYtWP9slgpfmxPF4B60NEQMVCsE65uojAl9Tarwh
JCGFUkS14OXnE/gXWiYMn0VlFoPPjgZlhBQgpXwicOnzHC2G3YkuD254s7KzGhA9
r6SdvA7XNqOw4AhM/nsnLwZdvuBtu+VYWDo4eUKqUmcIN46wvpsYqFwQQysylDlg
xk7xwq+M+f3XlU4D3HkCRK+1PmTFtVvIaNnjzqM4vwUhRdx719iXYPNSowGQ03u+
VVK2RQuzkLYvW0hGz2MT1pcxWiRoFC9dX91lbPHI9tzEghh5xWvxYzFTeIcrR9FA
RzUclwtUCJXmvMV0b8kP7qGFuJ+FsFnIuVvJdwQXjp5WmHZdUrn5nc8fem2WkYIy
mx0USYquzScxApXAHbtIIK6eiooOp4TPWj+NCH0S6uKwEU1AjiqsT+Rmx9pnoM5Y
ODrtQ/h/Jyca5eijczZlc0JknOYo/K3z3OFVbCnkkkJ4haddTDq0s5n66rXfgVL2
F6NsoQuRcm97vrizkOFXBLwJAjHidHaVV5e7AnCSkgtz/NXu9fxDlbhf0eKhMFMr
64XBDSzvrbE+mDNmnZAMCZBsi5eOITOSQ2yVTacjSS2STx4BaTz9OLhD1kipdOJC
Ud7Fs59jwQZFcFdSx/awocWVL4E07yvxhdYn3SB/vLi7wqnSLlBOFnaZVYF4aRmv
oXlLiMfLhahy75eEN0YIQIYchsRF/X/CacfHHLKOpqgL8tPY8ZYy4dhJl+DOeYAx
QAzEt/eOSSXhcd7qKPLB6ynjOxekeOyzqt7HOfTfcZBVy7P5AvXPvE8fO1Kt5X3F
oBugyI6o4LqBLmGHZlVvyya25LtAxzOa6v/mDL30E1ynOEDhLIW6CYjkfCNVdexh
MJyvoKTTESADwuSiuxHU8Ay6+pYWRUXaQohtCyA8Yuq7s/oyLLHfwfWcxXX5KXsr
cQBkaeQeOl/Jw4yQVInKgNg2dKIq6SvUBhU8W8SC9kvxnllS7IMOPs4J97cN5b5O
5KY9BH+WB7gtBW2x9y0nFZCjXY6DgigYmZqiMRlxgyES0CY7t3BkwbBEE1e1Pt56
vT6azkncrKaNyWGzinoqG/cxjX4H0VXRaUYXYQsegGgiwylpEYnLSiWTbydybQNd
WNUnYifnPupQmYP+vNfJk5GOzOWPZGDSrw/zW2RT9TIHLpHWc9bu2Aum++H4FskN
sPdqolBp7QbGD9DpnBQGL8t2TjJPx15tiiLTR9YHwlVxfBjZRqeurridCf4cCEC0
0A+u5qXxYM+ksXU/VHSic/mL4qcgGtgJrnrlcmzBbWo4+AfLf3huSqZBCZFiaISc
lIHi3UOWDY1PO0GP1++WHL7RiNXWqGDBbJdugki+Gk20LpsTGlu2ot9LHx2cWPZr
BGHp2wuHVU8thmuveehYLu3ukRc0Xg/ZWQ2WtK6cHqYG8dLCSb1GQRxL+GA+h9KB
/8nnzuGz2Ru+6tA4aeT8lfbS6VyZMy5HIwkbaV2t/wd17kTaljqB16p9sh7DQwCN
4lrqRkL6nf41aMTahZbRMQOAHrx4vLEdSMJ1zgwuLQ5D/mXtYUhhBSXOgle4gAMx
7xetMtw6AKN3OLJlFs+VSzt4QicgC2t7oSz0NqWkTvgZvNgAMp8pInFpI7Y7EcIW
/anNqL7Vz2y8+vYHw6JPRJDq6B7ZR6MLrZPSgHeG9oY/YT2IelnNE/3+UD2TVBA7
DxSxTM1KGrooGKH5W0T6VaYeFGIXyApPUatPvpV66KDDg26htybNEjTKxcBSDaGT
W7CC9JX3X84/f/+jw4FOim+XIQFiXpLnbYUeX1O2nW5pSikm0Q22KeuwRhrotcSz
9CphiysXymME3PsaB6yYIdlmoBf+dKGO0PwV3pJjNmlFxmspdcvHyhfErDsDC6hW
sF6F3BXbv8yEP1uAL6ht+veKLLBLsKDL1WndE5+PFESb4CZckUV5r4O/lwoeCPSi
QwZ0jEySqqcJQQCpF4eEqGRdAElkv9OoFat+DxQKwhcPlEIzCPLz82gFPQaOlN10
6Y4gwKADYEn9roGoJ9TfCVk6oi856o7R/WIIJ9bgh/xAuARifiBgEls1R88mlEkS
BcAkFB2pw0BIFgc+VOboIE0Pmb1dEl3XwIIHWXUk2f/pz1Xr9NLVCvMl4+ArUZIh
UUJFXOkXJ8+ipG+IlvEQ1FXmBD5KkWJvfV2rybbCAggvspsOZwPFnC41YHT3bZcx
BVncxq8tx8C7GxgADSq1aRzbNMGXNwkwfaAE3ClO/6c2aGj72iEBK1USplAIJH0t
9hD7htlEsbY8yRVaKcAlE9dP+TDAU+EkDwQ9odoryNNBT1DeQoI2KQhNZjrc2G6i
VZWsFct/Mql0Cxvx19zDYT6mwEVzGn9iQGbTi8TfSCaxYEw8/OI1BTBZhMnM7KG3
so4+kxgbbHyC2Dr86zKMOGWeC9bGtAQlK/Ed6AToP1BXMPn8LZoS/CkgNaaIeHo3
Jm0vwjqr5yo+FGYDhR2gmnH/qFjHB9cuqyBVFn8iarD7QFUxgybL78CLHm+smPop
tJzzzGr5qDSoTACp6bfdBwnWc4L+sfzSLUBfGxfROgfBYLSRi+/g20rwLOMJRUzH
kDgwbYFbm2AG0o1HUddBFF+tdJuOrfUo5qHiUi7QOnCfIX/CZdb6USZ256lBURZZ
NWgFa/St6UN7VkXne+jKvk5rG153wy2P3zUHHthQFDKaG924zcMdK0gcT6gbBAv/
Xm/PCF+KGukoovkUCt24CvBYVkWkBxsVQTvxYbj74RgrxXaw3Ty9RCg9lWOaiYmH
huOMIpj0OhpftEER9f41JRwJsmmGqrS+fSYM1bhTTOdgby/eDlwfZgOHCKJJJyB1
fXx7CbF99nECsjvWJAsc2P6Vg8WJIiJfos56pcjIhzeRIjWPTMWwnGumv7wMnYBV
E7OFXhn0Lj6QTBSUeerlyMXEuj5oQfFxLiOGsIYA4X4tgMlqlQZkb24K9hpIVm5y
Y2S8nBKvWPnncyalVMrZ4nTEDh1z+Vepd5RNyLz1mbhNNcJRdxAg+zJfkaC8lF1s
AUsA6TPX5LvrUDV4bcf7LVVM3jiRvh/X+SwVdI7mOrbh5AzBKm4YLd8cuWMZzC+l
4wtiwUL+gV67iQWqpJRwesKXEnuufLvgGZ3qOmWrpqnWltqid+N9ob4OKhW6VHlR
LgL1BPlzXyQqkXG/57C93sIMWLT1jWfu3Yf89bH5uFcOBaVYpF4pj9ux7Ykea3+k
Jz4WebR7Bn62MDkuGgOhkYZ3A8abnr9N/rn+Gpo6Vhge/KUUdr2m2xVWc/7LFumS
1HWMSQVf6QYPNPcxHetfnKAfeYorkRzeDE/n6EeIQet5oI9Z3stZoyi0xmSLrCLf
SiECe+483MGcYCNfRxuhW6DLQ475UfZ5x2JZ1sRAXs+//hHdiVVcTwkYLCxneQoL
eOmGUycb6+wO9WNhHdRi29S+btbAV6HZbqQQAzs2VYaeYoqyvY5aaDa+n9Eh4HSr
CTlRujEoapyWs0yLr7jzjNJf8TfZYEHRfyF/LUtKnKIaEbn/C/eWnWObX0/G3k4E
T6gMbz2lDwE7YN/p6BS5XGblK7itgBXAwYAsCM0/SEswscoNDc+kDX9+z2RmLS9f
X70G61r0f+KuuiAe125Vk82JDkq1KE5XdxrHStIxVqbkbbA6IIuFQCZAA6DVaSdj
+iVmNGMy3tqnCaILYiNeYHtlxIsMMG0zLejFl8QrrwqNnFIxLV6PMeBwibDadGNN
LG+HRdYZtsNzrjNogn9ZnlmRGqqIynOT3z7V8n4mVtrqh3jPmAJsUBcHotPgh4la
Q2xrA+2x9o8K8Oa8CeTggnvWOCoVZgH8M5t6Qaw53i1Y+3MH147AkRKTrZ2zvIOC
5jjHs2pB0m5AQt244JZHuRwrbPbRMdMKfFlJzlQWgp3RffFFdQZLOqhIuKC7q6MM
Odj9T+d254sZ4EsPbjzp2+7KhI8j2DrkJeds1C7Cvhr3nU2b3/KjcyYa0VwU8fRt
XYUdJYSLUzC4Pvj74eq27B5PPLSnYVpQI9Z3oNh8OIJ281wELYEyly7KaxV5JVda
qq0GAWeMC6/fBH8ZTfuL1K2VaMLhCBtHk2DPA6263AriZ3P9RSCCOC0N5T/7ZGJH
GXpLuRZhiRGDQb3QDg0pFMP8h4UpyIS3TFp/S2r/uPSqr5jghuJVKz4qfjFrufjf
u73+ZTW798k33B+6qzbq+K4IsykhJdxS3la3tF0RD+FzSL/sGdiAn30MMq2AztAr
ynBpIbLcomC86nRvNw9rfYIN3/7Ry5yhRaT9FznCSASGX0hKZBEdCb2xTB0yiPyD
2ACQK8b5T5K4HJ1773DIcT8u/9GXidIL26dZVkO7o1ygrZl4n4D97MDjH7r1GH4M
bVuJf2qSftfzj3e7SnVRqA0TAPT5d8XQSmfgS9mkg7ZJRfp5pCEp6BCvIJgOql28
5RskM66EaZe/KycEc1Tlfxxgb208uW2C3Zw8p/bTZWQd8db0s/DnTV6TDJEQ/O44
Z692xBI2qfAXj/qIK0YYk+V0ibZgEEUJZTVAgxevga/rgiW3h7+YjiIelPGu8RhC
IXeDG79vDlOsC0m5/M0unnk42kSmWKiL360s9BoI3xtMDbUnyqL/tKY7xWg2LFEG
1c/+q6es1nLwYyDl79FCCBfCnwQeG58SB66DfctqC0efPhixgaj+bgvHvfz1ncPP
JyLsQo613uHaXS1fSbor5WdZ0VlaZP4w5I7nLuh6cPmZUpU5B08Tmw6dpy3QJGf8
sskaPsCUTwZACDPMcIuAVin8OV5WKjn/4WziHcQcaGd3xmXlF3BmbAyiTeyzm/qO
A2mmeHMBthYQLbMHp7rzzizLbcsYkul6V0ZC8QFZu9FzukMHZSMhrOGJkq8uOYce
EqlNC+KGgqi6p4yyAufDwz0YedlZTxIMDRECZjgVBL4ua9ULkoFI9CdTFU4qDRBZ
hcmSs9y4TBBgvKlqawBREaWNPbOpeLFOypdaEyC3qZC1dFckAw3zOxrZ/UKO8HXs
bWWEtLYTNB1ecX9eGwDvdGgbwNJ6c6BuSBGXzmUePdVekjeCJvTK9oVpQ94Og0JV
+CIMr52wq8jGwMXSFe0DllG0bbe14DcMIUQ3mQXnnNzA2oHFJneTeqtHe/mSumIY
+fnKy4v1xwOPl/UQhXFj+nFhFpe3vdwnMZ39jFWBLTCfMpgMuyCXz8tw3FxBz+vN
PsM9pKs9YS6bBeshuxH7pw6NMSlN88QgTu/Rxt0VfqT6i5vQ2mR6fRN+gaIlUaIM
qPXb6XdcZs0SbmMbwpx7WFlFInSR8haEeWlwnYO8IrUtVPHb8WuNaKxB+JUAAkFb
LetWkOAd1hY9TuGif6btHK+2yuKgZBaPMTjpeGPL4zWIpFSGCOTiNnibnctdMqve
ai1k1KUbkId3ciDotN3i4V4EqUmvxInbO1Ia0o1lnuaj850qQZQsoG4awiDDRfhI
RQyzQQsm3kQzV9V0Ap7ww5zRyC2FCaeROZTfjOmzp3sIEIQrysfyjpffmzA0oIQo
eJHAzC54KwloYwujg+ViZ+n567YizHeiQka1zTc+uIGlYAVz4DkZ7xwjRGDGxnZB
4yWUcdc5BIL9kWydRtVWs6rCtjTOkKDVspjc4ZT6+64A34nI3YXIv5g1XO0zFK60
t63B9qVxmH1UR+ZkBSNv63wLDsTcCrHwHs4aYRbJlfW89zNRqy5CD1al1jCZx/OP
kvMd4oiIb9iixx4I6QO3hJUE4wU81daTwOc3MEwrTJvXGjqk+0DoWzx2Vn9+l5ge
/863piEPBtvvKYvQrPugCwitLf9yC9ZG2jgHLdx29LKA8U+12VtinMebeQ3YOph3
rCpN5Ib1aDw6Nb4D3Yuc54EvgGDgeOCK/oGJIGxH/8RWe08ollq7XXpjy04XZjTD
OvGx4g0xgN7WWkiLhyKoDcn6vucaBDH6ODbVHS6IKpy/k10/yhHzl1aSMvXxeW5X
HBm5M3SoiFCMYXZikJx5D17BeXDuIId/PfwE8fdlmWkgE6meuly537gAez8pxlgW
v6fkXwlPHVNv8Z66vjO0GUAVtTcZQwnLY1BWSFY26hrDgetAOOytF0tON1sC39KM
tfcq5NYn+wVNeCQPov3iaCkUjUN/3QZPWJoa7dNu9GokAI05ElXOacQacEt4d2Fn
QKDjMSp6WmZ7z1fA2BrFy7IBaZC2bWiLgECPdVD1gS/ScCHiplB6C/VDyCXU3muU
IKK05TNf+7ryXq4USlQ3k9O3dZbEO/0rkRM5t8oQC67n5CdPh8nRWh1qno1L91IW
HEssS8VMXBVz9HLiaWpgnDt9nHnsqPM4RmFsI/CSoWdaSoMkyJJmJgFVDgUBKfYJ
yri0Rm2GWAlQ8lE0P7hjd2jdcAQYHq8+nUOEcWAT6bouscR/GKetnazgbGDscFKC
+AxluD1CEiEkdUaLzjOpA6Uaq/TDkRQCG22IkWxzkdv/gB6soiTy6muN2dGbLY+B
sSDrIiB9jnQVibK57Pe7ySmbhO/xm1VxYG4akFx1IdeWrDDMysqpaZcIM27KPzHI
aUmfmdxm4b5FAcLE0rPXhKrWqjurSdMb1qzCImYNa6E2D4m9cia4mo7BHMp52H4N
iE+5nxMpqY72LRD1sLyYPEEYXpmH5DR8B0PzOynIzsf/A+ZUOi8pHx+mt2qVOH/M
QSdVscQ+kndoWBQkx5tzqTXGgYwZAB62urIU8p+yeuuktB62JaR3ZdSTTjbgKQ1n
JO3uyRXAawZ5S0dL/bqYOAMNTNMXN75Ekt8FWoqOhoStZInGqSXPTZSPIXlw3WDT
QS5P9rWeuZNatJ30jfRmhEH8W5C+qdy6jW1L6GUV/AgZ4PvpckX01EbxxDMS1FoN
+8tDAvIA2jghRv8g8YZOSpZe/rMvCqUuszKTsQl5sx02UuyGdpSqSIHwFeQ3W9hg
fuMFJ8PHExwNIHADxKseckZDLWxEy8dsSm1jK4izqXtX6ezleUvGrl1enC0IkL9z
3F89mwPvrhVDHffLKlfZrRo1DqDEesQZqikub5Ey2+TSbpHEhwLBXp5mJX4ibVIP
q+zcZ4a1OqVNadH9pwiqpLZEO3bCWaXK2aTylkbyYoXjEBp3GSkV6d8AkwIR4SoS
jL+lkmWwuPahlNmpQvyW//GU+jSl1PGn/6RY+JkuIlrG2yZ05hitn0IfDng5+iIT
/cgW2PTTWYdJLTWpxNLSBxFu+6d2M3oP6/t3c9vP9cNcxsOqrC8LGf6QbzwjZt3x
XelSSmmNHpROjNycuNMzBnxxWpH9L7brbDCE3gFHUmqAlK76nNNp17xhP7crYLvB
+Ysvj7QTb+SIsk6ATL3BL4y3UVhlh+JtZiq1lFF9SdyqTeiOU6JB2mhSab+KsQQC
g5jWJYIuiCM5Xy+8TxvTqRlObVXhVT2BYwpbSGaDEEcsaHsbjxjoEeJxKXKj9+bn
1LPacjQ9t37ZwLKwR3aLzAno8/Te/fZE4TRrE/0Ooj/HGeI+wOFZD+VUJo/6NXWG
ZSTZSuJiAms3IkZK7l6z7RSckiGinRE0LnLepku2f/eIALg4KHvn98rzIfFfh5rf
Y8RbSW9PrGxDzCq0R4J9Isp1I1VBLkS5Pqq5vOUpjrUaFl/vC52dzlSJ9Vg8V8Og
chjTCUqwXYklPs1/JFVRmX3EYNy6YH1V9LdfUkrDtyYzEQVJTsrnUyDw+9fBArZ8
GZ7KOtEDw6E6qut2SQgZXaE/RiqZlSTuejLynnKV5c/DSia8gVFlZGp3YIiD9T0s
9dTWEQTSwac64w0FAVo7Ea0B+2fpFg/iTM/6OnKWEW8fRxoycd8TJnkiK+eWiWDv
rfAzCs5JCGf3u8Nadoaca9uIcVtLAXws+fKHd5Vfh6hDLVASzWVBQUCpCgsEVGCE
yWPAc0RrY3ydRP5x46Yk4g2R7q6folTRAhql9FkI/f9VlDWX33Im2jxekqsdEo9C
duwkBl3LmFjRF/vQi1e5PHe/J3sSFl/I6h9t0vPJyqdD0EJeoXvPtBiLCscuEMvA
ggEFc675nutuxmGdHebJ7fK5f0ePvfm2/wNxNzbRQtq2FRPqux70F76FoEfBKdrg
GOF2d+zGmqN0MB659G3kanQMwOBuVsribttESXNo32kHDrl8l6YOt7LCUCVQoxkT
lpZR6ogHI3N9XgQqpRJPaWruUYPUKaau1lVGdtWVei971w9kgNkTQziNxRn4BfSo
mcR+mcXnw/iaGvpBTVjKYblfVPYB0M2QWE3uj5CX8MgZcvyqqJfmrIsKtYghpD2J
uB7BU+XIJ7O7Fc6LQ8jpQSu8XnnED2N1ujw1KsQbBVWy/p5WzVA7QKJJnxNcVVzz
oh/u79gc8GyEjcwhzFk8zJgk9p88mdlXy7KrUQRXjBykQJMv2oWW65DTHoThdDLo
n/BUPHPEd/p4rQRej7OHw2/O0UGfrmBLz8MUw3DQpSP9WCL3BpSv+YZDk2QQ/eQa
n1gyxQwZhIdqYQ3Aj0TnKVdQOOTVB3LeTL7GwS4VFThF4G1/XK5DuM+dsdZ4F0um
`pragma protect end_protected
